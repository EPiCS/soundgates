../../../../../basic/add/add.vhd