../../../../../basic/white_noise/PRBS.vhd