../../common/soundgates_v1_00_a/hdl/vhdl/soundgates_reconos_pkg.vhd