../../basic/square/square.vhd