../../../../../basic/sub/sub.vhd