../../../../../basic/adsr/adsr.vhd