../../../../basic/sawtooth/sawtooth.vhd