../../basic/sawtooth/sawtooth.vhd