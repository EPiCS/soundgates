../../../../sndcomponents/nco/nco.vhd