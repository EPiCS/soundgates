-- Derived from yay.raw
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity SampleDataRom is
Port ( clk    	 : in  STD_LOGIC;
	  	enable 	 : in STD_LOGIC;
	  	data_out : out std_logic_vector( 24 - 1 downto 0);
		rst    	 : in std_logic );
end SampleDataRom;
architecture Behavioral of SampleDataRom is
	type rom_type is array (0 to 42678) of std_logic_vector(24 - 1 downto 0);
constant rom_array : rom_type := 
( 0 => "111111000100111101011000",
1 => "111111000000101110000101",
2 => "111110111010000100110100",
3 => "111110111100111111100010",
4 => "111110111111010011011000",
5 => "111110111100010000000000",
6 => "111110110110101110011011",
7 => "111110110001100110110010",
8 => "111110110011101111110100",
9 => "111110111000000000011110",
10 => "111110110111001101101110",
11 => "111110110010011100011011",
12 => "111110101101100111000001",
13 => "111110100111101001111001",
14 => "111110011011100011001001",
15 => "111110010001010110011010",
16 => "111110010000000101011101",
17 => "111110010001100001001011",
18 => "111110010010011000000001",
19 => "111110010100100000101100",
20 => "111110010111101110100110",
21 => "111110011000010110011101",
22 => "111110010111011001010010",
23 => "111110011001000100101001",
24 => "111110011111100001010000",
25 => "111110101010100011000000",
26 => "111110110000010111100000",
27 => "111110101101101100000010",
28 => "111110101101100011101101",
29 => "111110110010010001010111",
30 => "111110110100111111001010",
31 => "111110110011010101100001",
32 => "111110110000101111010011",
33 => "111110110000001110100011",
34 => "111110110000101000010011",
35 => "111110101110010111110011",
36 => "111110101010110111101100",
37 => "111110101011101000011101",
38 => "111110101100111101011000",
39 => "111110101101010011001111",
40 => "111110101111110010110100",
41 => "111110101110000101000110",
42 => "111110100111110000011100",
43 => "111110100001100011101110",
44 => "111110011111011101100011",
45 => "111110100111101010100110",
46 => "111110110011000111001101",
47 => "111110111001011101111101",
48 => "111110111110011001110111",
49 => "111111000010111001100011",
50 => "111111000011110100111111",
51 => "111111000100100100001110",
52 => "111111001001011101100111",
53 => "111111001100001001110100",
54 => "111111001011000111000111",
55 => "111111000111111000110010",
56 => "111110111110101101100000",
57 => "111110111001110000000111",
58 => "111110111001011010001010",
59 => "111110110001001001010110",
60 => "111110101100111011111001",
61 => "111110110110100111111110",
62 => "111111000000000101000110",
63 => "111110111111001110101101",
64 => "111110111010110011001010",
65 => "111110111101101111101010",
66 => "111111000111110100100001",
67 => "111111001011100100000100",
68 => "111111000001001011111101",
69 => "111110111001100110000001",
70 => "111110111111011010000010",
71 => "111111000010100011101011",
72 => "111110111100110110001011",
73 => "111110111000000011010011",
74 => "111110111011010010110101",
75 => "111111000000010010011100",
76 => "111110111110111010001101",
77 => "111111000011011100110100",
78 => "111111001110101011100100",
79 => "111111010010001101001010",
80 => "111111010001000111101110",
81 => "111111010000110101000010",
82 => "111111010110000111001101",
83 => "111111100000101100111011",
84 => "111111100011000010100011",
85 => "111111100000111011011111",
86 => "111111100111100000001000",
87 => "111111110010001010001010",
88 => "111111111010111111001011",
89 => "000000000001111001000001",
90 => "000000000110111001001100",
91 => "000000001111100101101100",
92 => "000000011000100011000100",
93 => "000000010011100100011001",
94 => "000000000110101101000000",
95 => "000000000100111000011000",
96 => "000000001111010010010010",
97 => "000000010011101100111110",
98 => "000000001001101011000000",
99 => "000000000100101011110011",
100 => "000000001011100100000000",
101 => "000000001111101110000100",
102 => "000000010001101101011110",
103 => "000000010110000010001011",
104 => "000000011010010110000011",
105 => "000000011101001111001111",
106 => "000000100000001111100001",
107 => "000000101000001010100000",
108 => "000000110010010110001011",
109 => "000000111000001110110011",
110 => "000000110110100010011110",
111 => "000000101111100100110101",
112 => "000000101011010011000101",
113 => "000000101011000001101000",
114 => "000000101001101111110111",
115 => "000000100100110011101101",
116 => "000000100010111011101111",
117 => "000000101010010001001001",
118 => "000000110001111010111010",
119 => "000000110011001000100010",
120 => "000000110011101110110110",
121 => "000000111011010010000100",
122 => "000001000111100000110000",
123 => "000001010011001101101000",
124 => "000001011001110101101100",
125 => "000001010011001110111011",
126 => "000001001110100000010001",
127 => "000001010100000011101110",
128 => "000001010010101011000011",
129 => "000001011010101001101000",
130 => "000001110001010011101000",
131 => "000001110100101110011100",
132 => "000001100110100001011100",
133 => "000001100100001011000111",
134 => "000001110000111111101011",
135 => "000001110010111000001000",
136 => "000001100110100011110111",
137 => "000001100011101110110111",
138 => "000001101001100001111011",
139 => "000001101111111011010000",
140 => "000001110000110100001100",
141 => "000001101010000101011000",
142 => "000001101011100111110010",
143 => "000001110001100010010011",
144 => "000001110000110010110100",
145 => "000001110010110001110100",
146 => "000001111001111001011110",
147 => "000001111011101001011011",
148 => "000001110110000001001100",
149 => "000001110010000010001101",
150 => "000001101001100101111110",
151 => "000001010111010001010010",
152 => "000001001111110100011001",
153 => "000001100010001101110000",
154 => "000001111010101000001100",
155 => "000001111001001101111100",
156 => "000001101100001000010100",
157 => "000001101100011001010011",
158 => "000001101100000000101000",
159 => "000001101101111111101001",
160 => "000001110011111101000011",
161 => "000001101101111110001001",
162 => "000001100111010100110110",
163 => "000001100001010011100001",
164 => "000001010101000110110100",
165 => "000001001101001000101100",
166 => "000001001011011010011000",
167 => "000001001010100101000110",
168 => "000001000110010001100000",
169 => "000001000101010001111100",
170 => "000001010000101000111001",
171 => "000001011101111100111100",
172 => "000001011100001111111000",
173 => "000001001011011100101001",
174 => "000001000000101111001001",
175 => "000001000101100011111000",
176 => "000001001010111100110000",
177 => "000001000011110101001000",
178 => "000000110011000110101001",
179 => "000000100100101110101110",
180 => "000000011000101011000110",
181 => "000000001110010100010100",
182 => "000000001100100000111101",
183 => "000000010001110100101000",
184 => "000000011001101011100111",
185 => "000000010111111100110110",
186 => "000000001011010100011001",
187 => "000000000010111100010101",
188 => "111111111100111001010111",
189 => "111111110100101010010110",
190 => "111111101011100101011001",
191 => "111111100001100000000010",
192 => "111111011011001001101000",
193 => "111111011011101100010100",
194 => "111111100010110111101010",
195 => "111111101000011101100011",
196 => "111111101000110100000011",
197 => "111111100101100010100101",
198 => "111111011000110110001011",
199 => "111111001011101001000000",
200 => "111111000111100110001001",
201 => "111111000110110000100011",
202 => "111111000011010010111101",
203 => "111110111000110000000010",
204 => "111110101110001010001100",
205 => "111110101010110101110011",
206 => "111110101000100010010110",
207 => "111110100110000000000001",
208 => "111110101010010110111100",
209 => "111110110110010000010110",
210 => "111111000000111001000010",
211 => "111111000110000010011001",
212 => "111111000010010011111010",
213 => "111110110111101000010111",
214 => "111110110010000001010000",
215 => "111110101101011101010001",
216 => "111110100111000011101000",
217 => "111110100100011100101001",
218 => "111110100001011010001011",
219 => "111110011110000101100010",
220 => "111110011001001000011000",
221 => "111110010011101100111100",
222 => "111110010001001001101000",
223 => "111110001110100000111000",
224 => "111110010010000010111101",
225 => "111110010111111001100000",
226 => "111110011010010111001100",
227 => "111110011110101110111101",
228 => "111110011110001001111000",
229 => "111110011000110100011010",
230 => "111110010101101001010111",
231 => "111110010101011100010010",
232 => "111110010111011011101011",
233 => "111110010101111000001111",
234 => "111110010100010010110110",
235 => "111110010110101010001100",
236 => "111110011001010001110010",
237 => "111110011001000101101110",
238 => "111110010010010101111110",
239 => "111110001011110010011101",
240 => "111110001010100101110001",
241 => "111110001100000011110110",
242 => "111110010001101010001101",
243 => "111110010111100100100111",
244 => "111110011001111100101100",
245 => "111110011000110110100010",
246 => "111110010100000011001101",
247 => "111110010011101011100011",
248 => "111110011111110001100101",
249 => "111110101011011010000010",
250 => "111110101001001010100001",
251 => "111110101000101011110100",
252 => "111110101111011000010111",
253 => "111110101111000111101011",
254 => "111110101110101011001101",
255 => "111110110001010000101100",
256 => "111110101101110100001001",
257 => "111110101010001100101011",
258 => "111110101010110101010101",
259 => "111110101000111101100101",
260 => "111110100101010100100000",
261 => "111110100110110110110010",
262 => "111110100110001001110001",
263 => "111110011110111111010111",
264 => "111110011100010101001101",
265 => "111110011111000000111001",
266 => "111110101011010100010000",
267 => "111111000001100000110111",
268 => "111111001000101011101110",
269 => "111111000000111110001000",
270 => "111111000111100011111000",
271 => "111111010110110010001011",
272 => "111111001101110101110010",
273 => "111110110110011010111101",
274 => "111110111000001111010010",
275 => "111111001000100000101011",
276 => "111111000110111111000000",
277 => "111111000111100100001100",
278 => "111111011101011000001110",
279 => "111111101101000100100111",
280 => "111111101010110010000111",
281 => "111111100110110011001011",
282 => "111111101010001110101111",
283 => "111111111001101101101010",
284 => "000000000110100011111011",
285 => "000000000010011100001110",
286 => "000000000000100011101100",
287 => "000000000101101100001010",
288 => "000000000100101101110011",
289 => "000000000000000111000000",
290 => "111111111111011100101001",
291 => "000000001010001010001000",
292 => "000000010110111110000110",
293 => "000000010101001110000100",
294 => "000000001011110000110111",
295 => "000000001001110111111101",
296 => "000000010001000000011110",
297 => "000000010001011011100010",
298 => "000000000100110110111010",
299 => "111111111111000111000010",
300 => "000000001101100010001010",
301 => "000000011111101001111011",
302 => "000000011111110101001011",
303 => "000000011011000001101110",
304 => "000000100100000011101111",
305 => "000000101101111101000001",
306 => "000000101110000111111101",
307 => "000000101101111001000010",
308 => "000000111100000011101000",
309 => "000001001111101100101101",
310 => "000001001110101101001111",
311 => "000001000110000010110010",
312 => "000001001010001001001110",
313 => "000001001110100100100000",
314 => "000001001010111011111101",
315 => "000001000011111110001010",
316 => "000001000110000100011001",
317 => "000001010101000011000110",
318 => "000001011100101100011001",
319 => "000001011010011111001101",
320 => "000001100110100111100110",
321 => "000001111101110000111001",
322 => "000010000110101000111001",
323 => "000010000010100110111001",
324 => "000001111110100101000010",
325 => "000001111111100011010001",
326 => "000010000011011110101101",
327 => "000001111010111110110110",
328 => "000001101110000110000011",
329 => "000001110100011101000101",
330 => "000001111101001011011010",
331 => "000001110010010011100001",
332 => "000001101100110110100011",
333 => "000001111110111110010110",
334 => "000010000001111001010110",
335 => "000001110001011101010110",
336 => "000001111101011101000110",
337 => "000010010000001001000011",
338 => "000010001001111001011001",
339 => "000010000111111000010100",
340 => "000010000111000011110111",
341 => "000001111010101110010010",
342 => "000001110111110000100100",
343 => "000001111111110100001011",
344 => "000010000111100011110001",
345 => "000010001011101011011101",
346 => "000010000110101101100111",
347 => "000001110110001100000100",
348 => "000001100100100100011100",
349 => "000001100101001010011010",
350 => "000010000000001010111100",
351 => "000010011111100010101001",
352 => "000010100100000001010011",
353 => "000010010111100101110010",
354 => "000010011000101001111111",
355 => "000010011101110000100011",
356 => "000010010000110111101000",
357 => "000001111111001110100010",
358 => "000001111001100110101010",
359 => "000001110111001100001001",
360 => "000001110100101110110010",
361 => "000001110110001010111000",
362 => "000001111000111011000010",
363 => "000001111111011111011110",
364 => "000010000000010011001100",
365 => "000001111000100100011000",
366 => "000001111101001101000101",
367 => "000010001000010111011000",
368 => "000010001000011110111111",
369 => "000010000000111101110110",
370 => "000001110100111110011001",
371 => "000001100110100000000011",
372 => "000001011100011011101000",
373 => "000001011010111100011111",
374 => "000001010111101001001011",
375 => "000001001011101110110111",
376 => "000001000011001011001010",
377 => "000000111111110000101010",
378 => "000000111011000101011000",
379 => "000000110010100101000011",
380 => "000000101100000100111110",
381 => "000000110001100000110010",
382 => "000000110001001010101011",
383 => "000000100100101000110010",
384 => "000000100100001110010100",
385 => "000000101000001110010001",
386 => "000000011111001011010011",
387 => "000000010100110010101101",
388 => "000000001111010111000010",
389 => "000000000101101111110110",
390 => "111111110110101000010011",
391 => "111111110000010100100101",
392 => "111111111000110011000101",
393 => "111111111110010010111000",
394 => "111111110101011011000101",
395 => "111111101000010110111011",
396 => "111111100000110111110101",
397 => "111111100001000001000001",
398 => "111111100000010101000100",
399 => "111111010000110000001010",
400 => "111110111001101111011111",
401 => "111110101000101010101011",
402 => "111110011110010001101010",
403 => "111110011100010101011100",
404 => "111110011000011101101101",
405 => "111110010010000101111010",
406 => "111110011100010111001100",
407 => "111110101100001110111000",
408 => "111110110011100110100110",
409 => "111110111010001101011100",
410 => "111110111011000001000001",
411 => "111110110001010001011100",
412 => "111110100000101100101010",
413 => "111110001100101111010111",
414 => "111101111110110110011100",
415 => "111101111010101111001101",
416 => "111101111000001100111100",
417 => "111101110001100101010100",
418 => "111101110000000000010011",
419 => "111101111000111101011011",
420 => "111110000000000110111111",
421 => "111110000001101000110110",
422 => "111110000011110010011100",
423 => "111110000100101011100111",
424 => "111101111110110111111111",
425 => "111101110010000100101110",
426 => "111101101001000011001110",
427 => "111101101001010111100110",
428 => "111101100111101011000001",
429 => "111101100001011100111100",
430 => "111101100000110110001110",
431 => "111101100111000000110110",
432 => "111101101110110000010001",
433 => "111101110111001110111101",
434 => "111110000000111111011010",
435 => "111110000100110111001101",
436 => "111101111000101011100010",
437 => "111101100011011000001110",
438 => "111101010110010000000111",
439 => "111101010101011100111110",
440 => "111101011100000100001100",
441 => "111101100101001100011001",
442 => "111101101110011101010000",
443 => "111101110110110111111111",
444 => "111101111001110011101101",
445 => "111101111000111110101011",
446 => "111101111011010100010011",
447 => "111110000000101010111010",
448 => "111110000110010100101111",
449 => "111110001011101101000011",
450 => "111110010011000011011010",
451 => "111110011001001101001001",
452 => "111110010111110001101110",
453 => "111110010011011110011000",
454 => "111110010001001010101001",
455 => "111110010011101111101000",
456 => "111110011100010000111001",
457 => "111110100000011010111101",
458 => "111110011100011110010011",
459 => "111110010010100100111001",
460 => "111110000111100110011101",
461 => "111110010001110101101000",
462 => "111110110110001100010111",
463 => "111111010110010010101100",
464 => "111111011101001111101010",
465 => "111111010011100010001101",
466 => "111111001010110110010101",
467 => "111111000101111101111101",
468 => "111110111100110110011001",
469 => "111110110100110010100000",
470 => "111110110111000001001001",
471 => "111111000000111111101001",
472 => "111111001010100100000010",
473 => "111111001010000001010000",
474 => "111111000101000000100011",
475 => "111111000111000101011010",
476 => "111111000011101001111010",
477 => "111110111010011011101010",
478 => "111111000101101100011001",
479 => "111111100001110000010011",
480 => "111111110000100101011010",
481 => "111111101011101000011100",
482 => "111111100110010110100000",
483 => "111111101110110000000100",
484 => "111111111110110011101001",
485 => "000000001001101000010101",
486 => "000000001011011010011100",
487 => "000000010000010011111111",
488 => "000000011011000000100001",
489 => "000000010111111011101111",
490 => "000000001011100101111110",
491 => "000000001011110011010000",
492 => "000000010010101001111001",
493 => "000000010010111110010100",
494 => "000000001010110111010001",
495 => "000000000101111011011101",
496 => "000000010100111010111010",
497 => "000000100110011100010110",
498 => "000000100001110001111101",
499 => "000000011001011000110000",
500 => "000000100000000110101000",
501 => "000000100100000111010100",
502 => "000000011010100101000100",
503 => "000000011101101101101011",
504 => "000000111011100011101010",
505 => "000001010010111100010000",
506 => "000001001101101011000110",
507 => "000001000000011000010001",
508 => "000001000000010011100000",
509 => "000001001101100010010110",
510 => "000001010111011000101101",
511 => "000001010101111011100000",
512 => "000001010011111001110011",
513 => "000001001101011110001110",
514 => "000001000011010011000000",
515 => "000001001010000000101111",
516 => "000001011000111001100011",
517 => "000001011110000100111110",
518 => "000001100110010101000010",
519 => "000001110000001110011001",
520 => "000001101100000110111001",
521 => "000001110100001101110111",
522 => "000010011001101000100111",
523 => "000010100001011101000011",
524 => "000001110100001101110011",
525 => "000001100001010100110101",
526 => "000010000011100011001110",
527 => "000010010100111101110000",
528 => "000010000010111000000111",
529 => "000001111011100011110001",
530 => "000010000110001111100110",
531 => "000010000000100010000100",
532 => "000001101010110100111010",
533 => "000001101110110100111100",
534 => "000010001101000111101010",
535 => "000010010111110110110010",
536 => "000010001001001001000110",
537 => "000001111111000000101001",
538 => "000001111110110100011110",
539 => "000010000001000100110101",
540 => "000010000100101111110100",
541 => "000001111011111000000000",
542 => "000001011100101111011111",
543 => "000001001000011100110101",
544 => "000001100010111111111111",
545 => "000010010100101101000110",
546 => "000010101010000111101010",
547 => "000010010110111111110000",
548 => "000001111110111000001011",
549 => "000001111111100000100111",
550 => "000010000111010011001000",
551 => "000010000100100010011100",
552 => "000010000101001110010000",
553 => "000010000111100011010011",
554 => "000001111001011110000011",
555 => "000001011111111011100110",
556 => "000001010000111111100101",
557 => "000001010101110110011100",
558 => "000001011111010010111001",
559 => "000001100010111011001010",
560 => "000001101000011111000010",
561 => "000001110101110001010111",
562 => "000010001100101100010010",
563 => "000010011011001101010110",
564 => "000010000111110010101000",
565 => "000001100101111011101001",
566 => "000001010100100100010001",
567 => "000001010001001001010111",
568 => "000001001101111001011101",
569 => "000001000000011001100110",
570 => "000000110010101011110110",
571 => "000000110000000111000101",
572 => "000000100110101110001010",
573 => "000000010110010000000011",
574 => "000000010011100010001111",
575 => "000000011101110011001111",
576 => "000000101100010000011001",
577 => "000000110100000101010010",
578 => "000000101100101110000011",
579 => "000000100100101011011000",
580 => "000000100110011000010011",
581 => "000000100010100110010010",
582 => "000000010001010011111010",
583 => "111111111011110010000110",
584 => "111111101011111110011011",
585 => "111111101011101011101110",
586 => "111111110101110100010010",
587 => "111111110111110111111111",
588 => "111111110000000011010011",
589 => "111111100101100100000111",
590 => "111111011000000010110000",
591 => "111111001100001101101001",
592 => "111111001001100111101101",
593 => "111111001100011000110100",
594 => "111111001100001000010011",
595 => "111111000001010001010010",
596 => "111110101011001101110110",
597 => "111110010110101110001010",
598 => "111110001010000110111000",
599 => "111110000101110000100010",
600 => "111110001011110101101011",
601 => "111110010111100111111011",
602 => "111110100101010010101001",
603 => "111110101010100011100000",
604 => "111110100100011011100110",
605 => "111110100110100100111010",
606 => "111110101010110010111111",
607 => "111110011000111000011100",
608 => "111101111010110010001010",
609 => "111101101000000100110101",
610 => "111101100101000010111100",
611 => "111101100100000010100011",
612 => "111101011100001000100011",
613 => "111101011010000100100110",
614 => "111101100010100010010011",
615 => "111101101000011001010010",
616 => "111101101011100111010000",
617 => "111101110001010110011001",
618 => "111101110111010110110000",
619 => "111101111000111000011011",
620 => "111101101111101100001011",
621 => "111101100010100101110101",
622 => "111101011011011000110000",
623 => "111101011000010101010110",
624 => "111101010100111010011100",
625 => "111101001101001100111100",
626 => "111101001001110100110010",
627 => "111101010101101100111001",
628 => "111101100101110110011000",
629 => "111101101001101001100100",
630 => "111101100001110011001000",
631 => "111101011011111010100100",
632 => "111101011111111111010101",
633 => "111101101000110111000001",
634 => "111101101111111010000100",
635 => "111101110100111100101110",
636 => "111101110110010011011111",
637 => "111101110000101101100100",
638 => "111101101000111011001101",
639 => "111101101100101110101110",
640 => "111110000100010010011100",
641 => "111110011001001011001111",
642 => "111110010111000100011011",
643 => "111110010101101100111111",
644 => "111110100010011101011111",
645 => "111110100111001101010000",
646 => "111110100001000101001000",
647 => "111110100011011110011011",
648 => "111110101100010110110110",
649 => "111110101001010001100010",
650 => "111110011010011011011000",
651 => "111110001011110000011000",
652 => "111110000110010011110001",
653 => "111110010000010100100011",
654 => "111110101011110001111101",
655 => "111111010011010110011010",
656 => "111111100101101000011111",
657 => "111111010100011110100011",
658 => "111111010000010101110100",
659 => "111111100101100000010110",
660 => "111111101100111110011011",
661 => "111111100101101001011011",
662 => "111111100000110011111100",
663 => "111111100100001110101100",
664 => "111111100011010111101111",
665 => "111111001100111100001110",
666 => "111111000111000011101111",
667 => "111111100011000100011111",
668 => "111111101001011111001110",
669 => "111111011001101101101010",
670 => "111111011110011100000011",
671 => "111111110010010001111011",
672 => "111111111101111111111111",
673 => "111111110100100010101111",
674 => "111111101000110001111100",
675 => "111111110100101100010110",
676 => "000000000010100011101101",
677 => "000000000011001010101111",
678 => "000000000101100011111110",
679 => "000000001001010001011101",
680 => "000000001101101101100010",
681 => "000000010011111001011100",
682 => "000000010001110100011111",
683 => "000000010010001001110001",
684 => "000000100001000100010100",
685 => "000000100111110100111110",
686 => "000000011001101101111100",
687 => "000000001101001111110011",
688 => "000000010000000010001100",
689 => "000000011100000110111010",
690 => "000000100111111100110100",
691 => "000000100111101011101001",
692 => "000000100011000111110010",
693 => "000000101100110001110110",
694 => "000000110110111011111010",
695 => "000000110100011101001101",
696 => "000000111001010000101111",
697 => "000001001010011111100101",
698 => "000001010010011001000110",
699 => "000001001000010100111101",
700 => "000000111001111001101001",
701 => "000000110110001001111110",
702 => "000000110111101010100000",
703 => "000000110001111110000011",
704 => "000000110100011011111110",
705 => "000001000110101011110111",
706 => "000001001100110111101111",
707 => "000001001000001001101111",
708 => "000001010001010000110101",
709 => "000001011100101001110011",
710 => "000001011010011001001001",
711 => "000001010111011100110110",
712 => "000001011111001010111101",
713 => "000001101010100001100110",
714 => "000001111000110111110000",
715 => "000010001101110101110110",
716 => "000010010110011111100110",
717 => "000010000010100110101110",
718 => "000001101001001101110111",
719 => "000001101010000000111001",
720 => "000001110100100001100111",
721 => "000001110110010001011010",
722 => "000010000100000001110000",
723 => "000010001001001010111100",
724 => "000001111011011010100010",
725 => "000010000110000100011110",
726 => "000010000111111011100011",
727 => "000001110010111101000010",
728 => "000010001001010011010000",
729 => "000010011110111011001100",
730 => "000010000010001000011011",
731 => "000001110111001001010000",
732 => "000010000001110010110010",
733 => "000001101110110101010111",
734 => "000001010000100001110000",
735 => "000001001101001100001000",
736 => "000001110001101001110101",
737 => "000010101100100110100110",
738 => "000011001011100010001011",
739 => "000010110010100000001010",
740 => "000010001100001010011111",
741 => "000010000101110010000101",
742 => "000010001111101101111010",
743 => "000010001110001010010111",
744 => "000010000001111001100010",
745 => "000010000001010111010100",
746 => "000010001100100010110000",
747 => "000001111100100011111000",
748 => "000001011001000101111011",
749 => "000001011000100111111100",
750 => "000001101101111101000011",
751 => "000001101110000111100110",
752 => "000001110101101011100011",
753 => "000010001111000100011100",
754 => "000010010011100011101110",
755 => "000010001010111001000011",
756 => "000001111101111111101100",
757 => "000001101101011001101011",
758 => "000001110000110011111110",
759 => "000001111101010011011011",
760 => "000001111110011111001110",
761 => "000001111000010100000101",
762 => "000001101111001011100110",
763 => "000001011001011011010001",
764 => "000000111000001000000000",
765 => "000000100101011101110001",
766 => "000000100010011111011010",
767 => "000000101100001100001001",
768 => "000000111111101111011010",
769 => "000001001000001110101100",
770 => "000001001001001110010110",
771 => "000001000110100011010110",
772 => "000001000100111001100010",
773 => "000000111111110100010110",
774 => "000000100110100110010110",
775 => "000000010000001110001110",
776 => "000000000100111110011110",
777 => "111111111101011111100001",
778 => "111111111111001110100110",
779 => "000000000010101011110000",
780 => "000000000011001010101111",
781 => "111111111001000111010111",
782 => "111111101101010001010011",
783 => "111111100110111010001000",
784 => "111111010111001010111010",
785 => "111111001000001101100001",
786 => "111111000001010100110010",
787 => "111110111001010111110110",
788 => "111110110000000111111010",
789 => "111110101100000110100111",
790 => "111110101000000100010100",
791 => "111110011101101011100001",
792 => "111110100100100111110101",
793 => "111110110011110010011100",
794 => "111110110100101001000111",
795 => "111110110110100111011100",
796 => "111110101100110001000110",
797 => "111110010111110101100110",
798 => "111110010001010000000000",
799 => "111110000110001100000011",
800 => "111101101010100000010011",
801 => "111101010010100111110001",
802 => "111101001111110000110011",
803 => "111101011110100101000000",
804 => "111101101010101100001001",
805 => "111101101010010110001101",
806 => "111101100111111001001001",
807 => "111101101011100001111100",
808 => "111101101100010111101110",
809 => "111101101100111100101011",
810 => "111101111001111011101011",
811 => "111110000110110111010010",
812 => "111110000111110100011011",
813 => "111110000000100111111111",
814 => "111101110101010100110001",
815 => "111101110010101010100110",
816 => "111101111000001001110101",
817 => "111101110001110011000001",
818 => "111101100101101010010011",
819 => "111101101001100111111011",
820 => "111101110101111011100001",
821 => "111101110100101101100110",
822 => "111101101101111001111010",
823 => "111101110000101111101000",
824 => "111101101101000011100001",
825 => "111101101001000111000011",
826 => "111101111011100110001010",
827 => "111110001001011011100110",
828 => "111110000110011011101001",
829 => "111110000011111000010101",
830 => "111101111110111100001110",
831 => "111110000000011111101111",
832 => "111110001010010100011101",
833 => "111110010111010100100100",
834 => "111110101100101100010000",
835 => "111110110010000111110000",
836 => "111110101011111110010111",
837 => "111110111010001010110010",
838 => "111111000010001001101110",
839 => "111110110001111101001110",
840 => "111110100011110110001101",
841 => "111110011101101000000010",
842 => "111110011110001101001100",
843 => "111110101000001011010110",
844 => "111110101010110001101101",
845 => "111110011101001001000010",
846 => "111110010110110111111101",
847 => "111110101100011111001011",
848 => "111111001011110110101010",
849 => "111111011100010100110111",
850 => "111111011110110101001110",
851 => "111111100000001101011011",
852 => "111111100110000010110011",
853 => "111111011110010010010010",
854 => "111111001000000101111110",
855 => "111111000110011110100101",
856 => "111111001111000100101101",
857 => "111110111111101100110000",
858 => "111110101100011010111010",
859 => "111110101111011111011100",
860 => "111110111101101110010010",
861 => "111111000001001010001010",
862 => "111110111101001111111100",
863 => "111111001001100101000010",
864 => "111111100010110011100011",
865 => "111111110011110010001011",
866 => "111111111001011110001011",
867 => "111111111011110111100000",
868 => "111111111101101101010000",
869 => "111111111000001010001101",
870 => "111111101110011011001110",
871 => "111111110000010101101000",
872 => "111111111100101011000011",
873 => "000000000100101000001110",
874 => "111111111100110011001110",
875 => "111111101011100000110110",
876 => "111111101011011110001011",
877 => "111111111011001010110011",
878 => "111111111111100110101010",
879 => "111111111011101100001000",
880 => "000000000110010001001110",
881 => "000000100000001011010101",
882 => "000000101000010001101001",
883 => "000000011001000001101101",
884 => "000000011010010011111001",
885 => "000000101010010110100110",
886 => "000000101111110000101110",
887 => "000000110001101000100100",
888 => "000000110010111011011011",
889 => "000000110100111100101011",
890 => "000001000110101000000111",
891 => "000001010110110010011001",
892 => "000001001111110110010001",
893 => "000001001111001101010010",
894 => "000001010100000001011111",
895 => "000001001011110010001000",
896 => "000001000111011110110010",
897 => "000000111000001011011111",
898 => "000000110101010110000110",
899 => "000001001011001000000001",
900 => "000000111010011101111001",
901 => "000000110100101101110101",
902 => "000001101000110010110010",
903 => "000010001101000101100110",
904 => "000010010000011011000111",
905 => "000010010010101111111000",
906 => "000010010110100101000101",
907 => "000010010100000001010111",
908 => "000010010001001001000100",
909 => "000010001000000100100011",
910 => "000001111001000000001010",
911 => "000001111100110101011000",
912 => "000001111011110011010101",
913 => "000001111011011100100100",
914 => "000010010000001010010110",
915 => "000010001000100110101001",
916 => "000001111001101001101111",
917 => "000010000110000100110100",
918 => "000010000010001111111001",
919 => "000001111010010111100110",
920 => "000010010101111101101011",
921 => "000010011100111001111001",
922 => "000001110001101100100111",
923 => "000001100111000001011110",
924 => "000001101101011101111111",
925 => "000001010110000111011011",
926 => "000001111000110011011000",
927 => "000011000001110101001111",
928 => "000011000001110111001110",
929 => "000010010001101111000110",
930 => "000001111001110010100110",
931 => "000010001000010100111100",
932 => "000010011100010001010100",
933 => "000010010000011010100111",
934 => "000001110111001010100010",
935 => "000001111100001101110101",
936 => "000010000100011111100110",
937 => "000001101110111111100110",
938 => "000001101010100011101111",
939 => "000001110000111110111011",
940 => "000001011000000000010000",
941 => "000001001101111010010011",
942 => "000001101101010110111110",
943 => "000010001101011100101010",
944 => "000010011100001110010001",
945 => "000010011110010100100000",
946 => "000010010011010011100101",
947 => "000010001010111110001010",
948 => "000010001101101011001010",
949 => "000010001000011001011001",
950 => "000001111111010110110101",
951 => "000001110010000111011110",
952 => "000001010010010011101110",
953 => "000000111100010011110111",
954 => "000000110100011110010111",
955 => "000000100100101001001011",
956 => "000000100111000111011011",
957 => "000001000000100111110010",
958 => "000001001010101001000001",
959 => "000001000111110110100100",
960 => "000001010010000011011000",
961 => "000001011000011000010100",
962 => "000001000110011100010000",
963 => "000000101101100010110100",
964 => "000000010001110001010010",
965 => "111111110101001010010000",
966 => "111111101011110011011100",
967 => "111111110010000011011010",
968 => "000000000011011001101011",
969 => "000000001101011111001100",
970 => "111111111100001111010000",
971 => "111111110011111001111101",
972 => "111111111010011110001101",
973 => "111111101111111101110111",
974 => "111111011011111010010001",
975 => "111111001001101101101001",
976 => "111110110111001111111111",
977 => "111110100110111111100000",
978 => "111110011101111100110100",
979 => "111110010010111000101001",
980 => "111110001001011011001011",
981 => "111110011001010000100000",
982 => "111110101010001100110110",
983 => "111110101110111110011100",
984 => "111110111111110000001010",
985 => "111111000100100100101001",
986 => "111110110011100110010000",
987 => "111110101000010000011001",
988 => "111110011010011110010001",
989 => "111110000110011011110001",
990 => "111101111111110000010000",
991 => "111110000000001000010001",
992 => "111101111101110111101101",
993 => "111110000000001110010011",
994 => "111101111100001000011010",
995 => "111101101110011000111101",
996 => "111101101011100101011110",
997 => "111101101111111010010101",
998 => "111101110011001000001111",
999 => "111101111100010100010011",
1000 => "111110000011010111011001",
1001 => "111110000101101000100010",
1002 => "111110001101000001011000",
1003 => "111110010110011001111000",
1004 => "111110011101000111000000",
1005 => "111110011011110001101111",
1006 => "111110010001111100000000",
1007 => "111110010000001001100001",
1008 => "111110011001000011000011",
1009 => "111110011011111110101100",
1010 => "111110010010001101111011",
1011 => "111110001001000110000001",
1012 => "111110000110000111001010",
1013 => "111101111100010101101100",
1014 => "111101111001100010011000",
1015 => "111110001010101011110110",
1016 => "111110010110101101101011",
1017 => "111110010100100001100100",
1018 => "111110001011101110011011",
1019 => "111110000000101000010111",
1020 => "111110000101110001001101",
1021 => "111110011001110111100010",
1022 => "111110011011010000001110",
1023 => "111110001111001000000101",
1024 => "111110100000100000111010",
1025 => "111111000100101000100010",
1026 => "111111010001111010010101",
1027 => "111111001100000100011010",
1028 => "111111000010011001000010",
1029 => "111110111000010111010011",
1030 => "111110101110110111000101",
1031 => "111110011011001011111100",
1032 => "111110001101110100110101",
1033 => "111110011011001001111110",
1034 => "111110100000100011111101",
1035 => "111110001011010011101010",
1036 => "111101111110100010110010",
1037 => "111110010111111100001010",
1038 => "111110111110110010101010",
1039 => "111111000000010111100011",
1040 => "111110110101101110110011",
1041 => "111111010001101111000011",
1042 => "111111110100111010100011",
1043 => "111111101101000001101010",
1044 => "111111000101000011010000",
1045 => "111110110000011011101000",
1046 => "111110111011000010000100",
1047 => "111111000000100101001010",
1048 => "111110110000010000100001",
1049 => "111110101000110010001010",
1050 => "111111000100100111111011",
1051 => "111111010011000000011001",
1052 => "111110110101101010011110",
1053 => "111110100101011001101111",
1054 => "111111000010100001000001",
1055 => "111111101001110010001100",
1056 => "111111101100011001000110",
1057 => "111111011101110010011010",
1058 => "111111101110101101000101",
1059 => "000000000101001101000001",
1060 => "111111111000111101101111",
1061 => "111111011100011100111010",
1062 => "111111010110101111001010",
1063 => "111111101001000110100101",
1064 => "111111101100000001111101",
1065 => "111111010011100110010011",
1066 => "111111001010111110101110",
1067 => "111111100001010110001000",
1068 => "111111100101011100111000",
1069 => "111111001111010010010000",
1070 => "111111001111111111101101",
1071 => "111111110010011101000110",
1072 => "000000001101111010001101",
1073 => "000000001001101101110100",
1074 => "000000000011001000000000",
1075 => "000000001011011110100100",
1076 => "000000010001011111111011",
1077 => "000000001000111011100100",
1078 => "111111111100001010001101",
1079 => "000000001001111110101110",
1080 => "000000101001001001011111",
1081 => "000000110001001000011110",
1082 => "000000011100111010100011",
1083 => "000000011001011100100100",
1084 => "000000110111110011000110",
1085 => "000000110101111000001110",
1086 => "000000010100101010100001",
1087 => "000000011000111110010111",
1088 => "000000100101001100000011",
1089 => "000000010001011100010110",
1090 => "000000010011010111001100",
1091 => "000000110010011110000010",
1092 => "000000110100011001000011",
1093 => "000000111011001110100010",
1094 => "000001011100111000001110",
1095 => "000001101001100100111111",
1096 => "000001110111111000010101",
1097 => "000010001011101011000110",
1098 => "000010000000100010001110",
1099 => "000001011010111010001101",
1100 => "000001001010000010000100",
1101 => "000001101001101001000011",
1102 => "000001101100010011101110",
1103 => "000001001101000100111010",
1104 => "000001011011100000000001",
1105 => "000001101001000011000000",
1106 => "000001000111101010101110",
1107 => "000001001000111001110010",
1108 => "000010000110010011110101",
1109 => "000010001110101011011000",
1110 => "000001100101101010101100",
1111 => "000001011111010010000110",
1112 => "000000111011001111011001",
1113 => "000000010110111101110001",
1114 => "000001100010111011000010",
1115 => "000010111110010110111010",
1116 => "000010111011110111000011",
1117 => "000010100111001001100010",
1118 => "000010110101011000001001",
1119 => "000010101110010001000110",
1120 => "000010100011111110001011",
1121 => "000010110111010111100111",
1122 => "000010101111101010101010",
1123 => "000010001100010101000101",
1124 => "000001111000000001110111",
1125 => "000001110100100011011111",
1126 => "000001101010001111010010",
1127 => "000001001100000000000000",
1128 => "000001000000111010010011",
1129 => "000001010110101011010111",
1130 => "000001101010111110000010",
1131 => "000010000001100100010100",
1132 => "000010011101111100111111",
1133 => "000010011110001101000001",
1134 => "000010000100000010111001",
1135 => "000001110000100011101011",
1136 => "000001101110000000111011",
1137 => "000010000010010100001100",
1138 => "000010011110011101110001",
1139 => "000010010000000101101011",
1140 => "000001100100101110010110",
1141 => "000001011010000100011100",
1142 => "000001001101110101001000",
1143 => "000000100100010111000110",
1144 => "000000100000010000101110",
1145 => "000000110100100111000011",
1146 => "000000101101010010100000",
1147 => "000000101000111110011010",
1148 => "000000111110110001000110",
1149 => "000001001100110000001100",
1150 => "000001000011011010001000",
1151 => "000001000100101100111000",
1152 => "000000111011111001111011",
1153 => "000000010010011000101001",
1154 => "111111111101010001110011",
1155 => "000000000001000001001101",
1156 => "000000000011010111111100",
1157 => "111111111101000001100110",
1158 => "111111110110101110111010",
1159 => "111111111001111110110110",
1160 => "111111110001100001100110",
1161 => "111111110100010010101110",
1162 => "000000000101010110111010",
1163 => "111111111011001001001101",
1164 => "111111100010001000001100",
1165 => "111111001001110100110100",
1166 => "111110110010011100100011",
1167 => "111110011101101100100101",
1168 => "111110011000111011011110",
1169 => "111110100101110001011011",
1170 => "111110101101101011000001",
1171 => "111110111101001110001101",
1172 => "111111001101111000101000",
1173 => "111111010011101101110101",
1174 => "111111100000111110100010",
1175 => "111111100011011011010101",
1176 => "111111010001111111001001",
1177 => "111111000001111010100001",
1178 => "111110111001011111110010",
1179 => "111110101010100110001110",
1180 => "111110011010100110001110",
1181 => "111110100001111110000100",
1182 => "111110100011111010010101",
1183 => "111110010011001011111000",
1184 => "111110010100110011010011",
1185 => "111110011101111010010110",
1186 => "111110011010111011101001",
1187 => "111110010110010000011000",
1188 => "111110010011010100010110",
1189 => "111110010111101111010111",
1190 => "111110100111010101001011",
1191 => "111110111010110111100010",
1192 => "111111000111101011101001",
1193 => "111111001100100001111011",
1194 => "111111000110010101000001",
1195 => "111110101110110110100001",
1196 => "111110100100110110011001",
1197 => "111110101011000110111000",
1198 => "111110100010111101101100",
1199 => "111110011101001011110000",
1200 => "111110010110110110011010",
1201 => "111110010100110101000010",
1202 => "111110101010111001011010",
1203 => "111110101100011110011001",
1204 => "111110100000011000010000",
1205 => "111110101000110111010011",
1206 => "111110101001111100110110",
1207 => "111110011101100000110101",
1208 => "111110011100001100101100",
1209 => "111110110011110111101010",
1210 => "111111001100101110001000",
1211 => "111111001001011001100100",
1212 => "111110111000110101001101",
1213 => "111110111001101010000011",
1214 => "111111010100000100010110",
1215 => "111111110101101110001001",
1216 => "000000001010000110000101",
1217 => "111111110100000010100000",
1218 => "111111000100000000011100",
1219 => "111110101010101101000000",
1220 => "111110010010011101110110",
1221 => "111110000000111100011010",
1222 => "111110001101101010010011",
1223 => "111110010011010010011000",
1224 => "111110010010011101110011",
1225 => "111110011001111010100111",
1226 => "111110101011001011010010",
1227 => "111111001011110010111000",
1228 => "111111011010011100101001",
1229 => "111111010000001000111110",
1230 => "111111010001010001111110",
1231 => "111111011011111000101011",
1232 => "111111100011011010000110",
1233 => "111111101010100011011011",
1234 => "111111011111101111001101",
1235 => "111111000010110101111001",
1236 => "111110100111111000010100",
1237 => "111110011001001100011100",
1238 => "111110100110001110001111",
1239 => "111110110110100101110110",
1240 => "111110101011110110110011",
1241 => "111110100110011000101100",
1242 => "111110110010100101011111",
1243 => "111110111010000000100110",
1244 => "111111000001000101100010",
1245 => "111111001101000011001100",
1246 => "111111011111011100000001",
1247 => "111111111011000010101000",
1248 => "000000001010000101010100",
1249 => "000000000110101101101100",
1250 => "000000000100010010010011",
1251 => "111111111011001110001110",
1252 => "111111010101011101010100",
1253 => "111110101000100010011111",
1254 => "111110101011001111101110",
1255 => "111111001101110101011101",
1256 => "111111010101101110101011",
1257 => "111111001001110000010111",
1258 => "111111001011000110000001",
1259 => "111111100100001000000110",
1260 => "111111111111001110010001",
1261 => "000000000100001001110000",
1262 => "111111111101001111110001",
1263 => "000000000001101010011101",
1264 => "000000010010000000000010",
1265 => "000000000111101010000000",
1266 => "111111101101000000010011",
1267 => "111111110010010101110011",
1268 => "000000000000011000010110",
1269 => "000000000000101001010001",
1270 => "000000010011000011011001",
1271 => "000000110011000001000100",
1272 => "000000100011101110100100",
1273 => "000000000100110100011100",
1274 => "000000010010110111111110",
1275 => "000000000101000110001011",
1276 => "111111100001010100001111",
1277 => "111111110110100011110101",
1278 => "000000001110010110100010",
1279 => "000000000101011000011110",
1280 => "000000010100110001000010",
1281 => "000000111011101010011001",
1282 => "000001001011001100001101",
1283 => "000001100100110111010100",
1284 => "000010001100011101100000",
1285 => "000010000010110011011010",
1286 => "000001111000110010010111",
1287 => "000010000101110010111011",
1288 => "000001100000011111000110",
1289 => "000000110000100101001110",
1290 => "000000111111100101000010",
1291 => "000001001011100100101010",
1292 => "000000110101101110111011",
1293 => "000001010100000111000110",
1294 => "000001110101110100111010",
1295 => "000001010011000000110110",
1296 => "000001000000010110101111",
1297 => "000001001000010100010110",
1298 => "000000110000110010001010",
1299 => "000000011000010110011110",
1300 => "000001000011000011101000",
1301 => "000010011111111000100011",
1302 => "000011001110111001011010",
1303 => "000010111011110100001010",
1304 => "000010011111000001110111",
1305 => "000010010110000110011100",
1306 => "000010001110111111110000",
1307 => "000010001101000110101001",
1308 => "000010010011110100110011",
1309 => "000010000000011011101001",
1310 => "000001111011101001110100",
1311 => "000010001000111011011111",
1312 => "000001100110010111001011",
1313 => "000001000011100001011101",
1314 => "000001001011010111000010",
1315 => "000001011010001010010011",
1316 => "000001100011110010000110",
1317 => "000001111110001011010010",
1318 => "000010011001111001111000",
1319 => "000010001001001001011100",
1320 => "000001110000011111011010",
1321 => "000001110000010001010100",
1322 => "000001111000110011011101",
1323 => "000010011111000010011001",
1324 => "000011000110010001001000",
1325 => "000011000000000000010010",
1326 => "000010100110000110100011",
1327 => "000010001111001010110000",
1328 => "000001110001110100010001",
1329 => "000001000000110011010100",
1330 => "000000010110111010110010",
1331 => "000000011011100100110000",
1332 => "000000101101000011111010",
1333 => "000000110111011101001010",
1334 => "000001001111100110101111",
1335 => "000001011111110000010100",
1336 => "000001100111011000011010",
1337 => "000001110001001100100010",
1338 => "000001100101010111000101",
1339 => "000001000001101010100000",
1340 => "000000101010010111101100",
1341 => "000000110111011111111110",
1342 => "000000111100011001000101",
1343 => "000000110001010111101101",
1344 => "000000111000000100000011",
1345 => "000000110001010000100100",
1346 => "000000100100001101111101",
1347 => "000000101101000000010110",
1348 => "000000110011000011111101",
1349 => "000000100101110101001001",
1350 => "000000010001111100100111",
1351 => "000000000111111101100000",
1352 => "111111110011100000010000",
1353 => "111111011110111011110101",
1354 => "111111011111001101010110",
1355 => "111111011010000011000110",
1356 => "111111100010101000010100",
1357 => "000000000101010100000100",
1358 => "000000100000110000010010",
1359 => "000000101010101100111110",
1360 => "000000101111111000010100",
1361 => "000000110011001110001011",
1362 => "000000011111001010101011",
1363 => "111111111011010000110100",
1364 => "111111011001001010000011",
1365 => "111110111010101100100010",
1366 => "111110101001110000001010",
1367 => "111110100011100010010000",
1368 => "111110110010010101000000",
1369 => "111111010000101111011001",
1370 => "111111011100010010100011",
1371 => "111111010101110110011011",
1372 => "111111000101000111110001",
1373 => "111110110010011011001101",
1374 => "111110101110111000000010",
1375 => "111110100110010110001000",
1376 => "111110011011001000001100",
1377 => "111110111001101101001110",
1378 => "111111100111101111011101",
1379 => "111111110101001111110110",
1380 => "111111100110110011100111",
1381 => "111111001100000100001001",
1382 => "111111000010010010101111",
1383 => "111111000100100001001111",
1384 => "111110111100000011001110",
1385 => "111110101101011100000100",
1386 => "111110011101001101110100",
1387 => "111110011111000000100010",
1388 => "111110011011110101011000",
1389 => "111110000101010000000110",
1390 => "111110000001001100100001",
1391 => "111110000100111010110101",
1392 => "111110010010001010100111",
1393 => "111110101110110110010111",
1394 => "111111000000011110011000",
1395 => "111111000011001010111101",
1396 => "111110110100111011001100",
1397 => "111110100111111010100101",
1398 => "111110100100010111011110",
1399 => "111110100101101010100010",
1400 => "111110111000011101000011",
1401 => "111111000000100011110001",
1402 => "111110110110010001000011",
1403 => "111110111000101111100100",
1404 => "111110111001101100110010",
1405 => "111110011100000111110110",
1406 => "111101101001111010010000",
1407 => "111101001000111010001011",
1408 => "111101000000011000110101",
1409 => "111101000000001110000110",
1410 => "111101011001111100110110",
1411 => "111110001100010110001011",
1412 => "111110101011000010010011",
1413 => "111110100100111000110101",
1414 => "111110010111011010100000",
1415 => "111110100110010110111101",
1416 => "111111000001111100100100",
1417 => "111111001101001001100100",
1418 => "111111011001000000000100",
1419 => "111111011000011000001011",
1420 => "111110101111001111011010",
1421 => "111101111101111110100101",
1422 => "111101100001011110111000",
1423 => "111101010010111000010101",
1424 => "111101000111001011100101",
1425 => "111101000000111101011110",
1426 => "111101010001000101110000",
1427 => "111101110100101011110011",
1428 => "111110001110011011101000",
1429 => "111110010001100000101111",
1430 => "111110001100001010000111",
1431 => "111110010010100101100101",
1432 => "111110110011001111011000",
1433 => "111111010001100010101111",
1434 => "111111010000101111110101",
1435 => "111111001101111101110110",
1436 => "111111001111001011011000",
1437 => "111111000010101010110000",
1438 => "111110101010101111011011",
1439 => "111110001111101101001011",
1440 => "111110001111101011000001",
1441 => "111110100011000001011001",
1442 => "111110011001100011101100",
1443 => "111101111100110010011010",
1444 => "111101111100000000111000",
1445 => "111110011101000110010111",
1446 => "111110110010001100000111",
1447 => "111110101010000101000100",
1448 => "111110110010001110110001",
1449 => "111111010001101001010111",
1450 => "111111011101011010011001",
1451 => "111111010010011100010001",
1452 => "111111010010110011011101",
1453 => "111111111010011001000011",
1454 => "000000100100001111100110",
1455 => "000000011000100010000101",
1456 => "000000001010010110110000",
1457 => "000000010100001100110101",
1458 => "111111111100111001000111",
1459 => "111111100000100111110010",
1460 => "111111101111111101111001",
1461 => "111111110101111010010111",
1462 => "111111010010111101110111",
1463 => "111111100111110100101000",
1464 => "000000101000001011011010",
1465 => "000000001010011011101111",
1466 => "111111111001001101100111",
1467 => "000001001010100111100010",
1468 => "000001011111111000010001",
1469 => "000001000101100111010111",
1470 => "000001010110101000001111",
1471 => "000001101110010010001000",
1472 => "000010010000101011010011",
1473 => "000010100001101011001111",
1474 => "000001110101010000100011",
1475 => "000001011010111001100011",
1476 => "000001101110001000101111",
1477 => "000001110001010101000111",
1478 => "000001101011100110011000",
1479 => "000001011010111101001101",
1480 => "000000111010100110010100",
1481 => "000000101101101100010111",
1482 => "000000000100110011010011",
1483 => "111111000101111111010001",
1484 => "111111110100001011110110",
1485 => "000010010100011100000011",
1486 => "000100010000010100011110",
1487 => "000100010101110101010100",
1488 => "000011101000100001010100",
1489 => "000011010101001110101100",
1490 => "000011100000000011000001",
1491 => "000011011000001110111111",
1492 => "000010100010100100110010",
1493 => "000010010011010010101000",
1494 => "000010111001010001011101",
1495 => "000010011111110001011100",
1496 => "000001100011111011111001",
1497 => "000001011001111010111001",
1498 => "000001001111010100010110",
1499 => "000001010001010010111101",
1500 => "000010000010110110011010",
1501 => "000010100001111101111110",
1502 => "000010111010101111111110",
1503 => "000011011100101010001111",
1504 => "000011001101111101100001",
1505 => "000010101000100110001000",
1506 => "000010010011110011111110",
1507 => "000010010110001101001100",
1508 => "000010111001010111111111",
1509 => "000011010001100001101110",
1510 => "000011001000000001101010",
1511 => "000010111111111100100000",
1512 => "000010110010100000101001",
1513 => "000010001011011100000011",
1514 => "000001110000010101111000",
1515 => "000001110000010001100000",
1516 => "000001101000011100100010",
1517 => "000001011000110001101100",
1518 => "000001010011110111101001",
1519 => "000001011000110111100100",
1520 => "000001100101110101001000",
1521 => "000001111000011111000100",
1522 => "000001111011111010110100",
1523 => "000001100010111010010001",
1524 => "000001001101100001110110",
1525 => "000001001110000101001111",
1526 => "000001010110000011000110",
1527 => "000001100001001100010101",
1528 => "000001100101011001101100",
1529 => "000001100011111010111110",
1530 => "000001101111011110000010",
1531 => "000001110010101111100000",
1532 => "000001011100000010100001",
1533 => "000001010000000000001011",
1534 => "000001000110011101111000",
1535 => "000000011101011000011011",
1536 => "111111111010101010110001",
1537 => "111111101111011000111000",
1538 => "111111100101110101011110",
1539 => "111111101010110001110100",
1540 => "111111111011101010101011",
1541 => "000000000010110100100011",
1542 => "000000010010000100001011",
1543 => "000000100101111010011011",
1544 => "000000010111011001001000",
1545 => "000000010100110111110010",
1546 => "000000110000010100000111",
1547 => "000000100001000010000110",
1548 => "000000000001001001110101",
1549 => "111111101110011100101110",
1550 => "111111010101110100100000",
1551 => "111111001001100010110010",
1552 => "111110110101100110010101",
1553 => "111110101000011101101101",
1554 => "111111000101110011010010",
1555 => "111111011100110010001100",
1556 => "111111001101001110000110",
1557 => "111110110110001010111000",
1558 => "111110110111101101011011",
1559 => "111111000000001110110010",
1560 => "111111000100101011100000",
1561 => "111111011101101111011001",
1562 => "111111111110110001111000",
1563 => "000000010001011001111101",
1564 => "000000000011101101110011",
1565 => "111111010100001111000111",
1566 => "111110110100110100000001",
1567 => "111110110111000110101000",
1568 => "111110110011001100101100",
1569 => "111110010111110111110101",
1570 => "111110001001110011010010",
1571 => "111110011101111110000010",
1572 => "111110101000001011011000",
1573 => "111110010101000101100100",
1574 => "111110000111110001000010",
1575 => "111110001011100100011010",
1576 => "111110010100010101000111",
1577 => "111110001101011000011001",
1578 => "111101101100111110101001",
1579 => "111101100101011001101011",
1580 => "111110010000011111001110",
1581 => "111110110001101000110101",
1582 => "111110101011011100010001",
1583 => "111110011110011011100110",
1584 => "111110100101010011100111",
1585 => "111111000110111101101010",
1586 => "111111011110101011000010",
1587 => "111111000010111010100101",
1588 => "111110010111011010001110",
1589 => "111101111001101000100010",
1590 => "111101001000110101001100",
1591 => "111100001111111101110111",
1592 => "111011110110000101000000",
1593 => "111100000110011010111011",
1594 => "111101000100010001010000",
1595 => "111110000011010111111001",
1596 => "111110010100111010111101",
1597 => "111110010001010101100001",
1598 => "111110011000101001110000",
1599 => "111110100000010011001111",
1600 => "111110010001000110110011",
1601 => "111110000001001011100010",
1602 => "111110010011011010001010",
1603 => "111110101011010011111100",
1604 => "111110100110011111010111",
1605 => "111110001000110110100111",
1606 => "111101100000010101110100",
1607 => "111101000101111111011011",
1608 => "111100111101000101101000",
1609 => "111100101110011111011110",
1610 => "111100100011001100100111",
1611 => "111100110110001110000011",
1612 => "111101011010110000011111",
1613 => "111101101011011101100101",
1614 => "111101100110011111101000",
1615 => "111101101100010011101101",
1616 => "111110001001101010111010",
1617 => "111110011110110010001100",
1618 => "111110010001111101000101",
1619 => "111110001111001011101100",
1620 => "111110110010001010111000",
1621 => "111111000111010111011100",
1622 => "111110110111110011110100",
1623 => "111110011000011110001110",
1624 => "111110001000111110010011",
1625 => "111110011001000101101100",
1626 => "111110010000100011110000",
1627 => "111101011111101010110101",
1628 => "111101001110000101110001",
1629 => "111101110100010000001000",
1630 => "111110100011100111111101",
1631 => "111110101010010100101011",
1632 => "111110011010100110111011",
1633 => "111110101100100011000100",
1634 => "111111010111111110011100",
1635 => "111111101100000010001100",
1636 => "111111100100101111010010",
1637 => "111111101110000000010011",
1638 => "000000000010100000001011",
1639 => "111111110111100001000000",
1640 => "111111100001011100011011",
1641 => "111111010111100100001101",
1642 => "111111010111011110010000",
1643 => "111111101010110110001101",
1644 => "000000000010101111110011",
1645 => "000000000001101101000101",
1646 => "111111100101111111110010",
1647 => "111111100001101110011001",
1648 => "000000000111001011001111",
1649 => "000000010001000000101001",
1650 => "000000000110011010111111",
1651 => "000000100000011010010101",
1652 => "000001000100011111100111",
1653 => "000001011110000001110000",
1654 => "000001011011100001010110",
1655 => "000001010011010110000000",
1656 => "000010001100010101111000",
1657 => "000010101101111100110101",
1658 => "000010000011001010101001",
1659 => "000010001110110000110110",
1660 => "000010100101111110010000",
1661 => "000001100111110110001101",
1662 => "000000111100110000010001",
1663 => "000000100111111001001101",
1664 => "111111010101111100101010",
1665 => "111110011101010000010101",
1666 => "111111001111110111001111",
1667 => "000001010001101110001000",
1668 => "000011100101000101111010",
1669 => "000100100101111100110111",
1670 => "000100000011111011100100",
1671 => "000011101010011110010000",
1672 => "000011111001010001001100",
1673 => "000011110101000100000101",
1674 => "000011101010111111011001",
1675 => "000011110110001100101100",
1676 => "000011100000000010001110",
1677 => "000010110000000101101100",
1678 => "000010010111000011011101",
1679 => "000001101010011010001101",
1680 => "000000110110010010011110",
1681 => "000000111000110010010011",
1682 => "000001011111011101110001",
1683 => "000010100001101011011100",
1684 => "000011101000110101000011",
1685 => "000100000010011101011001",
1686 => "000100000011111110010111",
1687 => "000011110011100100110100",
1688 => "000011010010000010111001",
1689 => "000011011111110111011111",
1690 => "000100000011001111000100",
1691 => "000011101110101100000110",
1692 => "000011010110000010110011",
1693 => "000011011101010101001000",
1694 => "000010110100110110001000",
1695 => "000001101010001111011011",
1696 => "000001011001010100111100",
1697 => "000001101011011110101001",
1698 => "000001111010011111010010",
1699 => "000010011001000000001001",
1700 => "000010110110010100100110",
1701 => "000011001111000101111010",
1702 => "000011100000001111010101",
1703 => "000010111001100101001011",
1704 => "000001110000101111111001",
1705 => "000001000001101000010100",
1706 => "000000101101000000000111",
1707 => "000000110001101110010001",
1708 => "000001010001011000110101",
1709 => "000001110001101110110011",
1710 => "000001111110110101111001",
1711 => "000001111111100101011100",
1712 => "000010001000001111010110",
1713 => "000010010011101000110010",
1714 => "000010001011001101000001",
1715 => "000001110101101010011101",
1716 => "000001011101111011100111",
1717 => "000000111000001110011111",
1718 => "000000000011001110101110",
1719 => "111111010100001110010111",
1720 => "111110111000001010101010",
1721 => "111110100010110100100011",
1722 => "111110010010010001110010",
1723 => "111110011010011110000001",
1724 => "111110110111101110101111",
1725 => "111111011101011000100110",
1726 => "000000010011101011111000",
1727 => "000001000100110101010110",
1728 => "000001000110100110011111",
1729 => "000000100011101011110101",
1730 => "000000000000011000101011",
1731 => "111111110010011000111100",
1732 => "000000000000101100001100",
1733 => "111111111110100011010110",
1734 => "111111001011000100000100",
1735 => "111110011111101001010100",
1736 => "111110010000111101101011",
1737 => "111101110100101110010101",
1738 => "111101100011111110110001",
1739 => "111101111001000010010100",
1740 => "111110010011010000100101",
1741 => "111110100110101100000000",
1742 => "111110110111000011011100",
1743 => "111111010001010111111100",
1744 => "111111110111011011011110",
1745 => "111111110110111010100101",
1746 => "111111000010111111101000",
1747 => "111110001001101011010011",
1748 => "111101100110100111010001",
1749 => "111101100001001010000000",
1750 => "111101110000111010100111",
1751 => "111110000101001111101001",
1752 => "111110001100110111111001",
1753 => "111110000000000101110011",
1754 => "111101111100110000101001",
1755 => "111110010010000111101000",
1756 => "111110101011110011010110",
1757 => "111110111001101110110100",
1758 => "111110011011101000010100",
1759 => "111101001110010001111101",
1760 => "111100010111100010001100",
1761 => "111100011010011111110010",
1762 => "111100101101010111001001",
1763 => "111100110100101101000111",
1764 => "111100111011111111101110",
1765 => "111101010110101111000101",
1766 => "111110010100111100010110",
1767 => "111111010101011100011010",
1768 => "111111011111011101100100",
1769 => "111110111000000100101100",
1770 => "111101110000111000100111",
1771 => "111100011100000011100011",
1772 => "111011110010110100000001",
1773 => "111011111100011110110101",
1774 => "111100010101101010001010",
1775 => "111100100010101101111000",
1776 => "111100000101110001110111",
1777 => "111011110000111000011110",
1778 => "111100011110010000100101",
1779 => "111101010100011101101100",
1780 => "111101110000000111110011",
1781 => "111110010001010100010101",
1782 => "111110101111001100100010",
1783 => "111110100111101101011111",
1784 => "111110000010011011000011",
1785 => "111101110010011000101101",
1786 => "111101110101011000110111",
1787 => "111101001000001001101111",
1788 => "111100000001111100110110",
1789 => "111011111110101010000011",
1790 => "111100111101110110011100",
1791 => "111101110100101110001110",
1792 => "111101110001011000010111",
1793 => "111101001011000001011100",
1794 => "111101000100001101111001",
1795 => "111101101001100011001101",
1796 => "111110001000010111000100",
1797 => "111110000100011111110010",
1798 => "111110000001100000111011",
1799 => "111110011101001110111101",
1800 => "111110101001101110100000",
1801 => "111110010101011011110110",
1802 => "111110011101001000000011",
1803 => "111111000010001000000001",
1804 => "111111001101001101011100",
1805 => "111110101101111101001110",
1806 => "111110001001001011001111",
1807 => "111110011010011110010110",
1808 => "111111000111000001000100",
1809 => "111111000011000101100011",
1810 => "111110100101011011100101",
1811 => "111110101010010100111010",
1812 => "111111010100111101001100",
1813 => "111111110000010100111111",
1814 => "111111100001010000101010",
1815 => "111111101000110000110100",
1816 => "000000010110001110000111",
1817 => "000000100011111101011111",
1818 => "000000001010010010001100",
1819 => "111111111101101000111010",
1820 => "000000011010101101100111",
1821 => "000000111010110001100111",
1822 => "000000111001110001010010",
1823 => "000000110100000110110001",
1824 => "000000111101100111101100",
1825 => "000001011111001001000100",
1826 => "000001111110010011010100",
1827 => "000001101111101111101110",
1828 => "000001100111111010000010",
1829 => "000001111000011101110101",
1830 => "000001111010100000100010",
1831 => "000010001001110110011001",
1832 => "000010010010011000011000",
1833 => "000010000001011101100111",
1834 => "000010010100001111111111",
1835 => "000011000011001111001010",
1836 => "000011011011100000010100",
1837 => "000011010110110011111110",
1838 => "000011101110100110011011",
1839 => "000100110110001000110011",
1840 => "000100011011101110011101",
1841 => "000010011110000110111011",
1842 => "000010000001000110001000",
1843 => "000001110000100000010010",
1844 => "111111110000101111000011",
1845 => "111111110010100001101100",
1846 => "000011001010110110101100",
1847 => "000101100011010100100100",
1848 => "000101010010011100100010",
1849 => "000100101111010011010100",
1850 => "000101001000000001110110",
1851 => "000101100001100000011110",
1852 => "000101010101100100001110",
1853 => "000101001010111100100011",
1854 => "000101000000101000010111",
1855 => "000100100001100011010011",
1856 => "000100001001111101000010",
1857 => "000011100011000001101011",
1858 => "000010001100010111010000",
1859 => "000001000100010011010001",
1860 => "000001010000100110001001",
1861 => "000010010100111110111111",
1862 => "000010111011000111001010",
1863 => "000011011101001010010010",
1864 => "000100111010110101010011",
1865 => "000101110010101000100100",
1866 => "000101001011011010001011",
1867 => "000100100111110100110110",
1868 => "000101000011000001100011",
1869 => "000101110101101111010010",
1870 => "000101100000100010101010",
1871 => "000100000100110010110001",
1872 => "000011010111100111100111",
1873 => "000010111110101000101000",
1874 => "000001100110111011010011",
1875 => "000000100111010100101111",
1876 => "000001000100011111101100",
1877 => "000001110001110111011111",
1878 => "000010001001100001111111",
1879 => "000010111100001001001000",
1880 => "000011111100010100010100",
1881 => "000100011010111000010001",
1882 => "000100101011110111011000",
1883 => "000100100010011101101010",
1884 => "000011001110011100110111",
1885 => "000001101001011100111110",
1886 => "000001001001000000100110",
1887 => "000001010011011001101011",
1888 => "000001011000011000110110",
1889 => "000001101010100110110101",
1890 => "000010001011000111111111",
1891 => "000010010101011000111001",
1892 => "000010001001010110100101",
1893 => "000010000001010110100111",
1894 => "000010001010111010110011",
1895 => "000010001110011000110110",
1896 => "000001100011110010101101",
1897 => "000000001101011101011010",
1898 => "111110100101100000111100",
1899 => "111101001101011000111101",
1900 => "111100101101111111000110",
1901 => "111101000011000100101011",
1902 => "111101100011110110101001",
1903 => "111110000101010100001010",
1904 => "111110111011111111111101",
1905 => "000000001011111011110000",
1906 => "000001011101111110111100",
1907 => "000010000001101111010000",
1908 => "000001010101011101010100",
1909 => "000000010101000001010111",
1910 => "111111110001001011011111",
1911 => "111111001000101010001001",
1912 => "111110101101101000010110",
1913 => "111110101010111110000110",
1914 => "111110000111110011111011",
1915 => "111100111000001011010101",
1916 => "111011010111111111000110",
1917 => "111010101000111011101100",
1918 => "111011010110000111111011",
1919 => "111100010111010111010001",
1920 => "111100110010010101011101",
1921 => "111100111101011011011001",
1922 => "111101011111111111111100",
1923 => "111110010101100000011100",
1924 => "111110100000101000111101",
1925 => "111110000100100011100001",
1926 => "111101101010011100000111",
1927 => "111101000000111100011001",
1928 => "111100010010001110010110",
1929 => "111011111110101011110001",
1930 => "111100000100110001111011",
1931 => "111100010011100001101111",
1932 => "111100000110100101011010",
1933 => "111011011011011011111100",
1934 => "111011001011011000110100",
1935 => "111011101101101111111011",
1936 => "111100001100110011001011",
1937 => "111011110100100101100011",
1938 => "111010101100000110110100",
1939 => "111001100111101101011110",
1940 => "111001100011000110110110",
1941 => "111010001000011110100000",
1942 => "111010011011111010101110",
1943 => "111010110100101000001001",
1944 => "111011011000111001110111",
1945 => "111011100111111011100000",
1946 => "111011111010001101001100",
1947 => "111100010101101001010101",
1948 => "111100100101000110001111",
1949 => "111100100010011011100010",
1950 => "111011111100100101001110",
1951 => "111011001101100010011101",
1952 => "111011001001111001001000",
1953 => "111011101010001110110111",
1954 => "111011111000000010001110",
1955 => "111011001001010100001110",
1956 => "111001110111001001001000",
1957 => "111001000011110010111000",
1958 => "111001000101100000100011",
1959 => "111001101101111101000110",
1960 => "111011000000010010001010",
1961 => "111100101101111101001011",
1962 => "111101111011111110110011",
1963 => "111110011000000100100000",
1964 => "111110101001000100110000",
1965 => "111110110001001000001000",
1966 => "111110000110101100010100",
1967 => "111100101111010000111100",
1968 => "111011110110001010011100",
1969 => "111011111010110110011111",
1970 => "111100001000000110000101",
1971 => "111100000000001110000111",
1972 => "111011110100110001101001",
1973 => "111011111001011000110011",
1974 => "111100011010001011111001",
1975 => "111101001010000111010001",
1976 => "111101101100110110111110",
1977 => "111110000111000001101111",
1978 => "111110110101110100111100",
1979 => "111111011010011011111000",
1980 => "111111001000100100111001",
1981 => "111110110001010010101100",
1982 => "111110110011101101110111",
1983 => "111110101011000001010011",
1984 => "111110010000011100011100",
1985 => "111101110111011110010000",
1986 => "111110001001011101111011",
1987 => "111111001110010110011100",
1988 => "000000000010101101100110",
1989 => "000000010110101110110011",
1990 => "000000101111011010011010",
1991 => "000001000010011110001011",
1992 => "000000110110001010001101",
1993 => "000000011101011111101100",
1994 => "000000011001001100010101",
1995 => "000000011110011011100011",
1996 => "000000011011010101100111",
1997 => "000000001110011111011111",
1998 => "000000001111010000111011",
1999 => "000001000010010010001101",
2000 => "000001110011001000000111",
2001 => "000010001010111001110011",
2002 => "000011000011001000110111",
2003 => "000011100011100000011001",
2004 => "000011101011010100111000",
2005 => "000100100001100110011011",
2006 => "000100010011010110111111",
2007 => "000010111111001101100100",
2008 => "000011011100111010100110",
2009 => "000100100001000010111011",
2010 => "000011011001110001010010",
2011 => "000001101111010101111110",
2012 => "000010000000111101101001",
2013 => "000011001101011011011110",
2014 => "000011110110010001101111",
2015 => "000100010010101010001001",
2016 => "000100110010000011011010",
2017 => "000101011100100110101000",
2018 => "000101101010001111011100",
2019 => "000011100111011101100010",
2020 => "000000100010001011100001",
2021 => "111111111110011011001000",
2022 => "000010011011100111000011",
2023 => "000101011011111000000011",
2024 => "000110100101010101000110",
2025 => "000110000100100000111000",
2026 => "000110001000010000111110",
2027 => "000110100111101111110010",
2028 => "000110010010010001111101",
2029 => "000110001010100111010010",
2030 => "000110100000011011111000",
2031 => "000110011011101000001011",
2032 => "000110000101000110110101",
2033 => "000100101001111101110000",
2034 => "000010010111010111100110",
2035 => "000001100011010001100001",
2036 => "000001110001110101111001",
2037 => "000001100000011010010001",
2038 => "000010000000000110100001",
2039 => "000011111000011100100101",
2040 => "000101100111010101111011",
2041 => "000110010110000110000000",
2042 => "000110011011010110011110",
2043 => "000110001111111101000111",
2044 => "000110010010010110101111",
2045 => "000110111010000110110100",
2046 => "000111001011100011011000",
2047 => "000110010111100000010011",
2048 => "000101010010010101100001",
2049 => "000100001001010011100011",
2050 => "000010011111010101101100",
2051 => "000000111001110100001001",
2052 => "000000010111111010100000",
2053 => "000000111011110110010010",
2054 => "000001100111001100100100",
2055 => "000010001110100000100010",
2056 => "000011100110111001101100",
2057 => "000101011100100101000011",
2058 => "000110011100100101110000",
2059 => "000110000010101100111001",
2060 => "000100110111011110100011",
2061 => "000011110110011000000111",
2062 => "000011001110110010000010",
2063 => "000010101101010100110011",
2064 => "000001111010001000010000",
2065 => "000001011001100111000111",
2066 => "000010001000011110111011",
2067 => "000011001000101010011100",
2068 => "000011000010100011110011",
2069 => "000010001111110000100100",
2070 => "000001011011010100000101",
2071 => "000000110010011011001101",
2072 => "000000010010110100001111",
2073 => "111111100001110111001110",
2074 => "111110100010100010001111",
2075 => "111101111011111001000111",
2076 => "111101111100001101001011",
2077 => "111110100011010110011111",
2078 => "111111101110110001000011",
2079 => "000000101101101010100111",
2080 => "000000111010100111001000",
2081 => "000000110111101100111010",
2082 => "000000111101011100101000",
2083 => "000001001100100100110001",
2084 => "000001011111011001111101",
2085 => "000001000111111111101001",
2086 => "111111111001000001001111",
2087 => "111110101010010100001000",
2088 => "111110000011110110110010",
2089 => "111101110110111010011100",
2090 => "111101100110001001110111",
2091 => "111101001101000101010110",
2092 => "111100011011000001011011",
2093 => "111011001001011101000110",
2094 => "111010010011111010010111",
2095 => "111010010010000001010011",
2096 => "111010100110110100100000",
2097 => "111011011001001000011000",
2098 => "111100100101001110101010",
2099 => "111101110001011110011100",
2100 => "111110110011100000110010",
2101 => "111111011011100010100011",
2102 => "111111100100111100101111",
2103 => "111111001011101010100001",
2104 => "111101111010100100001010",
2105 => "111100010010100111101010",
2106 => "111011010111101010100011",
2107 => "111011000000100101001101",
2108 => "111010010111101111101100",
2109 => "111001010111000010011100",
2110 => "111000011111110011110100",
2111 => "111000011100100010011010",
2112 => "111001010001100001001100",
2113 => "111010001100101010000010",
2114 => "111010110011011011001011",
2115 => "111011001011010001000001",
2116 => "111011001111010010010100",
2117 => "111011000111000010010110",
2118 => "111011000010001101110010",
2119 => "111011000100011001001001",
2120 => "111011010000000100000011",
2121 => "111011100000010101101011",
2122 => "111011100111111111111000",
2123 => "111011101111001110111111",
2124 => "111100001011001111011000",
2125 => "111100101100110000011011",
2126 => "111100110000110011010000",
2127 => "111100000011000101111111",
2128 => "111010101000000000110010",
2129 => "111001100000000000010001",
2130 => "111001011100100000010001",
2131 => "111001100111111100001010",
2132 => "111001001100100111101101",
2133 => "111000100111101111101101",
2134 => "111000111100010011001110",
2135 => "111010011101101110100101",
2136 => "111100010100110110011001",
2137 => "111101111100011100001111",
2138 => "111111001010000010111110",
2139 => "111111100010101000000000",
2140 => "111111010111011011011111",
2141 => "111111001101011111001110",
2142 => "111110111100010110111011",
2143 => "111110010101100101010111",
2144 => "111101100101000011000100",
2145 => "111101000110100011010111",
2146 => "111100111110101100100001",
2147 => "111100110000011100100000",
2148 => "111100001100010001010000",
2149 => "111011100111001101100110",
2150 => "111011101100100010001100",
2151 => "111100100000010110000110",
2152 => "111101010101000101111111",
2153 => "111110001010011110000001",
2154 => "111111011000111011101110",
2155 => "000000100110111111110111",
2156 => "000001011110011111111110",
2157 => "000001111101000110011011",
2158 => "000001111110011000111000",
2159 => "000001101111011001110000",
2160 => "000001010001111101110010",
2161 => "000000101010000000111101",
2162 => "000000010011010011111000",
2163 => "000000000100000000001011",
2164 => "111111110011000010011000",
2165 => "111111110111010110110000",
2166 => "000000001000111001111100",
2167 => "000000101000010100000011",
2168 => "000001010011010100111001",
2169 => "000001101001011000010111",
2170 => "000001111101111110100010",
2171 => "000010010100100110000011",
2172 => "000010010001100011001000",
2173 => "000010010010111000010101",
2174 => "000010001111110000001011",
2175 => "000010000010100101101111",
2176 => "000010100001110001011110",
2177 => "000011000010000101011110",
2178 => "000011001100110001011111",
2179 => "000100011101001001100001",
2180 => "000110011000101011111000",
2181 => "000111001110111011110101",
2182 => "000110101111111101010000",
2183 => "000101101101100110010100",
2184 => "000100111011110100111000",
2185 => "000100001110011011000111",
2186 => "000010110000110110001000",
2187 => "000001100000110010001110",
2188 => "000001111100101011011101",
2189 => "000010110011001010110011",
2190 => "000010110001101111000011",
2191 => "000011001011010110111101",
2192 => "000011001010101000100010",
2193 => "000000100111001000100111",
2194 => "111111010100001010000101",
2195 => "000011010001000101100101",
2196 => "000111110011000011001000",
2197 => "000111111010011001000110",
2198 => "000110010010010011001010",
2199 => "000110010110111111000111",
2200 => "000110111100010000001010",
2201 => "000110000110111011010100",
2202 => "000100101111001011011010",
2203 => "000100010101001110001000",
2204 => "000100001011101000111010",
2205 => "000011011110000010000100",
2206 => "000010110000100000001010",
2207 => "000001101101010110100011",
2208 => "000000001100000011100010",
2209 => "111111111001011001101000",
2210 => "000001000100001011011111",
2211 => "000010001010010110001000",
2212 => "000011011101100010011011",
2213 => "000101101100101000101011",
2214 => "000111001010101101101000",
2215 => "000110010101111111000000",
2216 => "000100110001001011000111",
2217 => "000100101100010111110011",
2218 => "000101101111111100010100",
2219 => "000101111110011000001100",
2220 => "000101010110100010010011",
2221 => "000101001110110001010101",
2222 => "000100101101110000100111",
2223 => "000010100101110000111010",
2224 => "000000110011101011000000",
2225 => "000000110110111000000100",
2226 => "000000111001111000101010",
2227 => "111111111001001110101010",
2228 => "111111101110111110100000",
2229 => "000001011011000110100010",
2230 => "000011000110110100001100",
2231 => "000011101110101001100100",
2232 => "000100001010010111111111",
2233 => "000100010000110101001110",
2234 => "000011110101010011100101",
2235 => "000011110110100000001010",
2236 => "000100000111001111101010",
2237 => "000011110001000101101100",
2238 => "000010111000011101101001",
2239 => "000001110011101011011000",
2240 => "000000111010010000011000",
2241 => "111111110110110001101101",
2242 => "111110100111101000100001",
2243 => "111110100001110100111100",
2244 => "111111000101100011101101",
2245 => "111110110011110000000011",
2246 => "111110100110001001111001",
2247 => "111110111010100100100010",
2248 => "111111001110110101100001",
2249 => "000000000010101110001100",
2250 => "000000100100010010010100",
2251 => "111111111010011010111101",
2252 => "111111100000010100100111",
2253 => "111111111011100000110010",
2254 => "000000011001111000101101",
2255 => "000000110000110011010000",
2256 => "000000110010011110011111",
2257 => "000000011100001110111001",
2258 => "000000000000001000100111",
2259 => "111111010111010000010011",
2260 => "111110101011000000011011",
2261 => "111110000011010110111000",
2262 => "111101001101011010010001",
2263 => "111100010001011110011001",
2264 => "111011100011111000110100",
2265 => "111011000110010110010010",
2266 => "111010101101011011010100",
2267 => "111010001101010001111110",
2268 => "111001111011110110101010",
2269 => "111010001101110001011101",
2270 => "111010111010000010111010",
2271 => "111100001100111000011000",
2272 => "111101110110110010001100",
2273 => "111110111001010010001101",
2274 => "111111010100110000111010",
2275 => "111111001111110110011100",
2276 => "111110000000110011111001",
2277 => "111100011110110110001101",
2278 => "111011111000101011000110",
2279 => "111011010100101000100100",
2280 => "111010000100010011100011",
2281 => "111000101011010111010101",
2282 => "110111100101010011101010",
2283 => "110111010011000111001000",
2284 => "110111100011111101111111",
2285 => "110111011111100011100000",
2286 => "110111101101110101101010",
2287 => "111000101111101010101000",
2288 => "111001110110011000111100",
2289 => "111010111010010111111111",
2290 => "111011110010100111101010",
2291 => "111100000110000100110101",
2292 => "111100010000111110110111",
2293 => "111100100100111010001001",
2294 => "111100111010110001100101",
2295 => "111100111110101011101011",
2296 => "111100001101000101010110",
2297 => "111011001110000100111100",
2298 => "111010111110010010010000",
2299 => "111010111101100001000010",
2300 => "111010011011100100000001",
2301 => "111001010001000001101011",
2302 => "110111111101011011001001",
2303 => "110111011001011100100000",
2304 => "110111111001010110110110",
2305 => "111001001000100100111101",
2306 => "111010010011111010000100",
2307 => "111011000011000101110101",
2308 => "111100010110100001000111",
2309 => "111110001010100110110010",
2310 => "111110111000000100101110",
2311 => "111110100111000001111000",
2312 => "111110101001001000001000",
2313 => "111111001000000100011010",
2314 => "111111100100101100011000",
2315 => "111111100001011011001100",
2316 => "111111001000110001110111",
2317 => "111110111001100101011100",
2318 => "111110011101000010010011",
2319 => "111101011010010010000001",
2320 => "111100001101110111011000",
2321 => "111011100010111111011110",
2322 => "111011101100011011100000",
2323 => "111100010101110011011001",
2324 => "111101000100001110001101",
2325 => "111101110100001110000100",
2326 => "111110111011011101010000",
2327 => "000000110110010110011111",
2328 => "000010111101101101111011",
2329 => "000100000001001010110110",
2330 => "000100000000010000101001",
2331 => "000011110000101010000100",
2332 => "000011100010101101010010",
2333 => "000011000000110011000010",
2334 => "000010001001111111000101",
2335 => "000001011110101111001010",
2336 => "000000111001100110011110",
2337 => "000000001100000000001110",
2338 => "111111111110010101010001",
2339 => "000000100010010110000000",
2340 => "000001011111101100010000",
2341 => "000010010010011111001101",
2342 => "000010011011010101000011",
2343 => "000010100011011101111101",
2344 => "000010111011011001010000",
2345 => "000010100111111111110000",
2346 => "000010010010100100011101",
2347 => "000010111110001001111011",
2348 => "000100001010100001101000",
2349 => "000101011011011111011001",
2350 => "000110001010100000100010",
2351 => "000110001010101100110110",
2352 => "000110011001000011010100",
2353 => "000110100101100110100001",
2354 => "000110010100011110010001",
2355 => "000101110110011110001001",
2356 => "000100100000101110111000",
2357 => "000011001100000100101001",
2358 => "000011001000100001111011",
2359 => "000010001111001100001111",
2360 => "111111101000100000000111",
2361 => "111101000111010011010010",
2362 => "111011011100010100010101",
2363 => "111100011000000000001011",
2364 => "000000111000110110101000",
2365 => "000101000100011101101010",
2366 => "000110010000100101000101",
2367 => "000110100111001001101100",
2368 => "000111011111110000111011",
2369 => "001000010001110100111111",
2370 => "001000100101010111000101",
2371 => "000111111101101011011000",
2372 => "000110100110100111110011",
2373 => "000101010101000110011111",
2374 => "000011101001011010011000",
2375 => "000001000010001111100011",
2376 => "111110101001010111011100",
2377 => "111101010011000010010100",
2378 => "111100110101011001011110",
2379 => "111101010011100101001001",
2380 => "111110101010010001101001",
2381 => "000000110100000011110110",
2382 => "000011001110100100101010",
2383 => "000100101000111110100011",
2384 => "000101011010011111011110",
2385 => "000110101100010100001001",
2386 => "000111100110110001011010",
2387 => "000111100111101111001110",
2388 => "000111010100100110011110",
2389 => "000110001000011000001111",
2390 => "000100001000100111001101",
2391 => "000010011000010110011111",
2392 => "000000110000000000111110",
2393 => "111111110001010011111110",
2394 => "000000000110111101110010",
2395 => "000000010100111110001111",
2396 => "000000010000010100101101",
2397 => "000001011111100011001100",
2398 => "000011010110001000011001",
2399 => "000100011010110100100001",
2400 => "000100110111001110010100",
2401 => "000100100000000111011100",
2402 => "000011011010001001111100",
2403 => "000010001111001001100000",
2404 => "000000101101111100110000",
2405 => "111111011110011001110101",
2406 => "111111110101011010101100",
2407 => "000000111101000010001001",
2408 => "000001101111100100010001",
2409 => "000010010101111001111100",
2410 => "000010011110010110010100",
2411 => "000010010110100011111101",
2412 => "000010100100001010001011",
2413 => "000010101101001001110011",
2414 => "000010100011011010001101",
2415 => "000001110011000000101101",
2416 => "000000000010111000110001",
2417 => "111110100000100010010001",
2418 => "111101111001001110000011",
2419 => "111101010001010001100000",
2420 => "111100101101110110011011",
2421 => "111101000000000100111101",
2422 => "111110001010100001110110",
2423 => "111111111011100011110001",
2424 => "000001100100101011001011",
2425 => "000010011100110011010010",
2426 => "000010101001010001101111",
2427 => "000010010111001101101001",
2428 => "000001101001111100000100",
2429 => "000000100000101111000010",
2430 => "111111010110100000010011",
2431 => "111110100010111101101101",
2432 => "111101000111111101000101",
2433 => "111010101100101111010101",
2434 => "111000110100000111111100",
2435 => "111000010010101101000001",
2436 => "111000111001010001010110",
2437 => "111010100100111100010111",
2438 => "111100100101011011110111",
2439 => "111110001001011000111111",
2440 => "111111011001010010101100",
2441 => "000000001011101110111101",
2442 => "000000011000000010110111",
2443 => "000000001101111001101100",
2444 => "111111010100001110001110",
2445 => "111101100101001000011110",
2446 => "111100000010000110101010",
2447 => "111011001101001000100011",
2448 => "111010110101100011001000",
2449 => "111010101010000101100100",
2450 => "111010000110110000011110",
2451 => "111001010011011101001110",
2452 => "111001011111111000100010",
2453 => "111010101000001000100111",
2454 => "111011011011110100100101",
2455 => "111011110001110111101101",
2456 => "111011110001111100011011",
2457 => "111011010101010010011011",
2458 => "111011001011001110000010",
2459 => "111011101011111010101111",
2460 => "111100010111010100111010",
2461 => "111100111001101100000001",
2462 => "111101000010000011101101",
2463 => "111100110011001111001011",
2464 => "111100110010100010101001",
2465 => "111101001110111010100001",
2466 => "111110000000000001100100",
2467 => "111110110001101111111011",
2468 => "111111000011011000011010",
2469 => "111110100000110000101011",
2470 => "111101000010110110110010",
2471 => "111011001100101010001011",
2472 => "111010001000110001000000",
2473 => "111010000101011101011011",
2474 => "111010010011100001011100",
2475 => "111010101011110111000111",
2476 => "111011111100000101111001",
2477 => "111110000110110011001110",
2478 => "111111110111000001011000",
2479 => "000000100101000101011010",
2480 => "000001010010110111000110",
2481 => "000010011001001010001110",
2482 => "000011011000101010001100",
2483 => "000100000100010000110100",
2484 => "000011111010101001001110",
2485 => "000010110111101011101101",
2486 => "000001110001101110101110",
2487 => "000000100110000100101001",
2488 => "111110111101100101100001",
2489 => "111101101000110011001100",
2490 => "111101010100011001001011",
2491 => "111101110101111111100111",
2492 => "111110101010001011100001",
2493 => "111111011010100100111000",
2494 => "000000011110111110100101",
2495 => "000010001011101001101000",
2496 => "000100000011101010001100",
2497 => "000101100110110111011110",
2498 => "000110100110000010101101",
2499 => "000110111000001010110100",
2500 => "000110011100000010100110",
2501 => "000101100000001001111111",
2502 => "000100110011110010101001",
2503 => "000100011111010101111100",
2504 => "000011100001001101101011",
2505 => "000010001000000101100001",
2506 => "000001100111001010001110",
2507 => "000001101110101110100010",
2508 => "000010000011100010101111",
2509 => "000010110100000001001010",
2510 => "000011010101100111000001",
2511 => "000011101000110001111100",
2512 => "000100100000111011010110",
2513 => "000101010111111001000111",
2514 => "000101100001011110100100",
2515 => "000101001011001010001100",
2516 => "000100111111110101101101",
2517 => "000101110001110100001011",
2518 => "000110011000010101101010",
2519 => "000101101111011111110001",
2520 => "000101011101110110010001",
2521 => "000101011110110100100110",
2522 => "000100011011010011100010",
2523 => "000011100011000110000001",
2524 => "000010100111011110111101",
2525 => "111111100001001010010111",
2526 => "111011010100100111100100",
2527 => "111000111110011010000101",
2528 => "111010100001100001110000",
2529 => "111111000110001001001111",
2530 => "000010010110101001100110",
2531 => "000010100111111011011110",
2532 => "000010011110101001100000",
2533 => "000011000111010001000110",
2534 => "000100000111111110000101",
2535 => "000100111000100011101000",
2536 => "000100011100000111001100",
2537 => "000011101110000000010110",
2538 => "000011101000111000011100",
2539 => "000010100000001001100000",
2540 => "111111111011011100100001",
2541 => "111101110101010111101110",
2542 => "111100100000110101100010",
2543 => "111011001001100101010011",
2544 => "111010001111010110010011",
2545 => "111010101110111010001110",
2546 => "111100110000111010010010",
2547 => "111111001001110011000100",
2548 => "000000000000110000101111",
2549 => "111111101100111111100111",
2550 => "000000101100011111010110",
2551 => "000011000111100010100001",
2552 => "000101000010001101010000",
2553 => "000101101011101110011101",
2554 => "000100101011001011010100",
2555 => "000010000110110111010100",
2556 => "111111100011011010000010",
2557 => "111101110101100101001101",
2558 => "111100110100101010100111",
2559 => "111100011010010011001011",
2560 => "111011110110110010001100",
2561 => "111011100010111011100000",
2562 => "111101001101001010110011",
2563 => "000000011000000111100011",
2564 => "000010111011011101111000",
2565 => "000011110011010000100100",
2566 => "000011000100010001011001",
2567 => "000001100111000111001000",
2568 => "000000001000100001110111",
2569 => "111110011010011001010000",
2570 => "111100101100100100011000",
2571 => "111011101011011000110101",
2572 => "111011011101111011110111",
2573 => "111011111111001010101011",
2574 => "111100101111101101110001",
2575 => "111101010100010001101000",
2576 => "111110100011000110010010",
2577 => "000000110000110000001010",
2578 => "000010100110000111000010",
2579 => "000010111100000101010011",
2580 => "000001101001000111101101",
2581 => "111111101100100001111011",
2582 => "111110101011111000110011",
2583 => "111110001100001110001101",
2584 => "111100111011011111010000",
2585 => "111011101001101011111101",
2586 => "111011001000011101010100",
2587 => "111010111101001001010111",
2588 => "111011001110010110000111",
2589 => "111100000110011010010000",
2590 => "111101000111100010001010",
2591 => "111101101111000001111000",
2592 => "111101110011110110011110",
2593 => "111101111101100011000111",
2594 => "111110100010001001100101",
2595 => "111110111100011001100101",
2596 => "111110100010110110011000",
2597 => "111100111110000011100010",
2598 => "111010101111001011110100",
2599 => "111000111110100111101001",
2600 => "110111111110011000100101",
2601 => "110111101011001001100101",
2602 => "111000000111110100010010",
2603 => "111001000101010000010101",
2604 => "111010100011111001000010",
2605 => "111100010110000001000111",
2606 => "111110000101000110101010",
2607 => "111111100110111111010000",
2608 => "111111110010100000010101",
2609 => "111110001000001110111011",
2610 => "111100001011110100010101",
2611 => "111010111001111010000110",
2612 => "111010000100010100011100",
2613 => "111001001010001100110110",
2614 => "110111100101000110011111",
2615 => "110110010011011100101000",
2616 => "110110101011100111110000",
2617 => "111000000011101000011010",
2618 => "111001100011001011000010",
2619 => "111011000011011001110001",
2620 => "111100001110011110001001",
2621 => "111100110101111001001000",
2622 => "111101000011100011111001",
2623 => "111101010011100101010010",
2624 => "111101111011001000010111",
2625 => "111110010100010101010100",
2626 => "111101101110110001010001",
2627 => "111100101000111111101101",
2628 => "111100001001001111101100",
2629 => "111100001101001001010000",
2630 => "111100000010001010000010",
2631 => "111011110110001010001011",
2632 => "111100001100100101111010",
2633 => "111100110010001111110001",
2634 => "111100111111100010101001",
2635 => "111100100000111101110100",
2636 => "111100010011101011000110",
2637 => "111101100110110010101011",
2638 => "111111001110001101101001",
2639 => "111111010111110011011011",
2640 => "111110111011101010111111",
2641 => "111111101011110100111100",
2642 => "000001010100111001010111",
2643 => "000010000010111110000011",
2644 => "000001101000001101011001",
2645 => "000001101100000001011101",
2646 => "000010011111001010110010",
2647 => "000011000000110101001100",
2648 => "000011000110011111001111",
2649 => "000011000001101101000110",
2650 => "000010111100110111111111",
2651 => "000010110000110100010011",
2652 => "000010001000100010100111",
2653 => "000001010110011011100110",
2654 => "000000111101100011010110",
2655 => "000001000111111101000001",
2656 => "000001100000100110111101",
2657 => "000001100111011011000100",
2658 => "000001111010011111101001",
2659 => "000011001110001000110101",
2660 => "000101010101001010000111",
2661 => "000111100001000111010001",
2662 => "001001000010001000010100",
2663 => "001001100101110010100000",
2664 => "001001010111101100101000",
2665 => "001000100111000011011000",
2666 => "001000000101010101000001",
2667 => "000111110001110000111101",
2668 => "000110101100001011110010",
2669 => "000101000101100101100111",
2670 => "000011101000101001111010",
2671 => "000011000110000100010001",
2672 => "000100001000000111011001",
2673 => "000100111011100110110000",
2674 => "000100111101110111101101",
2675 => "000110010000011110111011",
2676 => "000111101011001000110101",
2677 => "000111110001001011000010",
2678 => "001000010101010010110011",
2679 => "001001110111000011001110",
2680 => "001010110010111111010101",
2681 => "001001101100100100000000",
2682 => "000111110101011011011101",
2683 => "001000100101110111110110",
2684 => "001001110100110000100001",
2685 => "000111011111110110110100",
2686 => "000100001000010011000100",
2687 => "000001001011001111111000",
2688 => "111100111110011110100010",
2689 => "111010100110001010110011",
2690 => "111100111011100001110100",
2691 => "000001001110010100001110",
2692 => "000011101101011101100010",
2693 => "000011110100101010011011",
2694 => "000100100110011100110010",
2695 => "000111011011111101001101",
2696 => "001001010001011000010100",
2697 => "001000111000100011001000",
2698 => "001000001110001010110100",
2699 => "000111101011111010010010",
2700 => "000110011110111000101100",
2701 => "000100010101111000110010",
2702 => "000001010100010100111110",
2703 => "111110000110101100001110",
2704 => "111011110111011001110101",
2705 => "111011010100011111100110",
2706 => "111100010000111000010000",
2707 => "111110000010110010011010",
2708 => "000000001011110100001101",
2709 => "000010001011001011000010",
2710 => "000011001011101001110010",
2711 => "000011001010010101110010",
2712 => "000100000001000000110010",
2713 => "000110011011101010110001",
2714 => "000111011000010111001101",
2715 => "000101101001010100000101",
2716 => "000011111100011000101110",
2717 => "000010111001110011111000",
2718 => "000001001011010011110000",
2719 => "111111011010011000110110",
2720 => "111110100001100111010111",
2721 => "111101111011000101101011",
2722 => "111101000000111101011010",
2723 => "111100111101011000100101",
2724 => "111111010100000111111011",
2725 => "000010100101010011000011",
2726 => "000100010111001110110010",
2727 => "000101001100111111000001",
2728 => "000101100111110000001101",
2729 => "000100001110100110111010",
2730 => "000001010100001000011101",
2731 => "111111001010010110101000",
2732 => "111110001110100010110100",
2733 => "111101000100110000100110",
2734 => "111011110001101101000100",
2735 => "111011010010110011011010",
2736 => "111011010110001001011011",
2737 => "111100001111101001111000",
2738 => "111110110010100000001100",
2739 => "000001110100100100000110",
2740 => "000011011001101010110101",
2741 => "000010111101011110001111",
2742 => "000001110010001010000000",
2743 => "000001010111000010011001",
2744 => "000000111101011100100010",
2745 => "111111010101000011011100",
2746 => "111100110101011000010010",
2747 => "111010100000110000100110",
2748 => "111001110010110110000010",
2749 => "111011000111001110001100",
2750 => "111100101010101011111010",
2751 => "111101001010010110101101",
2752 => "111101000100101001100011",
2753 => "111101001101011000100010",
2754 => "111101110101111000110000",
2755 => "111110010111100101110011",
2756 => "111110011011010101010110",
2757 => "111110000100100001100110",
2758 => "111100101110000010001100",
2759 => "111010100000010000001010",
2760 => "111000100010001111011011",
2761 => "110111010011111110101111",
2762 => "110110110011000111111010",
2763 => "110110011111110001110110",
2764 => "110110001111011011001000",
2765 => "110111001110111110000001",
2766 => "111001110101111100001101",
2767 => "111100011110101010011001",
2768 => "111110000001001001110111",
2769 => "111110110010100100111100",
2770 => "111111000001111111010101",
2771 => "111110001100110100011110",
2772 => "111100100100001111110010",
2773 => "111011010101111101001110",
2774 => "111010010110000010110111",
2775 => "111000100000000101100100",
2776 => "110110001000101101110000",
2777 => "110100011100111011010111",
2778 => "110100010100011100111101",
2779 => "110101100110111011001111",
2780 => "110111001100100000111011",
2781 => "111000011011110001111101",
2782 => "111001011001100110101001",
2783 => "111010001001101110110010",
2784 => "111011000000001100001100",
2785 => "111100000110100111110010",
2786 => "111101000101101001000101",
2787 => "111101110110000101011011",
2788 => "111110010001101111101000",
2789 => "111101111110111001111011",
2790 => "111101001010000110110010",
2791 => "111100101110001111100101",
2792 => "111101001011000000111110",
2793 => "111101100101101110000000",
2794 => "111100100000101100011011",
2795 => "111010010110100101100000",
2796 => "111001000100011110010110",
2797 => "111001000110011011001011",
2798 => "111001101110110011011011",
2799 => "111011001101000101000000",
2800 => "111101010000101101101000",
2801 => "111110011011110101111000",
2802 => "111110100111100011101010",
2803 => "111111001110011001110111",
2804 => "000000100000001000110011",
2805 => "000001000111001110100100",
2806 => "000000101110010000111010",
2807 => "000000111010000011010110",
2808 => "000010010011010111000010",
2809 => "000011100001011100010100",
2810 => "000011110101001010110100",
2811 => "000011101110001101110000",
2812 => "000011010000110101000110",
2813 => "000010010010111001010100",
2814 => "000001001101110000011110",
2815 => "000000100010111001101001",
2816 => "000000010110000100010111",
2817 => "000000010011110111001110",
2818 => "000000010000010101101100",
2819 => "000000001101111110001000",
2820 => "000000011101101110101101",
2821 => "000001100001000010010011",
2822 => "000011100000111110001010",
2823 => "000101011001011000111011",
2824 => "000101111110011100011110",
2825 => "000110001101111100001010",
2826 => "000111100010001011110000",
2827 => "001000101000010000011010",
2828 => "001000001110001101010111",
2829 => "000111001110010000111111",
2830 => "000110000010110011111110",
2831 => "000100111111100101110111",
2832 => "000100110011100000010101",
2833 => "000100100001011010010101",
2834 => "000011101111100100110111",
2835 => "000011011010100101000001",
2836 => "000010100100101000111000",
2837 => "000001000001111000110111",
2838 => "000001101110000111100101",
2839 => "000100101101101010000100",
2840 => "000101100111100001010101",
2841 => "000011100011010111010010",
2842 => "000011011011011001000100",
2843 => "000111001010110010001110",
2844 => "001001111101111011001110",
2845 => "000111111010011111101010",
2846 => "000010110010001111011000",
2847 => "111110010100100011010100",
2848 => "111100010000110101101011",
2849 => "111100100111001000001010",
2850 => "111110101100001110101000",
2851 => "000000010001011101000011",
2852 => "000000000000001110000010",
2853 => "000000011001110000101001",
2854 => "000010011000101001100100",
2855 => "000011001110111010111000",
2856 => "000011001101011010110000",
2857 => "000100010000111110000010",
2858 => "000101011101010001100010",
2859 => "000101011001001001110010",
2860 => "000011101011010111111110",
2861 => "000001000101100111000101",
2862 => "111110110111010000011000",
2863 => "111100010011111011001110",
2864 => "111001110010010010110110",
2865 => "111001101101100001001000",
2866 => "111011101001000010110110",
2867 => "111101110000110111100101",
2868 => "000000000100001010111101",
2869 => "000001111001010110011100",
2870 => "000010011000111010101011",
2871 => "000010111011011111001001",
2872 => "000101001111101111111111",
2873 => "001000000000001101001000",
2874 => "000111110101101010101100",
2875 => "000100100001110010100000",
2876 => "000001010111110100001011",
2877 => "111111110111101000101000",
2878 => "111110101110001101010010",
2879 => "111101011011010010101101",
2880 => "111100101011000111000001",
2881 => "111100001010111100000010",
2882 => "111011111000111101100000",
2883 => "111101101100011010101000",
2884 => "000001101001011010000001",
2885 => "000100111101010000000111",
2886 => "000110110000011111111010",
2887 => "000111111101010111001100",
2888 => "001000000001110011010000",
2889 => "000110100100111010000101",
2890 => "000100111011010100000000",
2891 => "000100000100110001101010",
2892 => "000011000000001101101101",
2893 => "000000100111000110101000",
2894 => "111101110011001001011011",
2895 => "111011101100010010000100",
2896 => "111010111010010110001100",
2897 => "111100001110010101100001",
2898 => "111110100101100010010110",
2899 => "111111111110101100010000",
2900 => "000000011001010100111000",
2901 => "000001000111110111010101",
2902 => "000010110011110100001001",
2903 => "000100010011000110101011",
2904 => "000100000100001001010000",
2905 => "000010110111001110100111",
2906 => "000001111100100100101010",
2907 => "000001100010111111101010",
2908 => "000001101110101111110010",
2909 => "000001101000010001101000",
2910 => "000000110011000000001010",
2911 => "000000000110001000111111",
2912 => "111111011100101010010110",
2913 => "111110110110110001101101",
2914 => "111111000010100001101000",
2915 => "111111100000001111100001",
2916 => "111111011011000100000000",
2917 => "111110011010011100111100",
2918 => "111100101001000011111010",
2919 => "111011001101111000111100",
2920 => "111010011101001100110110",
2921 => "111010000010101010000101",
2922 => "111010001000001000110010",
2923 => "111010000111010001011010",
2924 => "111001110010101100011011",
2925 => "111010100111011001101001",
2926 => "111101010001111011111010",
2927 => "000000010010111100011000",
2928 => "000001100110100000101000",
2929 => "000001000100011110001110",
2930 => "000000010101000110001110",
2931 => "000000000111111010010010",
2932 => "000000000100111101011110",
2933 => "111111011001111111101111",
2934 => "111101000100010000010110",
2935 => "111001100101001010001111",
2936 => "110110111010111001101110",
2937 => "110101111000011110111001",
2938 => "110101110100100010110101",
2939 => "110110001010001011010101",
2940 => "110110110001010011011010",
2941 => "110111010100001100001111",
2942 => "110111101111001111100010",
2943 => "111001000110011010111101",
2944 => "111011110011101001010011",
2945 => "111110100111110111110001",
2946 => "000000100101101000000100",
2947 => "000001101110111110001110",
2948 => "000010010110010111101110",
2949 => "000010011101010001110001",
2950 => "000010000001101001000110",
2951 => "000001100011100011000001",
2952 => "000000110101100000101100",
2953 => "111110100111101001001011",
2954 => "111011001100110010111100",
2955 => "111000100101010010000100",
2956 => "110111110110000010010110",
2957 => "111000001011101000111011",
2958 => "111000100111101111001100",
2959 => "111001101100100110001101",
2960 => "111011110010101001101001",
2961 => "111101110101001000111111",
2962 => "111111101001010010001110",
2963 => "000001111110010110100010",
2964 => "000011111101101101110100",
2965 => "000100011100001010001101",
2966 => "000100010100010010101111",
2967 => "000100111010101110111011",
2968 => "000101100010000110100000",
2969 => "000101001011100110110001",
2970 => "000100011010111000100100",
2971 => "000011011100000101100110",
2972 => "000001110011101111100000",
2973 => "000000000100001111011010",
2974 => "111111000000011000110011",
2975 => "111110111011001101111010",
2976 => "111111011001100101011011",
2977 => "111111100010010101110010",
2978 => "111111010101101001011101",
2979 => "111111011010001101110110",
2980 => "000000100101100010011101",
2981 => "000011010111011001110010",
2982 => "000101100111010110111100",
2983 => "000101001101101100100110",
2984 => "000100001010000110010101",
2985 => "000101001011000101111010",
2986 => "000111011100101101001011",
2987 => "000111110111001100000100",
2988 => "000101111011010111010110",
2989 => "000101011000001010010110",
2990 => "000110111110100001111110",
2991 => "000110101010011011001110",
2992 => "000100001010010110101010",
2993 => "000011000011111010100001",
2994 => "000011101111101001010101",
2995 => "000011100000000011000010",
2996 => "000000110001101000111000",
2997 => "111110000100010101111010",
2998 => "111110100010111110100110",
2999 => "111111110110110110001111",
3000 => "111111000011011100110101",
3001 => "111110110011010001100001",
3002 => "000000001001001010011000",
3003 => "111110111100010010011100",
3004 => "111011001000010010000000",
3005 => "111010110100100011110100",
3006 => "111111110100000111000001",
3007 => "000100000101100000100101",
3008 => "000011101111111101100010",
3009 => "000010010011000011000001",
3010 => "000011000000101011111111",
3011 => "000011110100111001111100",
3012 => "000010011000000001001000",
3013 => "111111111100111010000000",
3014 => "111110011111111110010000",
3015 => "111101111100100000001111",
3016 => "111101010101111101100111",
3017 => "111100000010011010111000",
3018 => "111010010111011001010001",
3019 => "111001011001100110010101",
3020 => "111001000000000010010001",
3021 => "111000101111011110001000",
3022 => "111001110101001110001100",
3023 => "111100100010100010111010",
3024 => "111110111011000011011110",
3025 => "111111101010010001001010",
3026 => "111111011111011111111101",
3027 => "000000101001100100011000",
3028 => "000100000000101100011010",
3029 => "000110100110101111001100",
3030 => "000110000100101110010111",
3031 => "000100011101000101111010",
3032 => "000011001101110101011110",
3033 => "000000110011011111001111",
3034 => "111101011001001100000111",
3035 => "111011011111010010001010",
3036 => "111011010011110011111010",
3037 => "111010100101110100110111",
3038 => "111001001100011100010101",
3039 => "111001101100010000010011",
3040 => "111100100111100000100111",
3041 => "111111111011100111101011",
3042 => "000010111110110110110100",
3043 => "000101101111100110101100",
3044 => "000110110101010010010110",
3045 => "000110000010110011100000",
3046 => "000101001010011001000101",
3047 => "000101101110011000010110",
3048 => "000111011111011110101010",
3049 => "001000001100111000100001",
3050 => "000110100000100110110100",
3051 => "000011110100001000101101",
3052 => "000001010111111011000000",
3053 => "111111101101011010011000",
3054 => "111111001000000000101011",
3055 => "111110001001011110010100",
3056 => "111011111101110000101000",
3057 => "111010011000011110101101",
3058 => "111010101010011110011110",
3059 => "111100101000001000100010",
3060 => "111111010001001001001011",
3061 => "000000110100000010010001",
3062 => "000001010100010010000001",
3063 => "000010100111010110001001",
3064 => "000100110110101011001100",
3065 => "000110100111001010011100",
3066 => "000110111101101010101101",
3067 => "000101110111001101000100",
3068 => "000100001011010111111011",
3069 => "000011001110001100111011",
3070 => "000011001011111100000101",
3071 => "000010111001111001111110",
3072 => "000001111000111100000110",
3073 => "000000100100001001000110",
3074 => "111110100001011111000101",
3075 => "111011101101000010001011",
3076 => "111001011110001110010011",
3077 => "111000010010100001100100",
3078 => "110111011000000001000100",
3079 => "110110101001110110100100",
3080 => "110110101011101000110000",
3081 => "110111110100101010100000",
3082 => "111001111111010000011001",
3083 => "111100100010000000111001",
3084 => "111110110000011001110111",
3085 => "000000010100111111001101",
3086 => "000001001010110111101111",
3087 => "000001110011000101100101",
3088 => "000011001000011000111010",
3089 => "000100011111101001001011",
3090 => "000011101011001001001110",
3091 => "000000100001100001100110",
3092 => "111101000111111010001111",
3093 => "111010011001010100011011",
3094 => "111000001101010110000111",
3095 => "110110011111101101110000",
3096 => "110100101011011111111011",
3097 => "110010101101110011100010",
3098 => "110001101000010101010000",
3099 => "110001111110010110001100",
3100 => "110011100011010110011110",
3101 => "110110010001110110100010",
3102 => "111010000000101111001100",
3103 => "111101101101110110010111",
3104 => "000000001101101010010101",
3105 => "000010001011111111100001",
3106 => "000101001110111101101100",
3107 => "001000101001000111000100",
3108 => "001001101111011000110100",
3109 => "000111110101000110000111",
3110 => "000101000011100100111110",
3111 => "000010100001010110011001",
3112 => "111111100001001011001011",
3113 => "111100111000000011100000",
3114 => "111011110101010110100100",
3115 => "111011001011110110010100",
3116 => "111001101010010001101100",
3117 => "111000011100101101111001",
3118 => "111001011010001101001000",
3119 => "111100010001100110100111",
3120 => "111111000010001111010001",
3121 => "000001000100001000100011",
3122 => "000011100101001000011001",
3123 => "000111010100110010101010",
3124 => "001011011110001111110101",
3125 => "001110001010110000110010",
3126 => "001110101001000110101110",
3127 => "001101111101101100110110",
3128 => "001100111010110101101000",
3129 => "001011011010101111000100",
3130 => "001001000100011011011000",
3131 => "000101111101000111011001",
3132 => "000011100101100011111101",
3133 => "000010010011110111101011",
3134 => "000000100110110001111101",
3135 => "111111100000001000000101",
3136 => "000001010101001100111100",
3137 => "000100011111101111001011",
3138 => "000101101001100101101110",
3139 => "000101010110000010110000",
3140 => "000110100111101110000000",
3141 => "001001010011000000100110",
3142 => "001011001001110000110010",
3143 => "001011111110111111111110",
3144 => "001011101010001101011001",
3145 => "001010001001010010101011",
3146 => "001001001101010100011001",
3147 => "001001010010101110111101",
3148 => "001001110101011011111101",
3149 => "001010100000111110111010",
3150 => "001001101101111100001110",
3151 => "000111110100100001000010",
3152 => "000110011000100111001001",
3153 => "000011111000000111101100",
3154 => "000000111000010010000000",
3155 => "000000001111110100000010",
3156 => "111111101011100110000000",
3157 => "111011100001010000000010",
3158 => "110101101000010111010110",
3159 => "110011010001011000011100",
3160 => "110110110010100011101011",
3161 => "111011111111110010000010",
3162 => "111110011000000000110000",
3163 => "111111101011000100110011",
3164 => "000010010111100001110011",
3165 => "000101001101000100101011",
3166 => "000110111010011000010110",
3167 => "000111100011000010000010",
3168 => "000111001110101100111101",
3169 => "000110000010001111000001",
3170 => "000011110010011111001100",
3171 => "000000011000110001001000",
3172 => "111100001101101000100001",
3173 => "110111100010000011010010",
3174 => "110010101100000000001110",
3175 => "101111000110101000001010",
3176 => "101110000100010011001000",
3177 => "101111001111001010001000",
3178 => "110001111110111011100000",
3179 => "110101100100001110011010",
3180 => "111000101101001101011000",
3181 => "111011111001001101000100",
3182 => "000000011111001111010001",
3183 => "000101100010001001101110",
3184 => "001000111110100100110100",
3185 => "001001100000111101101000",
3186 => "000111001100001110010100",
3187 => "000011100001011001000010",
3188 => "111111101001000100111101",
3189 => "111100010011101011111111",
3190 => "111010000001100011011000",
3191 => "110111010010011010110111",
3192 => "110011110000100100010100",
3193 => "110010010110110011110010",
3194 => "110100000110111100111100",
3195 => "110111010010010000011101",
3196 => "111010111110111110111110",
3197 => "111110011001100010001101",
3198 => "000000010111011101000011",
3199 => "000001001101111001001001",
3200 => "000010000110011110101101",
3201 => "000011011110011011000111",
3202 => "000101000100011101010111",
3203 => "000110000010101010001010",
3204 => "000101110010100010000111",
3205 => "000101000101110000010110",
3206 => "000100110110111010110010",
3207 => "000100110100010100000010",
3208 => "000100111110010110011110",
3209 => "000101010010011110010001",
3210 => "000100001000111010000001",
3211 => "000001001000101000110101",
3212 => "111110010011001010001010",
3213 => "111100011100011010111010",
3214 => "111010111000100100111100",
3215 => "111001011100101101110100",
3216 => "111000000100110110001111",
3217 => "110111010101101010001000",
3218 => "111000011110110011110110",
3219 => "111010111100101011001101",
3220 => "111101000111110011001100",
3221 => "111111001100000100101110",
3222 => "000001111011011001110100",
3223 => "000100110111110000011100",
3224 => "000111011000111000010110",
3225 => "001001001100110011001100",
3226 => "001010000100110000000110",
3227 => "001001110000001110010010",
3228 => "000111011001101001100100",
3229 => "000011001000110011110011",
3230 => "111111010011000000011000",
3231 => "111100101101100011001110",
3232 => "111001001110110011100001",
3233 => "110100011001101000010001",
3234 => "110000110000011011111010",
3235 => "101111101111000000110100",
3236 => "110000010100011000011110",
3237 => "110001100110100000111100",
3238 => "110011101000100001001100",
3239 => "110101110111010101101010",
3240 => "110111100011000000100001",
3241 => "111001001101111100100000",
3242 => "111011110001000001110111",
3243 => "111111000111000110111111",
3244 => "000001111100011101011010",
3245 => "000010100101000010001110",
3246 => "000001011100101101010010",
3247 => "000000100100110010010111",
3248 => "111111111111000001111100",
3249 => "111110010101100111001110",
3250 => "111011010011010010001011",
3251 => "110110111111101110001001",
3252 => "110010001100110000011000",
3253 => "101110101011100000001100",
3254 => "101101001000010100111000",
3255 => "101100110111010100000100",
3256 => "101101101010111111011000",
3257 => "101111011010110001100000",
3258 => "110001001011010001010100",
3259 => "110011010100101101111110",
3260 => "110111110101100100010000",
3261 => "111101111011101100000000",
3262 => "000001110011001001001100",
3263 => "000010100001100100000100",
3264 => "000010110111101000000000",
3265 => "000100000011010001100101",
3266 => "000100110000010111001001",
3267 => "000100010011100010000111",
3268 => "000011101001111111011001",
3269 => "000011011110101100101001",
3270 => "000010100101111010100110",
3271 => "111111111000110001101100",
3272 => "111100111001001110110100",
3273 => "111011011100001011000110",
3274 => "111010100010100010111110",
3275 => "111001000001100111101100",
3276 => "111000101010110101101100",
3277 => "111011010110010010111110",
3278 => "111111101010001000010011",
3279 => "000011001000111110010000",
3280 => "000101101010010010100011",
3281 => "001000101101001001111110",
3282 => "001100110111000110101010",
3283 => "010000110001000001110010",
3284 => "010010011100111100010100",
3285 => "010001110101100011110100",
3286 => "010000100010000110010110",
3287 => "001111010110111010011110",
3288 => "001101110010000101111000",
3289 => "001011000001100111110010",
3290 => "000111001101110111101011",
3291 => "000011111010100000100011",
3292 => "000010010101101000010000",
3293 => "000010000100101011110000",
3294 => "000010101011011001010001",
3295 => "000100011101000100111001",
3296 => "000111001000011110111011",
3297 => "001001011010111011010001",
3298 => "001010100010001001000100",
3299 => "001011001101100111000110",
3300 => "001011111111010000001010",
3301 => "001100101100101110010110",
3302 => "001101111101010010110100",
3303 => "001111000010010010110010",
3304 => "001101011000010000101100",
3305 => "001001101001010111010000",
3306 => "000111100100100100001110",
3307 => "001000001010100001110110",
3308 => "001000100010100001011110",
3309 => "000101100111100011110110",
3310 => "111111101101001001111110",
3311 => "111010010110101101101000",
3312 => "111000101111000011111011",
3313 => "111010110000101111010010",
3314 => "111101001110010000110101",
3315 => "111101101111001010000111",
3316 => "111101100110101001111100",
3317 => "111110001101001011010011",
3318 => "111111001100001010010011",
3319 => "000000110000001000110100",
3320 => "000010010000101001100011",
3321 => "000010011111101100000110",
3322 => "000010011111010101011010",
3323 => "000010101011110100110010",
3324 => "000001100011100001101000",
3325 => "111111100001010100110000",
3326 => "111110000001010011101000",
3327 => "111100001101011101111000",
3328 => "111001100011000000111000",
3329 => "111000000111101101100001",
3330 => "111000101000001011001101",
3331 => "111000100000010111100010",
3332 => "110110110000100111001101",
3333 => "110101001110110100100010",
3334 => "110101011000111000111000",
3335 => "111000001001000000110010",
3336 => "111100111011110101111000",
3337 => "000000110110000001000010",
3338 => "000010011011010111100111",
3339 => "000010110101101000010100",
3340 => "000010110011100100010111",
3341 => "000010010001000010011100",
3342 => "000001011001000111001001",
3343 => "000000101010011010011101",
3344 => "111111101111010000010011",
3345 => "111101110010010100001010",
3346 => "111100010000110110100010",
3347 => "111100110100100111110000",
3348 => "111101111001010000000111",
3349 => "111110011011001011100010",
3350 => "111111011100011111001100",
3351 => "000000100111010001001100",
3352 => "000000110111011011110011",
3353 => "000000101101001001110001",
3354 => "000001101110001110011111",
3355 => "000100011111000010100001",
3356 => "000111000011110111100100",
3357 => "000111101000111000010100",
3358 => "000111000110010001011110",
3359 => "000111001111010101000010",
3360 => "001000100110010110010000",
3361 => "001001111100110001000110",
3362 => "001010101000011010011000",
3363 => "001100000000011000111100",
3364 => "001101101010010010011010",
3365 => "001101110000100111001100",
3366 => "001101001001110100000000",
3367 => "001100011010101110011110",
3368 => "001010001100101011100101",
3369 => "000110100101000011110010",
3370 => "000010011001001011111110",
3371 => "111110110101010111000011",
3372 => "111101100010010110011001",
3373 => "111101010110111110110011",
3374 => "111100100101001100001101",
3375 => "111100101011110101000011",
3376 => "111111000010000101100101",
3377 => "000010101100001011010001",
3378 => "000110001100011101111000",
3379 => "001000101110111000101010",
3380 => "001010100010101010101111",
3381 => "001011100001011010100010",
3382 => "001011000100011110100111",
3383 => "001001111001111100111011",
3384 => "001000011111111111101100",
3385 => "000101110110001110101010",
3386 => "000001110011100111100001",
3387 => "111101100110101011001011",
3388 => "111010101110101100101001",
3389 => "111001110001010111101010",
3390 => "111001001010101000100010",
3391 => "110111010111010101101011",
3392 => "110101010001111001010110",
3393 => "110100001111101110101101",
3394 => "110100001001101011110111",
3395 => "110100011000011101110000",
3396 => "110100110110101100111110",
3397 => "110101111000011110001110",
3398 => "110111000010000010100111",
3399 => "110111011001110010110110",
3400 => "110111100100111010111010",
3401 => "111000111110100101101101",
3402 => "111011000100000001010100",
3403 => "111011101000011111101010",
3404 => "111010010110100101011001",
3405 => "111001001000101110111011",
3406 => "111000100000101101110010",
3407 => "110111010001001011011100",
3408 => "110101001001010101100110",
3409 => "110010100111111110110110",
3410 => "101111111100000100110000",
3411 => "101101100010111100111000",
3412 => "101100011101101011110100",
3413 => "101101111000000001000010",
3414 => "110001000010010101110100",
3415 => "110011000001111010000010",
3416 => "110010111111100101010110",
3417 => "110011011001010111100010",
3418 => "110101111010111110000010",
3419 => "111001010100101011100100",
3420 => "111011101000111111101100",
3421 => "111100111011001100110001",
3422 => "111110110010001110110101",
3423 => "000001010000001011100000",
3424 => "000010010100111011011111",
3425 => "000001010010111101010001",
3426 => "111111111100011011001010",
3427 => "111111100011101010110101",
3428 => "111111000111011111101110",
3429 => "111101111110101101000001",
3430 => "111101101110011100000000",
3431 => "111110111111111010100100",
3432 => "111111111111001111100010",
3433 => "000000000100011000011100",
3434 => "000001000000100111111100",
3435 => "000011101101001110011101",
3436 => "000110010111101111110001",
3437 => "000110111000000000011011",
3438 => "000110001001101101011001",
3439 => "000110110100001001000010",
3440 => "001000111100111000010100",
3441 => "001010110001101111001111",
3442 => "001011110100000000111001",
3443 => "001100101000011000111100",
3444 => "001101010110100101111110",
3445 => "001101110101001101110000",
3446 => "001110000000000011111110",
3447 => "001101101011111100010000",
3448 => "001100110000011111001000",
3449 => "001011000011101010100010",
3450 => "001000111011110100011010",
3451 => "000111110100101100101011",
3452 => "001000000010010000001110",
3453 => "000111111111110010101000",
3454 => "000111001110100001100011",
3455 => "000110100110010110110100",
3456 => "000110001100100010110000",
3457 => "000101101101101010100100",
3458 => "000101011100101101010010",
3459 => "000101001100001010100001",
3460 => "000011100011100100111001",
3461 => "111111110010100000110001",
3462 => "111011010100011001101110",
3463 => "111001000011000000010001",
3464 => "111010011111111010110011",
3465 => "111101010110011000101111",
3466 => "111110011110110011100100",
3467 => "111110101000001000111100",
3468 => "111111111101010111100101",
3469 => "000001011111011001001111",
3470 => "000001000010000011110100",
3471 => "111111001101010011000001",
3472 => "111110000111011110101110",
3473 => "111110000100110110000100",
3474 => "111101011010110000111000",
3475 => "111010100100101011001001",
3476 => "110110011110011111010100",
3477 => "110011011111001010011010",
3478 => "110010000111001101011000",
3479 => "110001010111100000010110",
3480 => "110000111010101011100110",
3481 => "110001011101110010111100",
3482 => "110010110101110100111100",
3483 => "110011011101101011000010",
3484 => "110011111101010100111110",
3485 => "110110011000100010110110",
3486 => "111010001010101010100001",
3487 => "111110000000010111011010",
3488 => "000000111001110111100100",
3489 => "000001000100101100100000",
3490 => "111111000000110101001010",
3491 => "111101010010010100000100",
3492 => "111100000101000010111010",
3493 => "111010010001100111001010",
3494 => "111000010110100100010000",
3495 => "110110011001000001011100",
3496 => "110100000000100010101000",
3497 => "110011000000101000110110",
3498 => "110100110100001101000010",
3499 => "111000001000011111110011",
3500 => "111011110001101010111111",
3501 => "111111011011110010010000",
3502 => "000010001111111000011000",
3503 => "000011101100000001101001",
3504 => "000100011011101101011000",
3505 => "000101001000010001110000",
3506 => "000101111000111010010010",
3507 => "000110011101111000100010",
3508 => "000101101011100101100011",
3509 => "000011110100101000000001",
3510 => "000011001011001000110010",
3511 => "000011110001111110000010",
3512 => "000100110011001111110010",
3513 => "000110011111010110101101",
3514 => "000111110100101111011110",
3515 => "001000101110100101111000",
3516 => "001010100010110101010100",
3517 => "001100100101010101010000",
3518 => "001110000000011100000110",
3519 => "001111000011000001000000",
3520 => "001111010100111000001100",
3521 => "001111001011010010001000",
3522 => "001111010110100111001100",
3523 => "001110101011111011110010",
3524 => "001100011111110101110000",
3525 => "001010001100110001000001",
3526 => "000111100100111001100100",
3527 => "000100001010101101111100",
3528 => "000010001110011111000110",
3529 => "000010000110001110100010",
3530 => "000001101100010110011111",
3531 => "000000111111001011001001",
3532 => "000000111010001100011100",
3533 => "000001100110001000010001",
3534 => "000010110001001000000101",
3535 => "000011100111100000101011",
3536 => "000011111110100010000101",
3537 => "000100101011001101100111",
3538 => "000101011111100101011110",
3539 => "000101010000110110100000",
3540 => "000100010011010011100110",
3541 => "000011000111110110000111",
3542 => "000000110100100011000101",
3543 => "111101110101100110110011",
3544 => "111011111000001001001010",
3545 => "111011011101110100111001",
3546 => "111011111111100001010110",
3547 => "111011111100001001110001",
3548 => "111010011111000100000000",
3549 => "111000011111111111100101",
3550 => "110110110010111101111100",
3551 => "110101011010010000001000",
3552 => "110011111001000000011010",
3553 => "110010001100000111010100",
3554 => "110000101010001011101000",
3555 => "101111001111000011011000",
3556 => "101110101001000011001000",
3557 => "101111111010000000101000",
3558 => "110010101011011100011110",
3559 => "110101101101110100110000",
3560 => "110111101011100000011001",
3561 => "111000110010100010100110",
3562 => "111010011111010100011111",
3563 => "111100100001100010000101",
3564 => "111101100101000010100110",
3565 => "111101001011010011101001",
3566 => "111011001101001111110100",
3567 => "111000000100110100010000",
3568 => "110101001110001101101110",
3569 => "110011101011000110110000",
3570 => "110011001100110111100010",
3571 => "110011101110000001101010",
3572 => "110101010001100000010100",
3573 => "110111011011111111110101",
3574 => "111001110001000001000110",
3575 => "111011101000011011001110",
3576 => "111101010100101100100101",
3577 => "000000000000101100111001",
3578 => "000011011000110111011110",
3579 => "000110010101011000010100",
3580 => "001000011000010010000110",
3581 => "001001111000000000010110",
3582 => "001011101000111011110011",
3583 => "001101001110100010011100",
3584 => "001101110101100001000110",
3585 => "001110010100101111100110",
3586 => "001111011111001110001010",
3587 => "010000000111001001110000",
3588 => "001110100010011100111000",
3589 => "001011111101010101101110",
3590 => "001010111111001110100110",
3591 => "001011010011011110000001",
3592 => "001011000101111110111111",
3593 => "001010000010011111100111",
3594 => "001000111001100111011011",
3595 => "001001000101010101000100",
3596 => "001011010001100111100010",
3597 => "001110000010000011101010",
3598 => "001111110100100111100110",
3599 => "010001001110001101000000",
3600 => "010011001100111111011000",
3601 => "010100111110100100101010",
3602 => "010101011111010011100110",
3603 => "010101000000000110100010",
3604 => "010100010110111011101100",
3605 => "010011101110001000101010",
3606 => "010001111011101000101110",
3607 => "001110100001110101000000",
3608 => "001011010100111110001010",
3609 => "001001001101110001101000",
3610 => "000110001001000011001100",
3611 => "000000100100000111111110",
3612 => "111001110111111100000001",
3613 => "110100100011011111111111",
3614 => "110010100101101110000110",
3615 => "110100001010111110000001",
3616 => "110110101000110011010001",
3617 => "111000100111101110111110",
3618 => "111100001010000011011000",
3619 => "000000110110001111010111",
3620 => "000011010000001010111001",
3621 => "000010110010100010101011",
3622 => "000010001011000101111111",
3623 => "000011001011010110000010",
3624 => "000011111001111011111010",
3625 => "000001011001100010000011",
3626 => "111100001001000000011001",
3627 => "110110011110001010101110",
3628 => "110001010100011110010000",
3629 => "101101001100000011000010",
3630 => "101010111111110010111010",
3631 => "101010101000001001010100",
3632 => "101010011111101000000100",
3633 => "101010000101010000100010",
3634 => "101010111110100001001110",
3635 => "101101100110011001110100",
3636 => "110000101110101101000000",
3637 => "110100011001100001000110",
3638 => "111000010110111100111001",
3639 => "111010001100000011110110",
3640 => "111001011000000110110010",
3641 => "111001000011010100010111",
3642 => "111010101110001101110100",
3643 => "111011111000111000010011",
3644 => "111010011010011001100100",
3645 => "110111100011111111110101",
3646 => "110101011110110111000111",
3647 => "110100100000110010111000",
3648 => "110100110100010111011010",
3649 => "110110100111011001110101",
3650 => "111000000110011100010101",
3651 => "111000011011111111010101",
3652 => "111001011010100011100010",
3653 => "111010111000011100001001",
3654 => "111011001101111001111001",
3655 => "111011011101011001010101",
3656 => "111101100101011101100011",
3657 => "000001000110101000001101",
3658 => "000011101001010100010101",
3659 => "000100010010010011000110",
3660 => "000100100100011111110100",
3661 => "000101101011101001111000",
3662 => "000111001001100010010010",
3663 => "001000011010000010001001",
3664 => "001001011101100001000100",
3665 => "001001111110100001001100",
3666 => "001001100110000100100000",
3667 => "001001011001111001111000",
3668 => "001010000010100011110010",
3669 => "001010000011010111110100",
3670 => "001001100100110000010110",
3671 => "001010101100011010000110",
3672 => "001100110010101000001000",
3673 => "001101100011101100110000",
3674 => "001101011001100111110100",
3675 => "001101110011101010100000",
3676 => "001110100001110111111100",
3677 => "001111001101001111111000",
3678 => "001111110010110010101110",
3679 => "001111100000101011011100",
3680 => "001101110010011100101100",
3681 => "001010100001110001110101",
3682 => "000110011010100011000001",
3683 => "000010110100100110111010",
3684 => "111111110010001010000010",
3685 => "111100111001100011111111",
3686 => "111010110011001110101110",
3687 => "111001101011000111000100",
3688 => "111001010111010111000100",
3689 => "111010000011010011011010",
3690 => "111011011000011101101100",
3691 => "111100100100110011001100",
3692 => "111101010110001011100000",
3693 => "111101110111000000011011",
3694 => "111110000011110000011000",
3695 => "111110001000111010110111",
3696 => "111110001110101010100010",
3697 => "111101010011001011110111",
3698 => "111011000101110100001110",
3699 => "111001000111011100100100",
3700 => "111000010001001001100110",
3701 => "110111111100100101001100",
3702 => "110111001000001001011000",
3703 => "110101001110101000100100",
3704 => "110010011000111011100100",
3705 => "101111001101000100111000",
3706 => "101100000011010001100100",
3707 => "101000111100001111010010",
3708 => "100110100110101000101001",
3709 => "100101101100010101100011",
3710 => "100101110111000011100010",
3711 => "100111100011011000101001",
3712 => "101010111000010010010110",
3713 => "101110011001110111001000",
3714 => "110010000010101001000110",
3715 => "110110001111111001010110",
3716 => "111001111001000101110101",
3717 => "111100101111100000111100",
3718 => "111111011111000101011111",
3719 => "000000111010100000000011",
3720 => "111111111100101001000001",
3721 => "111101111110110101010111",
3722 => "111100001000100100001111",
3723 => "111010010101100010000001",
3724 => "111000101110110010111000",
3725 => "110110111011110011011101",
3726 => "110101000110000100010001",
3727 => "110100100010110001010110",
3728 => "110101111100000001010011",
3729 => "111001001100010111110100",
3730 => "111101000000001100101111",
3731 => "111111111111100000110010",
3732 => "000011010010011111111100",
3733 => "000111101101000011000110",
3734 => "001100001000000111110110",
3735 => "001111111111001101101000",
3736 => "010011001100100000010100",
3737 => "010101101110100000000110",
3738 => "010111011101000100000100",
3739 => "011000000000001101000001",
3740 => "010111111110001011001100",
3741 => "010111011001011010100100",
3742 => "010100110100110111110000",
3743 => "010001000001011101001010",
3744 => "001110100010010010101110",
3745 => "001100111101000001100010",
3746 => "001010110100010000101101",
3747 => "001001011111111001111010",
3748 => "001001110110110001010000",
3749 => "001010001101110011000110",
3750 => "001010010101000000011000",
3751 => "001100001000110011000000",
3752 => "001111101101101100000010",
3753 => "010010010110000111111100",
3754 => "010011010000000110111000",
3755 => "010100010111101101100110",
3756 => "010101101110000000111010",
3757 => "010110000100101101010110",
3758 => "010100110110010011101010",
3759 => "010000100000111000101110",
3760 => "001001000011101101100111",
3761 => "000010000110101010101111",
3762 => "111111010111011110110001",
3763 => "000000000100011001111101",
3764 => "111111010101101101001111",
3765 => "111011111110101011111111",
3766 => "111010000110011001010111",
3767 => "111010100011011110001011",
3768 => "111010011001010011100111",
3769 => "111001010100110100101010",
3770 => "111001100111011010110110",
3771 => "111011110011111000000010",
3772 => "111101000101001100100011",
3773 => "111011011100010011000010",
3774 => "111001001100110011001010",
3775 => "111000001011011101111110",
3776 => "110111001011011011010001",
3777 => "110110010110011000111110",
3778 => "110110010101010010011010",
3779 => "110101011000100000000110",
3780 => "110011011101001110110100",
3781 => "110010101011010000101010",
3782 => "110010100011011000011110",
3783 => "110001110011111110101010",
3784 => "110001110001110101000010",
3785 => "110011110111000110110000",
3786 => "110110101001010010011111",
3787 => "110111110001010001000000",
3788 => "110111110010101011010000",
3789 => "111000001010010110101100",
3790 => "110111111100100011001010",
3791 => "110110110010101110001101",
3792 => "110101010111001101111011",
3793 => "110011101100111111001000",
3794 => "110010111100011011010110",
3795 => "110011101111111000011010",
3796 => "110101010001101010101010",
3797 => "110111101101100001001011",
3798 => "111011011100110110111100",
3799 => "111111110101000100100101",
3800 => "000011101110101100110111",
3801 => "000110001110111110001011",
3802 => "000111011110100000111111",
3803 => "000111111100101010110010",
3804 => "001000001001010000101001",
3805 => "001000101011011011010001",
3806 => "001000011011011000010010",
3807 => "000101110101100110011100",
3808 => "000010100001000110000100",
3809 => "000000111111110101000101",
3810 => "000001001011011001001100",
3811 => "000010010101110111110101",
3812 => "000100010101111000111010",
3813 => "000110100010000111001111",
3814 => "001001001010110110011101",
3815 => "001100100000001001010110",
3816 => "001111001111000001000000",
3817 => "010001000110111011010010",
3818 => "010010101101010011110110",
3819 => "010011110101111000000010",
3820 => "010100011000110111101100",
3821 => "010011111110010000011110",
3822 => "010010111010101010101110",
3823 => "010010011111011111010110",
3824 => "010010001011010100010110",
3825 => "010000110010101101110100",
3826 => "001111010010001010010100",
3827 => "001111001110100101001010",
3828 => "010000001101001011100010",
3829 => "010000101001000110100010",
3830 => "010000000100100111100000",
3831 => "001110010011010101110110",
3832 => "001011000101011001010000",
3833 => "000111000011011100100000",
3834 => "000010001111100111101101",
3835 => "111100100100000010100011",
3836 => "110111011100101011010010",
3837 => "110100010110110101000011",
3838 => "110011010010001101011110",
3839 => "110011000010011010101010",
3840 => "110010101011001101111110",
3841 => "110010011010010000010010",
3842 => "110011000001001011111100",
3843 => "110101000011110101000100",
3844 => "111000000111010110101010",
3845 => "111011000110111011001000",
3846 => "111100101101100100000000",
3847 => "111100001000111100001111",
3848 => "111010011100011010100000",
3849 => "111000010101101000110000",
3850 => "110101011000011110101110",
3851 => "110001110110101000001110",
3852 => "101101111111111100100000",
3853 => "101010101000101011101100",
3854 => "101000101101011100011110",
3855 => "100111000011110000001001",
3856 => "100101000001111110001111",
3857 => "100011101110111001000111",
3858 => "100011101110111111001111",
3859 => "100100100001011110000101",
3860 => "100101001101010001000010",
3861 => "100110000001110010000011",
3862 => "100111111010000100100000",
3863 => "101010100100000011111100",
3864 => "101100111100101111100110",
3865 => "101110111011001101111000",
3866 => "110001110001001101110100",
3867 => "110101110011110001110010",
3868 => "111001111110110010010001",
3869 => "111101111111010010100101",
3870 => "000001000001111100110110",
3871 => "000001110101110101110011",
3872 => "000000111110101010001101",
3873 => "111111011010010100101000",
3874 => "111100101000011101110110",
3875 => "111000110101000100010110",
3876 => "110110111100000100101100",
3877 => "110111111010101011000010",
3878 => "111000111111100101000011",
3879 => "111001111001110011100100",
3880 => "111011111111000100010100",
3881 => "111110101111111010101111",
3882 => "000001110111101100000111",
3883 => "000101010000110001000110",
3884 => "001001011100001010101011",
3885 => "001110010101110000111000",
3886 => "010001110110110010000010",
3887 => "010011101011010000011110",
3888 => "010101001000010101010100",
3889 => "010110101001110011001100",
3890 => "011000000101010001011011",
3891 => "011000101001101000110011",
3892 => "011000011111000001110001",
3893 => "010111110100101110111010",
3894 => "010101101000011010010100",
3895 => "010010101001011000110100",
3896 => "010000101000101010011110",
3897 => "001110100000111001101000",
3898 => "001011001010101101111000",
3899 => "001001000111001000100100",
3900 => "001000111010000001011011",
3901 => "000111010101100101001100",
3902 => "000101001001101011110100",
3903 => "000101001110001010110100",
3904 => "000111001001110101101100",
3905 => "001001011001001101001110",
3906 => "001001011010010011000011",
3907 => "000110001000101001101010",
3908 => "000010000011111010101001",
3909 => "000000001001010000011010",
3910 => "000010010001101111110010",
3911 => "000101110011101010000011",
3912 => "000101111011110001110100",
3913 => "000011110100011110100001",
3914 => "000010111010000000000101",
3915 => "000010111011011011101011",
3916 => "000001110000010011101110",
3917 => "111110100110011010011000",
3918 => "111010111110111100000111",
3919 => "111000000000001101110000",
3920 => "110100110011001001111100",
3921 => "110000011101111101101010",
3922 => "101100000110001000001100",
3923 => "101000111010111010100100",
3924 => "100110000001111110100001",
3925 => "100100011001101001010011",
3926 => "100110001000010111000000",
3927 => "101001111000000010100100",
3928 => "101110000111001111110010",
3929 => "110010001101010011000010",
3930 => "110101101011100101010100",
3931 => "111001001101011110111000",
3932 => "111100110011011111011001",
3933 => "000000000000001110110010",
3934 => "000001010110010010100010",
3935 => "111111011000101110100100",
3936 => "111100001011111110111101",
3937 => "111001101111111111100000",
3938 => "110111011111110111101110",
3939 => "110100110100000100111011",
3940 => "110010010101110110110110",
3941 => "110001010010110010110110",
3942 => "110001001111000010110000",
3943 => "110001101100101000110100",
3944 => "110011000011100101010100",
3945 => "110101000000100011000000",
3946 => "111000001111011111110001",
3947 => "111100101110001001011111",
3948 => "000000101100110100100000",
3949 => "000011101110111110101101",
3950 => "000110111100011110100100",
3951 => "001011100101010001001000",
3952 => "010000001011011100101100",
3953 => "010010011100101000100100",
3954 => "010010100111001110101100",
3955 => "010001001001000011101110",
3956 => "001111100101111100000100",
3957 => "001110111101011110011000",
3958 => "001101101000011010101000",
3959 => "001100010001100001100110",
3960 => "001011101010111101100000",
3961 => "001010100101010011011010",
3962 => "001001110100110100111010",
3963 => "001010101001011010101110",
3964 => "001100011011110110101000",
3965 => "001110001110111010010010",
3966 => "010000011110000001000000",
3967 => "010011011011010001101000",
3968 => "010101100011111010110000",
3969 => "010110100001101101110100",
3970 => "010111001111010111010100",
3971 => "010111111110011100101100",
3972 => "011000001000110001100010",
3973 => "010111001001001111011010",
3974 => "010110111110100110000000",
3975 => "011000000100000010001110",
3976 => "011000000001111001110111",
3977 => "010111010110101111000000",
3978 => "010110101001100010000000",
3979 => "010101011001100010011110",
3980 => "010011110100011111010000",
3981 => "010000101110100011110100",
3982 => "001011010100111101110000",
3983 => "000011111000001000101111",
3984 => "111011010000111101000011",
3985 => "110011011011101111011110",
3986 => "101101100000100011000010",
3987 => "101010100100011011011010",
3988 => "101010011101110100110000",
3989 => "101011011100100011001010",
3990 => "101101011100100011101110",
3991 => "110000101111010001010100",
3992 => "110101011001000000001100",
3993 => "111011001111100100100110",
3994 => "000000011110101110110001",
3995 => "000011010101101000001101",
3996 => "000011000010011110011001",
3997 => "000000011000100010000000",
3998 => "111100110010111010100111",
3999 => "111000110100110001100111",
4000 => "110100101111011101100111",
4001 => "110000000000011000101010",
4002 => "101011011111110101000000",
4003 => "101000110010011111010000",
4004 => "100110111100100000111001",
4005 => "100101111001111111100101",
4006 => "100101100100010100000111",
4007 => "100100110001010100000111",
4008 => "100100110101101100101001",
4009 => "100110100111101001110101",
4010 => "101000110101110010111010",
4011 => "101010101001011011111010",
4012 => "101101000111110101100000",
4013 => "110001101010011000101000",
4014 => "110110100111110111001101",
4015 => "111011100010001101101100",
4016 => "000001101101100110000110",
4017 => "000111001111000011100011",
4018 => "001011000010100011101101",
4019 => "001101111110000100111010",
4020 => "001110101110111010000110",
4021 => "001100001100001111100010",
4022 => "001000000001110111011110",
4023 => "000100100010011111101011",
4024 => "000001010011001010010001",
4025 => "111101111111101101001001",
4026 => "111100101001101011100100",
4027 => "111101101011111010101111",
4028 => "111111101010011010110001",
4029 => "000001000110100101101010",
4030 => "000010001011011101110000",
4031 => "000100011111110011000010",
4032 => "000111111001100111111011",
4033 => "001100001110101010010010",
4034 => "010000110001010100010100",
4035 => "010011010101110011000100",
4036 => "010101000101111011000100",
4037 => "010111100100000000011100",
4038 => "011001011000110001100001",
4039 => "011001101111001110001101",
4040 => "011000111010010110001001",
4041 => "010111110001100000100110",
4042 => "010110100110101011101100",
4043 => "010100110100100000101000",
4044 => "010001111100010000000000",
4045 => "001110000010000001000110",
4046 => "001010011100000010101110",
4047 => "000110111100000100111010",
4048 => "000010100111110010110000",
4049 => "111111100001001010010001",
4050 => "111110101101001101000101",
4051 => "111110010100111110011010",
4052 => "111011110111101000011101",
4053 => "110111010111111000110011",
4054 => "110100001100101001001010",
4055 => "110011010101011011001000",
4056 => "110100010000110111010010",
4057 => "110111101011000110011101",
4058 => "111011101001010110011111",
4059 => "111110000110100110011100",
4060 => "111111110000110010111111",
4061 => "000001010110100110100110",
4062 => "000010100111010100101111",
4063 => "000010101101110110100000",
4064 => "000000101111011010110000",
4065 => "111100100110010110111000",
4066 => "110111111100000100011100",
4067 => "110011010000101001100100",
4068 => "101100100011101011000100",
4069 => "100101010110100111110011",
4070 => "100001101110101001101001",
4071 => "100001101001100011110111",
4072 => "100010010100101110000001",
4073 => "100010110000001010010111",
4074 => "100011111010110010110101",
4075 => "100101000111001010111011",
4076 => "100110000111011100000101",
4077 => "101001111100110010010100",
4078 => "110000011001010111111110",
4079 => "110110110010011110110110",
4080 => "111100101001111111101010",
4081 => "000000110000110001101000",
4082 => "000010001101111101000010",
4083 => "000001111111111111000101",
4084 => "000000101010101100001110",
4085 => "111101110110110001110111",
4086 => "111001001101001111101010",
4087 => "110100100000100010110100",
4088 => "110001100101110110000000",
4089 => "101111110101101001001100",
4090 => "101111001100000011111010",
4091 => "110000101001001001111100",
4092 => "110011111111010110011110",
4093 => "110111010101010010101101",
4094 => "111001101011111111100110",
4095 => "111100010110110001010110",
4096 => "111111110101010011111101",
4097 => "000011011101010101110010",
4098 => "000110111011100011101110",
4099 => "001010100010101101100111",
4100 => "001110011101001100111110",
4101 => "010000110011011101010110",
4102 => "010000111100010000000000",
4103 => "010000111001001010011010",
4104 => "010001001001110000100010",
4105 => "010001010111010110010000",
4106 => "010000111101111000111000",
4107 => "001110111110000101101010",
4108 => "001100100010010000100110",
4109 => "001011010001110110111001",
4110 => "001010110001001100111111",
4111 => "001010001110101010101110",
4112 => "001010010111000110011110",
4113 => "001011110001100110101000",
4114 => "001101011010001011100110",
4115 => "001110100000111111111000",
4116 => "001111001010011011110000",
4117 => "001111111001101000000000",
4118 => "010001010111011100111110",
4119 => "010010011100110011100010",
4120 => "010010101000101101010000",
4121 => "010010111000101101101100",
4122 => "010010110000000010011010",
4123 => "010001101111010101001010",
4124 => "010000101111001000101010",
4125 => "010000100111010111101010",
4126 => "010000100001111101100000",
4127 => "001110100100010000111010",
4128 => "001010111110101001110010",
4129 => "000110101101000011111100",
4130 => "000000001111001111010011",
4131 => "110110101000000000001100",
4132 => "101100111001100110010110",
4133 => "100110101000111000110000",
4134 => "100011011110000110000001",
4135 => "100001111111100001101010",
4136 => "100001111011010101000001",
4137 => "100011010101001100000001",
4138 => "100111111001000111110111",
4139 => "101111011011111011101100",
4140 => "110110110111111000010101",
4141 => "111101001000100011101010",
4142 => "000001100001000011011001",
4143 => "000010011110010000011010",
4144 => "000000101010010011100000",
4145 => "111101101000010011011000",
4146 => "111001100101010011101011",
4147 => "110100011010011001101110",
4148 => "101111011110110101100000",
4149 => "101100001001110011100100",
4150 => "101001110110000000000110",
4151 => "100111110111100111000011",
4152 => "100110101010110001100010",
4153 => "100110110010010110100111",
4154 => "100111110001110010110101",
4155 => "101000100110000001010100",
4156 => "101001001100000101101100",
4157 => "101010101111001111110110",
4158 => "101110010010101010111010",
4159 => "110010110111101001110110",
4160 => "110111011010110110000111",
4161 => "111101000100001110110011",
4162 => "000011101101111101100000",
4163 => "001010001111011110000100",
4164 => "010000010010100000010010",
4165 => "010100100001111100011110",
4166 => "010110000100001111110110",
4167 => "010101001100100101000010",
4168 => "010010110000000110001010",
4169 => "001111110101011101011110",
4170 => "001100011110100101100110",
4171 => "001001011100100000100010",
4172 => "000111101101111111100111",
4173 => "000110010111010001001110",
4174 => "000101011000001111100110",
4175 => "000101101010100101111101",
4176 => "000110101011001110111010",
4177 => "000111100010010101001110",
4178 => "001000100111111101000011",
4179 => "001010110101011111010110",
4180 => "001110000110100111001010",
4181 => "010010000001010110000000",
4182 => "010110001000110001110000",
4183 => "011001110101101101100101",
4184 => "011100001110110100111101",
4185 => "011100010000100011110111",
4186 => "011011001001000110011101",
4187 => "011010011010011011001110",
4188 => "011001101010101100010011",
4189 => "011000100101101001111011",
4190 => "010110001110100000110000",
4191 => "010010111000100001011000",
4192 => "001111011000111100111010",
4193 => "001010000111101111110111",
4194 => "000100011111111110010011",
4195 => "000001010111011000011101",
4196 => "000000000010101110000110",
4197 => "111111001010010000000100",
4198 => "111101000011011101101101",
4199 => "111001110001111100110011",
4200 => "110110011100110011101001",
4201 => "110010101101011101100100",
4202 => "110000110111111101101010",
4203 => "110011000010110000000100",
4204 => "110111000111001010110001",
4205 => "111010100010101011101000",
4206 => "111100110101111001100001",
4207 => "111111010110111010111010",
4208 => "000001110110000011000100",
4209 => "000010111110110000100010",
4210 => "000011001010000011000001",
4211 => "000010001010100111100000",
4212 => "111111101010000101110110",
4213 => "111011001011110110100101",
4214 => "110100100101011000011101",
4215 => "101110011110100110110110",
4216 => "101010011000011000010110",
4217 => "100111001100101011011001",
4218 => "100100011110110100101111",
4219 => "100011001000010110000101",
4220 => "100011110001100011010001",
4221 => "100100111110110011001110",
4222 => "100110010111101100011100",
4223 => "101001100011110101000010",
4224 => "101110111000110101111100",
4225 => "110101010101010101101000",
4226 => "111011000001011000110001",
4227 => "111111110100101010101101",
4228 => "000101001000011111000000",
4229 => "001001111000110011000001",
4230 => "001100001000110111011000",
4231 => "001011010010111101100011",
4232 => "001000100111000000111101",
4233 => "000100111000010111100110",
4234 => "111111100011101111000111",
4235 => "111010101101101000011111",
4236 => "110111101010100100000000",
4237 => "110101101001010011000101",
4238 => "110101011111001101110000",
4239 => "110110111000101101001010",
4240 => "111001010000111011100010",
4241 => "111100011000111110111001",
4242 => "111111001110010011111010",
4243 => "000010000010001011101100",
4244 => "000100110110111000001101",
4245 => "001000101100011001101111",
4246 => "001101101100000010100110",
4247 => "010000101011110100000100",
4248 => "010001111100011010001010",
4249 => "010010111001001101110010",
4250 => "010010111101000011111000",
4251 => "010010110101100101111110",
4252 => "010010011101000111110110",
4253 => "010001101000011000011000",
4254 => "010000000111001001111110",
4255 => "001101100111011011011110",
4256 => "001011101010110000110010",
4257 => "001001101110100001011110",
4258 => "000111110100000110101111",
4259 => "000111011111001000010101",
4260 => "000111101000100101111011",
4261 => "001000011100101000101110",
4262 => "001010010111010011001000",
4263 => "001011101100110100100010",
4264 => "001011101111100000001001",
4265 => "001010100010011100110000",
4266 => "001001011101110101110101",
4267 => "001001011011000000001000",
4268 => "001001010100100001110000",
4269 => "001000111010100100111100",
4270 => "001000100111100110010011",
4271 => "001000100100111011101100",
4272 => "000111101100010100010010",
4273 => "000101001000001100110111",
4274 => "000001110000001001001101",
4275 => "111100111100110000100111",
4276 => "110110011101110101110111",
4277 => "110000000100100001001110",
4278 => "101010110111011001110100",
4279 => "100110111110101101011111",
4280 => "100011110111000000010010",
4281 => "100010001101000110101001",
4282 => "100010111011100110101101",
4283 => "100101010110110001011011",
4284 => "101001100111010110111100",
4285 => "101111000101010000000000",
4286 => "110100010001011000010110",
4287 => "111000011110011110111110",
4288 => "111010110100100010011111",
4289 => "111011111101111100111000",
4290 => "111100011001001100010000",
4291 => "111011100011000101110010",
4292 => "111010001111001101000011",
4293 => "111000011000101111101100",
4294 => "110101010010100010100110",
4295 => "110001010010110100100010",
4296 => "101101011111011010101000",
4297 => "101010110000111110100100",
4298 => "101000010010001011000010",
4299 => "100110100010101011101110",
4300 => "100110111000011010101100",
4301 => "100111111000110111101111",
4302 => "101000100001100100110000",
4303 => "101001111111011110110000",
4304 => "101110001011001000100110",
4305 => "110101000010101000111110",
4306 => "111100001010111110011000",
4307 => "000010100010111010010111",
4308 => "001000010111110000010110",
4309 => "001101111000000000010110",
4310 => "010010101011101001011100",
4311 => "010100111011001111000000",
4312 => "010100101100110100010000",
4313 => "010011011101001011100010",
4314 => "010001010001001001101100",
4315 => "001110001111101111001110",
4316 => "001010111010110101110011",
4317 => "001000011011100000101010",
4318 => "000110110101001001010101",
4319 => "000101000110010010000000",
4320 => "000011110010111101011010",
4321 => "000010101001110111001001",
4322 => "000001010001011100111110",
4323 => "000001100111101110110001",
4324 => "000100100111010110001011",
4325 => "001000101100111100111101",
4326 => "001100001110000100011010",
4327 => "001111101110001101100000",
4328 => "010011101000110110100000",
4329 => "010110001000110011101110",
4330 => "010111110010101010110100",
4331 => "011001111011000101010111",
4332 => "011010001101001011111000",
4333 => "010111011101111011011100",
4334 => "010011101011010111011000",
4335 => "010000010000001011001010",
4336 => "001100101100101101110110",
4337 => "001000001110100001010100",
4338 => "000011111011000001010000",
4339 => "000001001111111000001100",
4340 => "111111100010101110011010",
4341 => "111101011001000110111111",
4342 => "111011010010010010001001",
4343 => "111011001110011010111110",
4344 => "111100101111101000000101",
4345 => "111100001011101110111011",
4346 => "111000100001001011110110",
4347 => "110100011111011101111100",
4348 => "110001000010010110001110",
4349 => "101110101001001111100110",
4350 => "101111101110001001100100",
4351 => "110011010100011011110110",
4352 => "110110011000001100000001",
4353 => "111000100110000001110011",
4354 => "111010100000110001010111",
4355 => "111100011100111000001110",
4356 => "111110000111100011110011",
4357 => "111110110110000011111011",
4358 => "111110110000100011111110",
4359 => "111101010000100010011000",
4360 => "111010011011111001010101",
4361 => "110111010111001001111110",
4362 => "110011111001011000010100",
4363 => "110000001111011011010010",
4364 => "101100111011011101010010",
4365 => "101010110010001011000010",
4366 => "101010000011001001110110",
4367 => "101001011001010110111100",
4368 => "101010010010000000001000",
4369 => "101101101011011001001100",
4370 => "110000101101100101011110",
4371 => "110100001001110000100100",
4372 => "111010100000010111101010",
4373 => "000010001111000001000100",
4374 => "001001000010100101000011",
4375 => "001101100100010110001010",
4376 => "001111110000010110011010",
4377 => "010000010010110010110100",
4378 => "001110101110011101000010",
4379 => "001011010110010010110000",
4380 => "000111011111101100100000",
4381 => "000011100000001010011011",
4382 => "111111011010101011110111",
4383 => "111011110111000100011111",
4384 => "111010001010100010010001",
4385 => "111011011110101010011100",
4386 => "111110101001000001000101",
4387 => "000001010111011101010010",
4388 => "000011000110010100010010",
4389 => "000100110001011100110111",
4390 => "000111101011000010100001",
4391 => "001011010110111111101010",
4392 => "001101110111001110100010",
4393 => "001111110011111010110010",
4394 => "010010000101010101111110",
4395 => "010010110110000101111010",
4396 => "010010011100111111001010",
4397 => "010011001100100000110000",
4398 => "010100101110001010001100",
4399 => "010101000100101100111100",
4400 => "010100000011010000011010",
4401 => "010011001110001001000110",
4402 => "010010000110011110001010",
4403 => "001111100001011011100100",
4404 => "001100111110010101101010",
4405 => "001011011001010011001110",
4406 => "001010101101111011001100",
4407 => "001010110111100000111111",
4408 => "001010110101000010000100",
4409 => "001010011011101000000010",
4410 => "001001100010010111110110",
4411 => "001000000000010000100110",
4412 => "000111000011111001000101",
4413 => "000110111111101100001100",
4414 => "000111101000101001101001",
4415 => "001000000000100101001000",
4416 => "000101110100000011010011",
4417 => "000001111000001111001101",
4418 => "111110100101111100111011",
4419 => "111011101011100111011000",
4420 => "111000001111000111011001",
4421 => "110100100100011101011110",
4422 => "110001101001110100010010",
4423 => "101111110100000000010100",
4424 => "101110110111100001111100",
4425 => "101111001100110010000010",
4426 => "110000101111000100110110",
4427 => "110010101110001011100100",
4428 => "110100011010001110011101",
4429 => "110101110000010000001110",
4430 => "110111101000110010100010",
4431 => "111001100101000010100000",
4432 => "111010001100100001111011",
4433 => "111001101000100110011011",
4434 => "111000010010110101100000",
4435 => "110110101110101100001110",
4436 => "110101110111101011100100",
4437 => "110100111111000110000011",
4438 => "110011100101010010111100",
4439 => "110010100011010101110010",
4440 => "110001000001001100000000",
4441 => "101110000111011010100000",
4442 => "101011101010010100111100",
4443 => "101010110010111001110100",
4444 => "101011000111011011011000",
4445 => "101100011111010110011010",
4446 => "101110000000010111110110",
4447 => "101111001001100100100100",
4448 => "110001101101000011000010",
4449 => "110110011010000000101100",
4450 => "111011000000111111110010",
4451 => "111110001000110101111000",
4452 => "000001000001011010010001",
4453 => "000100011100000011110110",
4454 => "000111010011010011101110",
4455 => "001001001100110010001010",
4456 => "001011000011011001001110",
4457 => "001100011010101000001000",
4458 => "001100000010100010100010",
4459 => "001010110011110111010001",
4460 => "001001101011101100001110",
4461 => "000111011111100011010000",
4462 => "000100000110111001100101",
4463 => "000001101011100001101001",
4464 => "000001001001000010001000",
4465 => "000001001000101101110001",
4466 => "000001010101001001001110",
4467 => "000010011110111011101100",
4468 => "000100010011100011111100",
4469 => "000111010011001111100110",
4470 => "001011100101101111010111",
4471 => "001111000010001010010000",
4472 => "010001100001111101011010",
4473 => "010011110101110110110010",
4474 => "010100000001011011110010",
4475 => "010001101100110101010010",
4476 => "001111000000111111110110",
4477 => "001100100011000100001000",
4478 => "001001010000111011111000",
4479 => "000101010000001000000001",
4480 => "000010011000011000111001",
4481 => "000001010010100100111101",
4482 => "000000100110000010111001",
4483 => "000000001011111100001011",
4484 => "000001000000001100100000",
4485 => "000010010010111000110100",
4486 => "000010110110010110010000",
4487 => "000010111111100110001100",
4488 => "000011000111011011101011",
4489 => "000010110111101110110110",
4490 => "000010001110100101111111",
4491 => "000000110110111100000111",
4492 => "111101101010100111001100",
4493 => "110111111011101111000001",
4494 => "110001001001001011011010",
4495 => "101100011100110001001000",
4496 => "101011000011111100100000",
4497 => "101100000001110111110110",
4498 => "101110001001110101000000",
4499 => "110000011001000000100000",
4500 => "110010011001000000100100",
4501 => "110100000001101001000101",
4502 => "110110000100011001000011",
4503 => "111001000110011110001010",
4504 => "111010111110110100100010",
4505 => "111010111101110101000111",
4506 => "111010101111111010010000",
4507 => "111010001111101101110110",
4508 => "111000011001010101111110",
4509 => "110101001111010010011101",
4510 => "110010100010001011000010",
4511 => "110001000010011100100100",
4512 => "101111100011100101111100",
4513 => "101111001010111110101100",
4514 => "110000001011100001010000",
4515 => "110000110101110111110100",
4516 => "110010010111110001000000",
4517 => "110101100111100111101110",
4518 => "111001010101101001011010",
4519 => "111100110101011100111001",
4520 => "111111111101011111010011",
4521 => "000011100101111011010111",
4522 => "000110111111011110111110",
4523 => "001000001110001110001001",
4524 => "001000000010101010110111",
4525 => "000111100010110011010111",
4526 => "000110100010111001111111",
4527 => "000100011111010100111010",
4528 => "000001110101001000000111",
4529 => "000000101110110011011100",
4530 => "000000111110110111111110",
4531 => "000000111010010011100111",
4532 => "000001011010110101101101",
4533 => "000010111101110101011101",
4534 => "000100100000110101110101",
4535 => "000101110000000110011111",
4536 => "000110100001110101110001",
4537 => "000111010011001111100111",
4538 => "001001011011001101011010",
4539 => "001100101010000110011010",
4540 => "001111011101101110111110",
4541 => "010001010110010000110010",
4542 => "010010001000101001000110",
4543 => "010010010000010110110000",
4544 => "010010110010001100011000",
4545 => "010011001100111000110000",
4546 => "010011000001100000001010",
4547 => "010010100001000010000110",
4548 => "010001011110010110001000",
4549 => "010000101001000100001000",
4550 => "001111111110111011110110",
4551 => "001110011011000100110110",
4552 => "001100101011110011110110",
4553 => "001011101100100000110111",
4554 => "001011100000111101010011",
4555 => "001011101010100101011101",
4556 => "001011011010001011011011",
4557 => "001010110011000110100111",
4558 => "001001010110110100110000",
4559 => "000110011101011000011000",
4560 => "000010010110001110001101",
4561 => "111101001011011000000010",
4562 => "111000001000011001101011",
4563 => "110100011000101111011011",
4564 => "110001011100101110100000",
4565 => "101111011000010011011100",
4566 => "101111010110011000001110",
4567 => "110001110010001111000110",
4568 => "110101100111110100110010",
4569 => "111001110011111010100010",
4570 => "111110010110010001110011",
4571 => "000010101000110001110010",
4572 => "000101011111011111010110",
4573 => "000110010110010110010100",
4574 => "000101001101111010101110",
4575 => "000010011101100011000000",
4576 => "111110000110000000010110",
4577 => "111001000010110011001001",
4578 => "110101110100100001111101",
4579 => "110100110100011111110011",
4580 => "110100010100010010011110",
4581 => "110100001101111110101011",
4582 => "110100110001111010111001",
4583 => "110100100100011011110011",
4584 => "110010110010001111010110",
4585 => "110000011110010101100000",
4586 => "101110110001011111101110",
4587 => "101101111000000011111010",
4588 => "101110000001101111001110",
4589 => "101111101001010110010100",
4590 => "110001111110000011000110",
4591 => "110100101011110110000111",
4592 => "111000100111110101101111",
4593 => "111100111001000001000000",
4594 => "000000110110011010100000",
4595 => "000101010110111011111100",
4596 => "001001010010110010100110",
4597 => "001011101100010111100111",
4598 => "001101000110110000001100",
4599 => "001100111111011100001100",
4600 => "001011110100110100001100",
4601 => "001010101110111110010101",
4602 => "001001000100111001111110",
4603 => "000111000011001010000100",
4604 => "000101010010010011010111",
4605 => "000011010011011111001000",
4606 => "000001110110111100100100",
4607 => "000001010001100111100100",
4608 => "000000001111011010010011",
4609 => "111111110010100000011000",
4610 => "000010000000000010000011",
4611 => "000110100111011011000100",
4612 => "001100010110010110101010",
4613 => "010001011010000110011010",
4614 => "010100110110011000010100",
4615 => "010111010001101111110000",
4616 => "011000011100001000111101",
4617 => "010111111010100101011110",
4618 => "010101100111100111110010",
4619 => "010001111010110100010110",
4620 => "001110010111010110011110",
4621 => "001010101011000000010111",
4622 => "000101111101101001111100",
4623 => "000001101011010001111011",
4624 => "111110110011110001110111",
4625 => "111101010111101111110110",
4626 => "111101000001001001010000",
4627 => "111101001001001100000010",
4628 => "111101101110010101110010",
4629 => "111110110111111110101011",
4630 => "000001001010000101110001",
4631 => "000011111001000000110010",
4632 => "000101001011000001011010",
4633 => "000101010110100010010010",
4634 => "000101010000101010111111",
4635 => "000100111000111001011010",
4636 => "000100100000101110011010",
4637 => "000011110111010000000111",
4638 => "000001111101101101110101",
4639 => "111100110010111110111111",
4640 => "110100011100011010100000",
4641 => "101100111010001100101110",
4642 => "101000100111100011111110",
4643 => "100110101000011001011100",
4644 => "100101010011101101011111",
4645 => "100100101101000101100011",
4646 => "100110000111000110000110",
4647 => "101000010111100001010000",
4648 => "101010011011010100001000",
4649 => "101101101101001000111010",
4650 => "110010000100100110000000",
4651 => "110101111100011001111001",
4652 => "111000101101100001100100",
4653 => "111010110010110001100000",
4654 => "111100001101001111010000",
4655 => "111011110011010101010111",
4656 => "111001011010110111100100",
4657 => "110110010101110100000000",
4658 => "110011111101000000101110",
4659 => "110010101110101001011000",
4660 => "110001101100111000111000",
4661 => "110000001001111000010110",
4662 => "101110110010111100010000",
4663 => "101111010011000000001010",
4664 => "110001110101010000100110",
4665 => "110100110001100101100100",
4666 => "111000101001000011000101",
4667 => "111101111101010010100010",
4668 => "000010100000010100110000",
4669 => "000101000011110100010001",
4670 => "000110010100001010111010",
4671 => "000111010110001001010110",
4672 => "000111101110101001101101",
4673 => "000101111000100111111110",
4674 => "000010101100111111010100",
4675 => "000000010101100011101110",
4676 => "111111111010111100010010",
4677 => "000001001110111101100111",
4678 => "000011000001100111100101",
4679 => "000101101001011001011101",
4680 => "001001010001011010000010",
4681 => "001100001100010011011110",
4682 => "001101111001101111110010",
4683 => "001110111010110000001110",
4684 => "001111100001111100010100",
4685 => "001111101011101001000100",
4686 => "001111001010000001000110",
4687 => "001110010001110010111100",
4688 => "001101000010111100011000",
4689 => "001011100111101011000010",
4690 => "001010110011000011001101",
4691 => "001011001110100001000010",
4692 => "001100110110110111110100",
4693 => "001110000101000110000110",
4694 => "001110001000101001101000",
4695 => "001101111111100101001110",
4696 => "001101100101000010010000",
4697 => "001100100100001011100000",
4698 => "001011011011100100000110",
4699 => "001011000101101111101000",
4700 => "001011011110000101111100",
4701 => "001010010001110101010101",
4702 => "000110011001111010100100",
4703 => "000000100111011010111111",
4704 => "111001110000100110110011",
4705 => "110011001011011001100110",
4706 => "101100111110000001111100",
4707 => "100111011111000001100011",
4708 => "100101001001111101010101",
4709 => "100110000110110011000001",
4710 => "101000011100100000100010",
4711 => "101100000110101001010000",
4712 => "110001010101011010011000",
4713 => "110110110010111000000100",
4714 => "111011010111101001010101",
4715 => "111111010111000011001100",
4716 => "000010000011101000010111",
4717 => "000001110101111110010111",
4718 => "111111101100011101001101",
4719 => "111101110111010111111100",
4720 => "111100101010000000110011",
4721 => "111011010010101111010101",
4722 => "111001101000001011100111",
4723 => "111000000001011111111001",
4724 => "110110010100000100000001",
4725 => "110011110001011010011110",
4726 => "110000011010010000111110",
4727 => "101100110110111111101100",
4728 => "101001100101100101001110",
4729 => "100111100111111011010001",
4730 => "100111101011101011010001",
4731 => "101000011101010101111000",
4732 => "101001010011000010011010",
4733 => "101100010111100011100110",
4734 => "110010010010010001010010",
4735 => "110111101111000111100110",
4736 => "111011010101010010011010",
4737 => "111111011011001001000010",
4738 => "000100100100010110011110",
4739 => "001001111110101001111010",
4740 => "001111010000001011111010",
4741 => "010010001111110111101100",
4742 => "010010011111111101010110",
4743 => "010001111011111101100100",
4744 => "010000111111001000011110",
4745 => "001111101101001100000000",
4746 => "001101010000011011000010",
4747 => "001001000000010011101000",
4748 => "000101101000101010000110",
4749 => "000011110010100001110010",
4750 => "000001001100001111010001",
4751 => "111110100101011111110101",
4752 => "111110010111000110110000",
4753 => "000001001001011011100110",
4754 => "000101101100011101001111",
4755 => "001010100101010000100000",
4756 => "010000000110111110001000",
4757 => "010110010100110001000110",
4758 => "011011010110111011101110",
4759 => "011101100101011111000000",
4760 => "011101010101100100100001",
4761 => "011100010111110110111010",
4762 => "011011101001000110101111",
4763 => "011001100110111011111111",
4764 => "010101000000000010011010",
4765 => "001111111100001011110100",
4766 => "001100010111100010101010",
4767 => "001000101001100100100110",
4768 => "000011011101010101011110",
4769 => "111110101010111101010001",
4770 => "111100001101101010100111",
4771 => "111011010101111011001001",
4772 => "111011001011110110101001",
4773 => "111101000001011010100110",
4774 => "000001011100011111110101",
4775 => "000110100010011110001110",
4776 => "001010101010011000010011",
4777 => "001110101101000101100000",
4778 => "010010011100100000001010",
4779 => "010010011111001001111010",
4780 => "001111000001000010111010",
4781 => "001011010110000100101111",
4782 => "000111001101001100100111",
4783 => "000000111100110101110100",
4784 => "110110110001001110101111",
4785 => "101010000111110001111100",
4786 => "100010100011100101011111",
4787 => "100001101010011000111111",
4788 => "100010011011100101101001",
4789 => "100100010000110110100101",
4790 => "100111010100011000111101",
4791 => "101001101010110011000110",
4792 => "101011000011001100010010",
4793 => "101100111010011110110100",
4794 => "110000111010100001011000",
4795 => "110101110110000000100110",
4796 => "111001000100001101101101",
4797 => "111010111000000011000100",
4798 => "111101010101010110001011",
4799 => "000000110101010100000001",
4800 => "000010111011111001111001",
4801 => "000001110000010110100001",
4802 => "111110100000010011101011",
4803 => "111011001100101110100101",
4804 => "111000000011011000111011",
4805 => "110011101011110111110110",
4806 => "101111011101110111011110",
4807 => "101110101011101010000100",
4808 => "110001000001110110000000",
4809 => "110101001101111100101111",
4810 => "111010111111001001011100",
4811 => "000001101001100010011001",
4812 => "001000110001110111101100",
4813 => "001110011010100100110100",
4814 => "010000101011001011101100",
4815 => "010000010001011000110010",
4816 => "001101100111101001110100",
4817 => "001001010000100100111110",
4818 => "000100111001110100011001",
4819 => "000010000010011110110010",
4820 => "000010000010111010010001",
4821 => "000100111110111110100111",
4822 => "001001100000001011110111",
4823 => "001110111110011000110110",
4824 => "010100101100001001010010",
4825 => "011000010101011110110101",
4826 => "011000010001000100101101",
4827 => "010110000100010100110110",
4828 => "010100001011000000011100",
4829 => "010010011011001011010100",
4830 => "001111101000111001100100",
4831 => "001100110000011001001110",
4832 => "001011000010000100001011",
4833 => "001001100000001011111001",
4834 => "001000000010001101000101",
4835 => "000111111111000111101111",
4836 => "001000111111101111011000",
4837 => "001001110000000001000001",
4838 => "001001001110000101100001",
4839 => "000111011101010010010111",
4840 => "000110000001000110111111",
4841 => "000101000100110100000001",
4842 => "000011011110011000100000",
4843 => "000000111011001101110101",
4844 => "111101110101001011101111",
4845 => "111010110001101110000110",
4846 => "110111011101100110011110",
4847 => "110011011001000100000100",
4848 => "101111100100010101010010",
4849 => "101101001101011111111000",
4850 => "101011111010001111111100",
4851 => "101010101000110110000000",
4852 => "101010011101000111100110",
4853 => "101100100001100101000110",
4854 => "101111100000100010110000",
4855 => "110010011001000100010010",
4856 => "110100010010010010001000",
4857 => "110100010110001111011010",
4858 => "110100001101000001001100",
4859 => "110100011100111101000110",
4860 => "110100010100101000110101",
4861 => "110100101000100001000111",
4862 => "110101011100001111100100",
4863 => "110110010101100111100111",
4864 => "110111011101010110110101",
4865 => "110111111000101100011010",
4866 => "110110111010101100010111",
4867 => "110100010011111010011010",
4868 => "110000001010000111110110",
4869 => "101100001100000001000110",
4870 => "101001111010111110011100",
4871 => "101001000001110110010000",
4872 => "101000100000100101010100",
4873 => "101000011001010011101110",
4874 => "101001111011010110100010",
4875 => "101101001001100010110010",
4876 => "110001001100010101110010",
4877 => "110110000110001100100000",
4878 => "111010110111101011010110",
4879 => "111110010001001110010000",
4880 => "000001001000000110110111",
4881 => "000100000101001100111011",
4882 => "000111000011000110101010",
4883 => "001010010100111010000000",
4884 => "001101111011111011110010",
4885 => "010001010000000101000010",
4886 => "010010010001110011000010",
4887 => "010000001101001100101000",
4888 => "001101011010011101101100",
4889 => "001010101111110110100110",
4890 => "000110111110001000001011",
4891 => "000010110011001110000000",
4892 => "000000000011101111100001",
4893 => "111111101001100001001101",
4894 => "000001010000011000001011",
4895 => "000100001000110011110001",
4896 => "001000001101101110111100",
4897 => "001101000101110000111010",
4898 => "010001000101100010100010",
4899 => "010010101010000000100010",
4900 => "010010100100000011110100",
4901 => "010010101100111110111110",
4902 => "010011000110011111000100",
4903 => "010010011001110000111010",
4904 => "010000001001111010001000",
4905 => "001110000101111011100010",
4906 => "001101101111011101011100",
4907 => "001101100010100101100010",
4908 => "001100010010110010000000",
4909 => "001010110001111010101110",
4910 => "001001000110011101100010",
4911 => "000111000010000101000111",
4912 => "000100011010001110011001",
4913 => "000001011111011100011101",
4914 => "111110110101111010001011",
4915 => "111100011101000100011100",
4916 => "111011101110101100011011",
4917 => "111110001011001100101000",
4918 => "000011001000100000101011",
4919 => "001001010100111000000000",
4920 => "001110001100010011010110",
4921 => "001111010101000110110010",
4922 => "001100111100100000101100",
4923 => "000111110010001011001011",
4924 => "000001110100010111011110",
4925 => "111100101110011110010001",
4926 => "110101000010101100110011",
4927 => "101001100101001000011010",
4928 => "100001101110010000100110",
4929 => "100001001011001011101011",
4930 => "100010100111100100011001",
4931 => "100011001000100000010111",
4932 => "100100010111110011011011",
4933 => "100110110101011111001111",
4934 => "101001110000001001010000",
4935 => "101011111101110010110010",
4936 => "101101110010101110000100",
4937 => "110001001011010101000110",
4938 => "110101110011011000100100",
4939 => "111001011111001101111000",
4940 => "111100001110111001110110",
4941 => "000000010101010101100101",
4942 => "000101010011001111100001",
4943 => "000111011110010100001010",
4944 => "000110000010001010100100",
4945 => "000010100100101010011110",
4946 => "111110101000001000011101",
4947 => "111011011001001100101100",
4948 => "110111011101011100101001",
4949 => "110011000011011111101100",
4950 => "110010100111000010111100",
4951 => "110111101100000001000110",
4952 => "111111110110011110011000",
4953 => "001000110111001000100111",
4954 => "010001001011110100111000",
4955 => "010111001100000100100110",
4956 => "011001101100111110010011",
4957 => "011001010000111010110101",
4958 => "010110110110000001111110",
4959 => "010010110111001000011100",
4960 => "001110010001001110011110",
4961 => "001010110000101001011010",
4962 => "001010010100010000000000",
4963 => "001100111100111110010000",
4964 => "010001001110011010111100",
4965 => "010110100110110000010110",
4966 => "011010110010010110010001",
4967 => "011011010101010100110000",
4968 => "011010000100000110011000",
4969 => "011001011001100100000011",
4970 => "011001010111001100011101",
4971 => "011000100011111011000000",
4972 => "010101101110111100110100",
4973 => "010010000101000101000010",
4974 => "001111100100001100101010",
4975 => "001101111010111001111000",
4976 => "001100001110010111010000",
4977 => "001010101100110011010010",
4978 => "001001101000110111111000",
4979 => "001000011011001011110001",
4980 => "000101110100100100011100",
4981 => "000001000101100100001000",
4982 => "111011011011101100101001",
4983 => "110110100111110100000000",
4984 => "110010100111000011101000",
4985 => "101111010011101111111010",
4986 => "101101111111010011111110",
4987 => "101111010100101011101100",
4988 => "110001111101101010000110",
4989 => "110100001001101010010101",
4990 => "110110011011100011100000",
4991 => "111001001100011111101000",
4992 => "111001110100000011101100",
4993 => "110111100101000101000110",
4994 => "110101101000100011100101",
4995 => "110101001001011100000001",
4996 => "110100000000011011101110",
4997 => "110001000000011100100100",
4998 => "101101010111100010110000",
4999 => "101010101101100100010010",
5000 => "101001010100010101101100",
5001 => "101000101101101111111110",
5002 => "101000111110010110010110",
5003 => "101010000111001111011100",
5004 => "101011110000111001010000",
5005 => "101110001100010111000110",
5006 => "110001000100010011000000",
5007 => "110011001100001011010100",
5008 => "110100110111111010101110",
5009 => "110110110100001001110010",
5010 => "111000100101011110100010",
5011 => "111001110011000101010001",
5012 => "111010011101100111000000",
5013 => "111010110010001011101110",
5014 => "111001111111111000011011",
5015 => "110111101000111010001111",
5016 => "110110000110100110100000",
5017 => "110110100100000001100000",
5018 => "110111001101010001000110",
5019 => "110111101010011111111111",
5020 => "111000011110110001000011",
5021 => "111001010110001000000000",
5022 => "111010000011001010001100",
5023 => "111010101111110110101101",
5024 => "111100100101111101100001",
5025 => "111111111011110111110101",
5026 => "000011001011101101001010",
5027 => "000101111011100011010010",
5028 => "001000010100111010110101",
5029 => "001001100011111111010110",
5030 => "001010000001111101101110",
5031 => "001010010011010001000011",
5032 => "001010000101011110001110",
5033 => "001001101110100011111100",
5034 => "001001101011000000001011",
5035 => "001010011110000111110010",
5036 => "001011111101011001010110",
5037 => "001100011011000001110000",
5038 => "001100000011100111100000",
5039 => "001100011001110101100010",
5040 => "001100101001111010100010",
5041 => "001011011110010011111010",
5042 => "001000100110000001000010",
5043 => "000100100010101101010011",
5044 => "000001001110000100100100",
5045 => "000000010101100111001100",
5046 => "000001010110101100011001",
5047 => "000010001100111000110000",
5048 => "000010011110101101011011",
5049 => "000011111000110000101110",
5050 => "000110011001101010011000",
5051 => "001000100111000111000001",
5052 => "001010000011111001111001",
5053 => "001010000010010110111100",
5054 => "001000001110011000110010",
5055 => "000101110110000111111010",
5056 => "000100001100111111110011",
5057 => "000011101110111110110111",
5058 => "000011011100000011110011",
5059 => "000010111100011110010001",
5060 => "000100010100011101001100",
5061 => "000111011001010111010000",
5062 => "001000011011000000100010",
5063 => "000101001000111011010011",
5064 => "111110010010100011011111",
5065 => "110111110111101010101010",
5066 => "110100101001011011100110",
5067 => "101111001000011000101000",
5068 => "100101011111100001010110",
5069 => "100001001000110100011111",
5070 => "100011011010100000101001",
5071 => "100100110001000111010100",
5072 => "100101011011010011100101",
5073 => "100110110000010101011101",
5074 => "100111011010110101110011",
5075 => "101010001000011011000000",
5076 => "101110100000011001010100",
5077 => "110010000111000110111100",
5078 => "111000000010101110110100",
5079 => "000000000110101111110101",
5080 => "000100110110110111100001",
5081 => "000101100111001011011000",
5082 => "000101100111100110001101",
5083 => "000110000100000001101111",
5084 => "000101001000010110010101",
5085 => "000000111110101000111100",
5086 => "111011100100010101000100",
5087 => "110111101111100100001100",
5088 => "110100110100110101010100",
5089 => "110001110111110101011000",
5090 => "110000011001100101011000",
5091 => "110010100000010001011000",
5092 => "111000100110001100001100",
5093 => "000000101100101100100111",
5094 => "001001111000111011000100",
5095 => "010100001111000110110010",
5096 => "011100001000101001010001",
5097 => "011110101011110111101001",
5098 => "011110000110011011100111",
5099 => "011100011010111010000111",
5100 => "011001111111110010100111",
5101 => "010110111001011000100100",
5102 => "010010100010000011001000",
5103 => "001110110100010010000110",
5104 => "001110011111111011000110",
5105 => "010000001010001101110110",
5106 => "010010100011001110011100",
5107 => "010110101100110100100100",
5108 => "011010011011001101010011",
5109 => "011010111111111111111101",
5110 => "011001101100000100111111",
5111 => "010111010010111101101000",
5112 => "010011011001110101011000",
5113 => "001111101011110101101100",
5114 => "001101100111111100001110",
5115 => "001100111001111100010100",
5116 => "001100010111000100011010",
5117 => "001010010001010010101111",
5118 => "000110011101110100011100",
5119 => "000010001110010111110101",
5120 => "111101011111100110000001",
5121 => "110111111101100011011010",
5122 => "110010101110001110100100",
5123 => "101110101001100011111010",
5124 => "101100000010001110011000",
5125 => "101011101100001101110000",
5126 => "101101110110000101001100",
5127 => "110001101110100000110000",
5128 => "110111000101101100110010",
5129 => "111100110110100101000111",
5130 => "111111111111101010101010",
5131 => "111111011101010101101010",
5132 => "111101110001011000101101",
5133 => "111100010110001111101111",
5134 => "111001001010101110101011",
5135 => "110011100010111111101100",
5136 => "101111001000000010101100",
5137 => "101110110000000010000000",
5138 => "110000100011100111101110",
5139 => "110001101101001101111110",
5140 => "110010000111111101111000",
5141 => "110011010111001101011110",
5142 => "110101011010111100101000",
5143 => "110101111110010111010000",
5144 => "110100001001000010101001",
5145 => "110010011100111010110000",
5146 => "110011000110111110011110",
5147 => "110101110011011101101100",
5148 => "111001100001010010100100",
5149 => "111101100001000101101110",
5150 => "000001011110001110001010",
5151 => "000101010010100111111100",
5152 => "001000001100011001111001",
5153 => "001001100110010101000001",
5154 => "001010000111101100001000",
5155 => "001010000010011001110010",
5156 => "001000110010101111011000",
5157 => "000110101100010111010011",
5158 => "000101001110011000111000",
5159 => "000101000111101010100000",
5160 => "000101010100000011111110",
5161 => "000100101000001101101000",
5162 => "000010111011101001010100",
5163 => "000000010010101011011101",
5164 => "111101001100000101100110",
5165 => "111010110111000010001011",
5166 => "111001111110011100000100",
5167 => "111010011010010111011011",
5168 => "111100010101110111011011",
5169 => "000000000100010000010001",
5170 => "000101000000001101001011",
5171 => "001010000010010010010101",
5172 => "001110110111000000010110",
5173 => "010011010011010111010010",
5174 => "010101111101101111001110",
5175 => "010110000101100100100100",
5176 => "010100100101011110110110",
5177 => "010001101101001101001010",
5178 => "001101001111101110110100",
5179 => "001000010101111111000000",
5180 => "000100010110111111010101",
5181 => "000001101011101011010010",
5182 => "111111101001101000100111",
5183 => "111101100101011011100001",
5184 => "111100001011101111110000",
5185 => "111011111100001000110000",
5186 => "111100010001001010100101",
5187 => "111101000011010101011011",
5188 => "111110001110111001110001",
5189 => "111111101010001111111110",
5190 => "000001011001110000111010",
5191 => "000010100100111100101101",
5192 => "000010101010011011101010",
5193 => "000010110111000010110111",
5194 => "000011101010010011001101",
5195 => "000100000110101100000101",
5196 => "000100000101101011011000",
5197 => "000100010011001001010000",
5198 => "000100001100110110010000",
5199 => "000010101010101101111010",
5200 => "000000000100001101010110",
5201 => "111110000110101011100001",
5202 => "111101101000010001011110",
5203 => "111101001000000001100101",
5204 => "111010110101110000000000",
5205 => "110111100101010100101110",
5206 => "110100000010010000000110",
5207 => "101101111110010111110110",
5208 => "100101110010111111001010",
5209 => "100001000011011000111100",
5210 => "100001010000000111001110",
5211 => "100010000110100001111111",
5212 => "100011000000011110001001",
5213 => "100101000110100000110111",
5214 => "100101111101000011111111",
5215 => "100110100011111110010001",
5216 => "101011011111111101101110",
5217 => "110011111000110110111100",
5218 => "111011111010111000101001",
5219 => "000011100111110011110000",
5220 => "001010100100010101001110",
5221 => "001100110001100000100100",
5222 => "001010000101011101001011",
5223 => "000110111101110111001100",
5224 => "000100000011001110101111",
5225 => "111111010100111010000111",
5226 => "111001111110100011100001",
5227 => "110110001101100101001100",
5228 => "110100100011101111101010",
5229 => "110011111111100111111000",
5230 => "110010111111111100011010",
5231 => "110010001111010100101000",
5232 => "110100010000001000111011",
5233 => "111001100010101111011100",
5234 => "000000000000100010001111",
5235 => "000110100000100111101001",
5236 => "001101100010110011011110",
5237 => "010100001110111111110010",
5238 => "011000110010111110011001",
5239 => "011011010001101001001001",
5240 => "011100011001111000111001",
5241 => "011011101011011011010111",
5242 => "011000101100011101100111",
5243 => "010100100100101001011010",
5244 => "010001011100001100110010",
5245 => "010000110101000010100100",
5246 => "010001010100010001011000",
5247 => "010000100101100111010100",
5248 => "001111111001010110000100",
5249 => "010000000101111001100010",
5250 => "001110011101111100100100",
5251 => "001010100111111100010010",
5252 => "000110101110110001011110",
5253 => "000011101001111111011100",
5254 => "000001110000010101100101",
5255 => "000000010101010010101011",
5256 => "111101111111111100111011",
5257 => "111010010101011100000110",
5258 => "110100101110010010100010",
5259 => "101101110101101000010110",
5260 => "101000011111001111010110",
5261 => "100101110101100011101111",
5262 => "100100111101011111001101",
5263 => "100101011010011111010111",
5264 => "100111010010100001000110",
5265 => "101010110111011001001100",
5266 => "110000011100101011110000",
5267 => "110110111010101101110111",
5268 => "111100110101110011100000",
5269 => "000010010010101100011101",
5270 => "000101101100000001000100",
5271 => "000100010111010010011000",
5272 => "111111110110010110110111",
5273 => "111011000010110010111010",
5274 => "110110001000100111111110",
5275 => "110001000111001010000000",
5276 => "101101000111110111100010",
5277 => "101011110010001101110110",
5278 => "101101011110111001011010",
5279 => "101111101011101010010110",
5280 => "101111101011100111111100",
5281 => "101101111011011100111100",
5282 => "101100110111111011110000",
5283 => "101101110100001000010110",
5284 => "110000001100100011011110",
5285 => "110011101001001101111100",
5286 => "111000110111011101100011",
5287 => "000000010101001110000011",
5288 => "001000010111010100110011",
5289 => "001110010011011000111010",
5290 => "010001111100111001111110",
5291 => "010100100110101000010110",
5292 => "010110000011001110000000",
5293 => "010101001001001000101010",
5294 => "010001111111001001100000",
5295 => "001110010110000001001110",
5296 => "001010111111110101100000",
5297 => "000111100010010001000100",
5298 => "000100111010101001100111",
5299 => "000100001101011101100010",
5300 => "000100100100101110100010",
5301 => "000011110111100110100111",
5302 => "000001011001010011110110",
5303 => "111111000100000011100100",
5304 => "111101010011101111101111",
5305 => "111011011000111001110101",
5306 => "111011000101010100111111",
5307 => "111101101000101100001101",
5308 => "000010010010111100111110",
5309 => "001000010110010101001011",
5310 => "001110100010110110101100",
5311 => "010011101000101111011010",
5312 => "010111001100011101111000",
5313 => "011000111111001011110110",
5314 => "011000111101111111110011",
5315 => "010111101011101101110010",
5316 => "010101111000010101011110",
5317 => "010011010100000101001010",
5318 => "001111101011100101000000",
5319 => "001011100010010100111100",
5320 => "000111100000010011101101",
5321 => "000100011010010011010100",
5322 => "000001111010010101010010",
5323 => "111110111101000100001101",
5324 => "111100100110001111100010",
5325 => "111011111000110010001001",
5326 => "111011111111000001011100",
5327 => "111011111001110010000011",
5328 => "111011100101000001100110",
5329 => "111100000111010111000110",
5330 => "111110010111100110010110",
5331 => "000010000011101011100011",
5332 => "000110001010110100010011",
5333 => "001001100001010111011100",
5334 => "001100010010011111111010",
5335 => "001110100011110001000110",
5336 => "001110110001001110100000",
5337 => "001100011011000111001010",
5338 => "001000101111100001101000",
5339 => "000100100011001100010100",
5340 => "000000000100110110101001",
5341 => "111100000110100000101010",
5342 => "111001010110100101010001",
5343 => "110111100010010111101000",
5344 => "110110010010011101110011",
5345 => "110101000010110110111110",
5346 => "110011000111101011111010",
5347 => "101111100001111111101000",
5348 => "101000111010110011110000",
5349 => "100010101010111011000101",
5350 => "100001110001101101000101",
5351 => "100011101100000001111000",
5352 => "100100100011101010001101",
5353 => "100101001001110111000101",
5354 => "100110111100101000110000",
5355 => "101011011111110110101000",
5356 => "110010001010111100111010",
5357 => "111000110001111110010111",
5358 => "111111110101010010110010",
5359 => "000110101011111001001100",
5360 => "001010110110111010010110",
5361 => "001011110010111100101000",
5362 => "001010000011100000101111",
5363 => "000111111000111000011011",
5364 => "000111100001110110101111",
5365 => "000111000101000110001000",
5366 => "000100011000101001110100",
5367 => "000000111001010111010001",
5368 => "111110001110000111001101",
5369 => "111100011000110110110001",
5370 => "111010111100111011101110",
5371 => "111001010111001101010000",
5372 => "111001010001010100111110",
5373 => "111101001110010011001001",
5374 => "000100000001011011101000",
5375 => "001011001111000110011000",
5376 => "010010001101000110000000",
5377 => "011000001101110111010001",
5378 => "011011111110011010101000",
5379 => "011100011011001011110001",
5380 => "011011000110000110010000",
5381 => "011001110110111001000011",
5382 => "010110110011111001111110",
5383 => "010001100001001110101100",
5384 => "001100011110011100000010",
5385 => "001001000111011011111000",
5386 => "001000101010010001111100",
5387 => "001010001100101000111010",
5388 => "001011100011101100001100",
5389 => "001100011000001011101100",
5390 => "001011010111011001110010",
5391 => "001000001000100010010110",
5392 => "000011101110100001100010",
5393 => "111101110101011011100011",
5394 => "110111001111111001111101",
5395 => "101111111011001011010010",
5396 => "100111011100001010100111",
5397 => "100001110110101011011011",
5398 => "100001000110010010001101",
5399 => "100001101000000100111000",
5400 => "100001111010101100010001",
5401 => "100011000000010111111111",
5402 => "100101110000101010100011",
5403 => "101011010100111000111110",
5404 => "110010010101000111101100",
5405 => "110111110010111100001000",
5406 => "111100011110010100100111",
5407 => "000000111011110000110001",
5408 => "000010100010000100011111",
5409 => "000001010111011101101100",
5410 => "111111001100001111000011",
5411 => "111100010011010110111110",
5412 => "111001001101010101100000",
5413 => "110101010001100100110100",
5414 => "110000011110010011100110",
5415 => "101100100110001001111110",
5416 => "101001111010100110001110",
5417 => "101000100000011000011010",
5418 => "101000110001000110000000",
5419 => "101010000111111100011010",
5420 => "101011110101010011000000",
5421 => "101101100011010000001100",
5422 => "110000101100111011001100",
5423 => "110101110010101110100101",
5424 => "111010101110100111001101",
5425 => "111111000111111111100100",
5426 => "000011111100010010100001",
5427 => "001001100000001011011010",
5428 => "001111000001000011100000",
5429 => "010010100111110101110000",
5430 => "010100111011000111000010",
5431 => "010111001101111100000010",
5432 => "011000011001001011101111",
5433 => "010111110001111111011100",
5434 => "010101000001110101111000",
5435 => "001111110101010000001010",
5436 => "001001111101001001110010",
5437 => "000101101010110100011010",
5438 => "000010111110010010011100",
5439 => "111111111110000000100011",
5440 => "111100000110101110111010",
5441 => "111000010111111100110000",
5442 => "110101101101001110100100",
5443 => "110101001101011010101001",
5444 => "110110111010101100000010",
5445 => "111010100101011000001010",
5446 => "000000011111000010000111",
5447 => "000111011011111010111000",
5448 => "001110000110110111101000",
5449 => "010011010111001000001010",
5450 => "010110010100000110001010",
5451 => "011000001110010000001011",
5452 => "011001100111100000101100",
5453 => "011000111001100111100011",
5454 => "010101010111001010001110",
5455 => "010000011000010011100110",
5456 => "001011101111110101100011",
5457 => "000111001111101001010101",
5458 => "000010011001001000000011",
5459 => "111110001000101110100010",
5460 => "111011001110010001110010",
5461 => "111010001001011000011111",
5462 => "111010010000110111100100",
5463 => "111010000111011011110000",
5464 => "111001011000000111000011",
5465 => "111000100001110111000110",
5466 => "111000101111100111011000",
5467 => "111001111000100110111100",
5468 => "111011000010110011100001",
5469 => "111101011100010011110010",
5470 => "000001001101100111110011",
5471 => "000101001011100100101101",
5472 => "001000110101001101001010",
5473 => "001010111101010001011011",
5474 => "001011100111010011111101",
5475 => "001011110001010001111110",
5476 => "001011111110010010011000",
5477 => "001100100100010111100000",
5478 => "001011011101101000111011",
5479 => "000111111011000011100010",
5480 => "000100101111010101011000",
5481 => "000010101100011000001011",
5482 => "000000100010010100101101",
5483 => "111101101110101010111010",
5484 => "111010101100000010011110",
5485 => "110110010110001100011111",
5486 => "101101101101000101110000",
5487 => "100100001110010100011001",
5488 => "100001101110100000100010",
5489 => "100100001111001010100111",
5490 => "100100111001000110010111",
5491 => "100101111010110000101001",
5492 => "101011111101100100101110",
5493 => "110100000101111011010011",
5494 => "111011000001111010101100",
5495 => "000001101010011000110010",
5496 => "001000000100100010000100",
5497 => "001101011110001001111100",
5498 => "010000100110011100100000",
5499 => "010000110001101001100100",
5500 => "001111101100101101111000",
5501 => "001101101010000010011010",
5502 => "001011000111100110010010",
5503 => "001010000100110110111100",
5504 => "001001100101010000110000",
5505 => "001000111100110110010001",
5506 => "001000111001000100110100",
5507 => "001000100010111011000101",
5508 => "000111001100011111001110",
5509 => "000100111001001011001001",
5510 => "000011101110110110011010",
5511 => "000101001001011010110101",
5512 => "000111000000000101011100",
5513 => "001001100111110110010101",
5514 => "001110010011000000011100",
5515 => "010011000110001011110010",
5516 => "010110111000110000111010",
5517 => "011000111010011000111111",
5518 => "011000110011110100101001",
5519 => "011000001101101011001101",
5520 => "010111010001011001010000",
5521 => "010100111000110111001100",
5522 => "010001101011100110010110",
5523 => "001110111101000100001110",
5524 => "001100100111100101011110",
5525 => "001010001011111010010111",
5526 => "000111110101001111000000",
5527 => "000100101100010010111101",
5528 => "111111101001101010100000",
5529 => "111000101101000110011001",
5530 => "110000110110001011101010",
5531 => "101001111100011001110010",
5532 => "100100011110110111111000",
5533 => "100001000000101110110101",
5534 => "100000101101011010011100",
5535 => "100001010000000010111001",
5536 => "100000101100110110100110",
5537 => "100001100011101000110101",
5538 => "100101110100110001000001",
5539 => "101011001010011100100100",
5540 => "101110000101101111011010",
5541 => "101111110010111110110110",
5542 => "110001111010010001101100",
5543 => "110010000011010011111100",
5544 => "110000110000110011011000",
5545 => "110000111110011101010010",
5546 => "110010111101101010011100",
5547 => "110110000000100011000000",
5548 => "111001000111100111000111",
5549 => "111011101111111011111110",
5550 => "111100100000101110101110",
5551 => "111001010001001101011100",
5552 => "110011001100101000100010",
5553 => "101100010000100110010100",
5554 => "100110001100100110000001",
5555 => "100011110010001000011001",
5556 => "100100011000001111111011",
5557 => "100101001011011101111001",
5558 => "100110100111010000011011",
5559 => "101011110010011100110110",
5560 => "110100111000001010001110",
5561 => "111101010010011011000101",
5562 => "000011001111111000110000",
5563 => "001001010011001100000110",
5564 => "001111011000110101011100",
5565 => "010011010011011001111000",
5566 => "010100101101010001100110",
5567 => "010100110100000110001110",
5568 => "010011111110100000101000",
5569 => "010010011111100011111100",
5570 => "010001100100010011101110",
5571 => "010000001101111011100000",
5572 => "001100111100101111111000",
5573 => "001000010010001111100010",
5574 => "000011001111101001001101",
5575 => "111111111011100101101000",
5576 => "111110111001011010011110",
5577 => "111110100001100100101110",
5578 => "111110110110101001011001",
5579 => "111111100001110110010000",
5580 => "111111101101011001001010",
5581 => "000000000010010111101111",
5582 => "000001000010111010100101",
5583 => "000010111011101010010011",
5584 => "000101000001001000111000",
5585 => "000110101011010001110001",
5586 => "001000000101110101001100",
5587 => "001001010010111001001100",
5588 => "001011000010100010001001",
5589 => "001100001110000101001110",
5590 => "001010111001011101000111",
5591 => "001000111111011001010011",
5592 => "001000000101110101010000",
5593 => "000110110010111001100110",
5594 => "000011100010101011001100",
5595 => "111110110011100011000111",
5596 => "111011011100101011101100",
5597 => "111010001100001101011001",
5598 => "111001010100000000000000",
5599 => "111000010011010001010101",
5600 => "110111010001100000010010",
5601 => "110110101110110110101110",
5602 => "110110100101111001001111",
5603 => "110110100100001000011001",
5604 => "110111011010100111110000",
5605 => "111000101001001010011010",
5606 => "111001101001110010000111",
5607 => "111010101001101010111110",
5608 => "111011100111111100011000",
5609 => "111101011111010111011010",
5610 => "000000001110100011110110",
5611 => "000011000000111111101000",
5612 => "000101101001011011010101",
5613 => "000111010110110000010110",
5614 => "001000001011011000101011",
5615 => "001000010111010111000100",
5616 => "000111111100001110000101",
5617 => "000111100010100010101111",
5618 => "000110100111000110000111",
5619 => "000101000111101011011000",
5620 => "000011100111111011111001",
5621 => "000001010101010100100001",
5622 => "111110010001000101100110",
5623 => "111010001100111111100010",
5624 => "110011110110100110011100",
5625 => "101100010111000111000010",
5626 => "100111110010010111011001",
5627 => "101000001101011011011010",
5628 => "101011001100100010010010",
5629 => "101111011101010110000010",
5630 => "110101010001110101100001",
5631 => "111010101111011100000110",
5632 => "111111010001000010110011",
5633 => "000011001000100011110101",
5634 => "000111000111111000111100",
5635 => "001101010000100111011000",
5636 => "010010100100011100100110",
5637 => "010011101011101010010010",
5638 => "010011000111010100111110",
5639 => "010010110110100001001010",
5640 => "010011000001100011000110",
5641 => "010011011000110001111100",
5642 => "010011010010010101100100",
5643 => "010011010000101100101110",
5644 => "010011010100111000100010",
5645 => "010011001001111010111000",
5646 => "010010100001011101111110",
5647 => "010000101000011101011010",
5648 => "001110111010010111110110",
5649 => "001111101100010101000010",
5650 => "010010001011111100001110",
5651 => "010100010001000010111100",
5652 => "010110001100011101111000",
5653 => "011000010101101011110111",
5654 => "011000110011111000101011",
5655 => "011000001010110111010011",
5656 => "010111111000101100001010",
5657 => "010110001010101010110010",
5658 => "010010110001000010011100",
5659 => "001111100001101101100010",
5660 => "001101101111001101101110",
5661 => "001101001011110000101100",
5662 => "001011011001110101000101",
5663 => "001000100100111111001101",
5664 => "000101110001101110011110",
5665 => "000000100100010001110100",
5666 => "111000100110100101001000",
5667 => "110000001000000001011000",
5668 => "101001001010000001001100",
5669 => "100101010011111001010011",
5670 => "100011111010110001101101",
5671 => "100100000010110010111011",
5672 => "100101100001110101100001",
5673 => "101000001111001101011000",
5674 => "101100100000000000010010",
5675 => "110001001101110011111000",
5676 => "110101001110101100111100",
5677 => "111000001110110000110100",
5678 => "111000110110101011100000",
5679 => "110110110110111111100100",
5680 => "110100001110100001010011",
5681 => "110010101100101100110100",
5682 => "110001110100000111000000",
5683 => "110001101110110010110000",
5684 => "110100100010011010000100",
5685 => "111000001000010010111100",
5686 => "111001000000101011110110",
5687 => "111000110100101100101100",
5688 => "111001000000110010001100",
5689 => "110111110011101100011100",
5690 => "110011111000000110011000",
5691 => "101111100001110010111100",
5692 => "101110010000111001011000",
5693 => "101110111011000000101000",
5694 => "110000001011011101101110",
5695 => "110011001111010111110010",
5696 => "110110100011011001010010",
5697 => "111001000111111111010011",
5698 => "111101001101100011000000",
5699 => "000011110001101100110000",
5700 => "001010001100101101011001",
5701 => "001101101101000101000010",
5702 => "010000001100110111001000",
5703 => "010011011011101101001100",
5704 => "010100110110100110000010",
5705 => "010011011000100101101100",
5706 => "010000110010100111001110",
5707 => "001110101110001011100100",
5708 => "001100101000010100101010",
5709 => "001000100100010100001100",
5710 => "000010110111110110110011",
5711 => "111101100001111101001111",
5712 => "111011000101000010111100",
5713 => "111100101001100001111110",
5714 => "111111101001011011110101",
5715 => "000010010111110100111000",
5716 => "000100111110100100010011",
5717 => "000110110000101101011110",
5718 => "000111000110100011100110",
5719 => "000101110101010111011011",
5720 => "000100010010100011101010",
5721 => "000011100000000100010010",
5722 => "000010010110010011110101",
5723 => "000000011011001110001000",
5724 => "111110000000001000110100",
5725 => "111100001110110100100010",
5726 => "111100001010111001111111",
5727 => "111100011010000110001110",
5728 => "111100010110010010101101",
5729 => "111100010100011010010111",
5730 => "111100001100100111001101",
5731 => "111100000001101010010001",
5732 => "111010100100001011010101",
5733 => "111000000100101011111001",
5734 => "110110010010100001001110",
5735 => "110100110110110001011111",
5736 => "110011001110001000100110",
5737 => "110001010101011111110010",
5738 => "101111111101001110100100",
5739 => "110000001101101000001100",
5740 => "110001010110001101110100",
5741 => "110010101100000111010010",
5742 => "110100010000101100000111",
5743 => "110110011100011000010100",
5744 => "111001010111110011110100",
5745 => "111011000100101111100010",
5746 => "111011100111000101011010",
5747 => "111101101011000110010101",
5748 => "000001010100001100101010",
5749 => "000011111111110101111100",
5750 => "000011111001001100110001",
5751 => "000010100101010110001100",
5752 => "000001111111110011011110",
5753 => "000001011101101010000101",
5754 => "000000111000000011000100",
5755 => "111111110100001011011110",
5756 => "111110001010000110100010",
5757 => "111101110110100001010011",
5758 => "111110101111101101111001",
5759 => "111111011110100100000001",
5760 => "111111001110110010110001",
5761 => "111100110000110101101000",
5762 => "111000100110000001010110",
5763 => "110100010000100111101000",
5764 => "110001000000000110011110",
5765 => "101111111010111010001000",
5766 => "110001000010010100001100",
5767 => "110011011101101110101110",
5768 => "110101110100111011110010",
5769 => "110111111010110110011010",
5770 => "111010010000001101000010",
5771 => "111101011000001101111010",
5772 => "000011001111000001011001",
5773 => "001010110010100011110000",
5774 => "010000100001100101111000",
5775 => "010011111110010001011010",
5776 => "010101100111100000010010",
5777 => "010110001101110111010010",
5778 => "010110010100110011110100",
5779 => "010101001110110001111100",
5780 => "010011111010111111110000",
5781 => "010010111101001011101010",
5782 => "010001110000101111100100",
5783 => "010000001111001001011110",
5784 => "001101011111010010011010",
5785 => "001011000000001010010110",
5786 => "001011000101111110111110",
5787 => "001101000000001100000100",
5788 => "010000000101000001110100",
5789 => "010011011011001111111010",
5790 => "010101010000010000111110",
5791 => "010101100000000111011110",
5792 => "010101001000000011001110",
5793 => "010011111010110011000110",
5794 => "010000100000110100110100",
5795 => "001011100000100000111000",
5796 => "000110110001100011000011",
5797 => "000010101111011111100011",
5798 => "111111101011101000011010",
5799 => "111100100011011000101101",
5800 => "111000101001010010001000",
5801 => "110110000110111011111010",
5802 => "110101000011001000011110",
5803 => "110011001100110101001100",
5804 => "101111111101000100000000",
5805 => "101101000000111110011100",
5806 => "101100100000000010110100",
5807 => "101101111100011100001110",
5808 => "101111110111001101000100",
5809 => "110001100001101110110010",
5810 => "110011001100111011001000",
5811 => "110110000111010000010111",
5812 => "111000010101100000011110",
5813 => "110111101100001011011010",
5814 => "110110100011000110010110",
5815 => "110110110001001011011001",
5816 => "110111001010100011100111",
5817 => "110101011110010111011011",
5818 => "110010011110001010001100",
5819 => "110010010011001001001100",
5820 => "110100010010001111101100",
5821 => "110101000000110000000011",
5822 => "110101001110010010010111",
5823 => "110110010011000010001010",
5824 => "110111111001010011001110",
5825 => "111001011110010111010100",
5826 => "111011101011110010101011",
5827 => "111110010111110001000001",
5828 => "111111000110111111001001",
5829 => "111111011111101011111110",
5830 => "000011001011001010010011",
5831 => "000111110010010101011001",
5832 => "001001011000001100110011",
5833 => "001000100100000010000011",
5834 => "001000100010101101101001",
5835 => "001010001011001110110100",
5836 => "001011110101001010000011",
5837 => "001101010000110111011010",
5838 => "001110101101110110100110",
5839 => "001111111101100010111010",
5840 => "010001001001111100100100",
5841 => "010001111111001111110010",
5842 => "010001101111111101001110",
5843 => "001111101100000000010000",
5844 => "001101011010010110100000",
5845 => "001100110101111001000010",
5846 => "001011011011011011110110",
5847 => "001000010001011100100110",
5848 => "000110000001011111111110",
5849 => "000100110000110111101101",
5850 => "000100001000111110001100",
5851 => "000101010100111110000011",
5852 => "001000010000001001110100",
5853 => "001010100111000011100000",
5854 => "001010101101001110100000",
5855 => "001001101110111101011110",
5856 => "000111101111111000001110",
5857 => "000100010000110010000010",
5858 => "000000111100010101100100",
5859 => "111101111111111000001000",
5860 => "111011010111000000101011",
5861 => "111001010000101011101101",
5862 => "110110110010101010101010",
5863 => "110100111010000101001010",
5864 => "110100000101100001001000",
5865 => "110011010110100000011110",
5866 => "110011011111011111010000",
5867 => "110100110100111110011001",
5868 => "110110010011100001110111",
5869 => "110110111111110111001110",
5870 => "110110011101001011000000",
5871 => "110100110110100100011000",
5872 => "110011000101111011001010",
5873 => "110010100011100001101000",
5874 => "110010011110010000100000",
5875 => "110010000001100001111110",
5876 => "110010101101101000100010",
5877 => "110011100001101101111010",
5878 => "110011001110100010001000",
5879 => "110011110001100011101100",
5880 => "110101100100011110111001",
5881 => "110111001101111101100101",
5882 => "111000000010001011100100",
5883 => "111000101111101111110001",
5884 => "111010010101001001011010",
5885 => "111100010001101010110011",
5886 => "111110010011110101001111",
5887 => "111111011001011010001110",
5888 => "111110101100100100000001",
5889 => "111110101010100011001101",
5890 => "111111101101111101100100",
5891 => "111111110001110001010111",
5892 => "111111100000110001000101",
5893 => "000000000100100110010111",
5894 => "000001000100110000111111",
5895 => "000010001111000000000111",
5896 => "000011101101000110100011",
5897 => "000100110101011011111010",
5898 => "000100001000011101011101",
5899 => "000000011111100000111011",
5900 => "111001111100010101011000",
5901 => "110011110010000101100100",
5902 => "110000101111010111111110",
5903 => "101111000101011111011100",
5904 => "101111001011001011011000",
5905 => "110001101110111100010100",
5906 => "110011111001111101100100",
5907 => "110101110010011011110010",
5908 => "111001001101001010110111",
5909 => "111110111011110010001000",
5910 => "000111010101000110011110",
5911 => "001111001011000010100000",
5912 => "010011101011011000001010",
5913 => "010101111100111010100100",
5914 => "010111010111110000100000",
5915 => "011000011111100000000110",
5916 => "011000101010011100011111",
5917 => "010111011010000101000000",
5918 => "010101100110010100011100",
5919 => "010011111110000100101010",
5920 => "010010110101111101000100",
5921 => "010000111111110010001110",
5922 => "001101100101010011111110",
5923 => "001011001001011101001111",
5924 => "001011100110010100100100",
5925 => "001100110111011100011110",
5926 => "001100111000101111010000",
5927 => "001101000110001000011100",
5928 => "001101110010000000111000",
5929 => "001100010100100001011010",
5930 => "001001000001110000100010",
5931 => "000101001011101101101010",
5932 => "000000001100110101111001",
5933 => "111010111111100100010110",
5934 => "110110100110111110011111",
5935 => "110011000110010110010110",
5936 => "110000000111100001011010",
5937 => "101101101001010011111100",
5938 => "101101101011100000001110",
5939 => "110000001101011000000110",
5940 => "110010100100000111101110",
5941 => "110011101101011111000110",
5942 => "110011101000011001110110",
5943 => "110011010101000100001110",
5944 => "110100010101101101111101",
5945 => "110110100000100010100000",
5946 => "110111100100010100100100",
5947 => "110100111111101100011000",
5948 => "110001000011111000001000",
5949 => "101111001110010101011010",
5950 => "101101111011000101101000",
5951 => "101100101011001110000000",
5952 => "101101101111110111001000",
5953 => "110000101001100011010100",
5954 => "110010110001101111101010",
5955 => "110011001001010111101100",
5956 => "110011101110000110001100",
5957 => "110101001011011110001101",
5958 => "110101011001000111011000",
5959 => "110100010100111000001110",
5960 => "110100001111000000001010",
5961 => "110110101001100000000010",
5962 => "111010100000101001100100",
5963 => "111101101100001100001000",
5964 => "000000101100011101111110",
5965 => "000011110110010101000111",
5966 => "000101101101110111011111",
5967 => "000111001000100011100111",
5968 => "001010011001000010101110",
5969 => "001111001010010111101110",
5970 => "010010001110001001101010",
5971 => "010010010000010001011010",
5972 => "010001110101111001111000",
5973 => "010010111101111110100110",
5974 => "010100110001111011010000",
5975 => "010101010011000110110010",
5976 => "010100101110101100101100",
5977 => "010100011110000001001110",
5978 => "010010111010000000000110",
5979 => "001111011110110111000110",
5980 => "001100010110110011001010",
5981 => "001010011100110000010011",
5982 => "001010110000011000010100",
5983 => "001100110100110011000110",
5984 => "001110011011110110110110",
5985 => "001111100110010010111010",
5986 => "010000111011110000010000",
5987 => "010010100110110010011010",
5988 => "010100000010011101011110",
5989 => "010100001110101001001000",
5990 => "010100011011000011011110",
5991 => "010100010011000110000010",
5992 => "010001001011110100100110",
5993 => "001011100110110001011110",
5994 => "000110010011110001110001",
5995 => "000010110111100111110101",
5996 => "000000101001101111010110",
5997 => "111110000110100000101110",
5998 => "111011000011110101110011",
5999 => "111000010100111111100011",
6000 => "110110110101101101100111",
6001 => "110110100111110101111100",
6002 => "110110110011101101101110",
6003 => "110111001100110011011011",
6004 => "110111110100010100011010",
6005 => "111000010100101011000000",
6006 => "110111110000101101001010",
6007 => "110110001101101000100001",
6008 => "110101101001011111001111",
6009 => "110101111101101010101100",
6010 => "110110001001100011111110",
6011 => "110110111010100100101010",
6012 => "110111111110111110101010",
6013 => "111000011111010000010100",
6014 => "110111111110111010101111",
6015 => "110110110101101000000000",
6016 => "110110100111101110101110",
6017 => "110111101010011100110001",
6018 => "111001000001110011001001",
6019 => "111001000111101001000110",
6020 => "110111101111111010110111",
6021 => "110111111110111000000010",
6022 => "111010011100101110101110",
6023 => "111100110111010011111001",
6024 => "111101111110100110111100",
6025 => "111100111110010101101101",
6026 => "111100000011111110000101",
6027 => "111101101101101000000000",
6028 => "111111100011010000001000",
6029 => "000000100000110111010111",
6030 => "000010000111111011010101",
6031 => "000011011000000011010110",
6032 => "000011010100101000110001",
6033 => "000011011010100010010010",
6034 => "000100000111001100011110",
6035 => "000011000100111101101010",
6036 => "111101100110010110101000",
6037 => "110100101000000100010000",
6038 => "101101101001010010110010",
6039 => "101011111100010101010000",
6040 => "101100111011101001101010",
6041 => "101111011000010110111010",
6042 => "110011110100101100000010",
6043 => "111000000010010010001010",
6044 => "111011001011000001001111",
6045 => "111110001110100111100011",
6046 => "000010010101111101111111",
6047 => "001000110010100011000110",
6048 => "001110110110011001101110",
6049 => "010001001010001001111110",
6050 => "010000101010100010000010",
6051 => "010000000010110100110110",
6052 => "010001100000110001001010",
6053 => "010011000001000001101000",
6054 => "010001100010100111001100",
6055 => "010000010001010001001110",
6056 => "010001101000100010111010",
6057 => "010011010001010000010010",
6058 => "010011100000010110101100",
6059 => "010010001000110101101010",
6060 => "010000101101100100110100",
6061 => "010000110011100101111100",
6062 => "010000101001000101111000",
6063 => "001110110110100000101000",
6064 => "001100110101101110011100",
6065 => "001010010010010100011101",
6066 => "000101000111001010100010",
6067 => "111110101100101001011010",
6068 => "111001011110101100011011",
6069 => "110011010000111011001010",
6070 => "101010011011100111001000",
6071 => "100011011011101011100101",
6072 => "100001100010110001001110",
6073 => "100001100001010110100010",
6074 => "100010000110101010000000",
6075 => "100111010101011011011101",
6076 => "110000101100110101001100",
6077 => "111000111110000100000100",
6078 => "111101000111101101111111",
6079 => "111100110100101001011100",
6080 => "111100000011101011101000",
6081 => "111101110101001011011001",
6082 => "111101100100111100110001",
6083 => "111000100011011000100111",
6084 => "110010011101010011000100",
6085 => "101110010100101110100100",
6086 => "101011010111001010000100",
6087 => "100111111011111011000100",
6088 => "100110110000001001100011",
6089 => "101001011101111110011010",
6090 => "101011000011011001011010",
6091 => "101001100101000111000100",
6092 => "101000010001000010101110",
6093 => "101000001011110000001010",
6094 => "101000100110001011010000",
6095 => "101000101011111100100100",
6096 => "101001110111010000110000",
6097 => "101110101000010100010100",
6098 => "110101011010011110110001",
6099 => "111100001110011100111110",
6100 => "000011001101011111010100",
6101 => "001000100000011001001110",
6102 => "001011000111001100110111",
6103 => "001101010000101100110000",
6104 => "001111010111010110111100",
6105 => "010000101011010111101110",
6106 => "010010000110001001100010",
6107 => "010010100110010101110100",
6108 => "010000100010100101010000",
6109 => "001101110011110101010110",
6110 => "001100111001100011001010",
6111 => "001101101001011001101000",
6112 => "001100110011110100100110",
6113 => "001000100011110111000001",
6114 => "000101000101011111010000",
6115 => "000101001001101111011110",
6116 => "000110000100010100010011",
6117 => "000110100011111011101101",
6118 => "000111111010110010011111",
6119 => "001011000110111011110010",
6120 => "001111011111011000011110",
6121 => "010011100011111111001100",
6122 => "010110101111111110011100",
6123 => "011000000001000000110101",
6124 => "010111011101000100110010",
6125 => "010110110111011110111010",
6126 => "010101111111000101000010",
6127 => "010100010010101000000010",
6128 => "010001011001110111000100",
6129 => "001100100010100001000100",
6130 => "000111110000100110000111",
6131 => "000100010000011001001010",
6132 => "000000101101101111101000",
6133 => "111101100011000001111100",
6134 => "111011000010110110000111",
6135 => "111000111010100110010010",
6136 => "110111111101100001010110",
6137 => "110111101111100011101100",
6138 => "110111000000100000000001",
6139 => "110101110101010011110010",
6140 => "110101010010100110111110",
6141 => "110110010110001000100111",
6142 => "111000010110110011101011",
6143 => "111001011001001010001010",
6144 => "111001000110011111001110",
6145 => "111001011001000110100110",
6146 => "111011100001111110101010",
6147 => "111110011100110101111100",
6148 => "000000011101000101010011",
6149 => "000001100100111101000010",
6150 => "000010110101011011000001",
6151 => "000011101001101100001110",
6152 => "000011010110110010110010",
6153 => "000010100001101111101011",
6154 => "000001010101101011000001",
6155 => "000000010011100110111011",
6156 => "111111001110100100100110",
6157 => "111101000111001001010101",
6158 => "111011110110101100010100",
6159 => "111100011101000111010011",
6160 => "111100110110101101011000",
6161 => "111101101001100000100101",
6162 => "000001001000101101111011",
6163 => "000110111000111001101100",
6164 => "001011100011110111011110",
6165 => "001100100101110011111100",
6166 => "001011101101000110011000",
6167 => "001010111011001011000000",
6168 => "001010000010111010110111",
6169 => "001000111100000101001100",
6170 => "000111100011011110100000",
6171 => "000110010001100101100000",
6172 => "000010110100011011010100",
6173 => "111001111101101011110110",
6174 => "110001101010101010011100",
6175 => "110000111111001100000000",
6176 => "110011101000001000101000",
6177 => "110100101001010000000100",
6178 => "110110000110001100111011",
6179 => "111010000111110010010100",
6180 => "111111100010101000101001",
6181 => "000010111010011011110000",
6182 => "000011010010101000010011",
6183 => "000100110001010111010110",
6184 => "001000110011000101101000",
6185 => "001011101000010010100101",
6186 => "001011110011110111011000",
6187 => "001011010111111000110011",
6188 => "001100001111010000111000",
6189 => "001110011110111011011010",
6190 => "001111101010110100110100",
6191 => "001111001101000111101110",
6192 => "001111111001000110100110",
6193 => "010001111100010001111000",
6194 => "010010110010110000111110",
6195 => "010001010011010100110000",
6196 => "001110010111110111011000",
6197 => "001011101001010101110100",
6198 => "001001011000110100001101",
6199 => "000111100111101111010000",
6200 => "000110110011110011010110",
6201 => "000101001011011000101110",
6202 => "000000111010100111110001",
6203 => "111011011100100010001010",
6204 => "110111010100010010110111",
6205 => "110011011111010111001000",
6206 => "101100001100011011001000",
6207 => "100100000010110000000111",
6208 => "100001000110100111110101",
6209 => "100001101111111000011010",
6210 => "100011001101100111011001",
6211 => "100111011111010111110000",
6212 => "101110001010001001101010",
6213 => "110100001110100100100001",
6214 => "111000000010010101001011",
6215 => "111010000010011110001000",
6216 => "111011110111001001010110",
6217 => "111100111100110011111110",
6218 => "111100010111010110110110",
6219 => "111011001000011101110010",
6220 => "111001000101010010010100",
6221 => "110101111001011100111001",
6222 => "110010111110101000101000",
6223 => "110001000000001100000110",
6224 => "101111110000001111000110",
6225 => "101110100000101110010000",
6226 => "101100110011101100011010",
6227 => "101011011110000011000000",
6228 => "101001100100110100111000",
6229 => "100110100101110010011100",
6230 => "100101111001001011001110",
6231 => "100111010011010010100111",
6232 => "101000000100001100110010",
6233 => "101011100100100010011010",
6234 => "110011101111000010000000",
6235 => "111100000110010010001010",
6236 => "000010000111001111000011",
6237 => "000110100110001011000110",
6238 => "001011010001000011011111",
6239 => "001111111011111001110010",
6240 => "010001010101111110010010",
6241 => "010000000010110110110100",
6242 => "010000001100001100110000",
6243 => "010001111001011000000000",
6244 => "010010000100001001111010",
6245 => "001111011001110110100100",
6246 => "001100110000101000011110",
6247 => "001100100010001000100100",
6248 => "001011110000101100011010",
6249 => "001000110000010101001111",
6250 => "000101111011010101111000",
6251 => "000011111001101101000001",
6252 => "000010111000110101011000",
6253 => "000011100110011010011100",
6254 => "000100101000100100001110",
6255 => "000101111010100100001101",
6256 => "001000110101110101110110",
6257 => "001100011001011100001000",
6258 => "001110110000100000001100",
6259 => "001110111101100110110010",
6260 => "001101011101011101000110",
6261 => "001100100101011100100100",
6262 => "001100111100110000101110",
6263 => "001101000010101011011010",
6264 => "001100011111001110100100",
6265 => "001010100100001010110010",
6266 => "000110011011010000110110",
6267 => "000001101100111000011010",
6268 => "111101101101011010101000",
6269 => "111010000000100111111000",
6270 => "110110101010110011000011",
6271 => "110011111011110100110110",
6272 => "110001101101001110000110",
6273 => "110000000100010101000110",
6274 => "101110110111101010110010",
6275 => "101110000010010101101100",
6276 => "101110010111011001010100",
6277 => "110000101001100101101110",
6278 => "110011110110001110101000",
6279 => "110110000010110000110110",
6280 => "110111100001010100110100",
6281 => "111001111010001111100010",
6282 => "111100111110010101010110",
6283 => "111111010100100010010100",
6284 => "000000111011101010110110",
6285 => "000010101101000110001001",
6286 => "000100011110000101101110",
6287 => "000100111101011000011111",
6288 => "000011100100111011110100",
6289 => "000001111110100011110011",
6290 => "000010100110010101111100",
6291 => "000100110001100110001100",
6292 => "000101111010101001001101",
6293 => "000110000001000001100101",
6294 => "000110000100001010000011",
6295 => "000101111001110011101110",
6296 => "000110001111001110101101",
6297 => "000111111100000100111001",
6298 => "001010100010110111111110",
6299 => "001100111001100101100110",
6300 => "001101101011101000000000",
6301 => "001101010011011101010100",
6302 => "001101101010010100001000",
6303 => "001110101010001111110110",
6304 => "001110110100110011100100",
6305 => "001110000111101110010010",
6306 => "001101100111011000011100",
6307 => "001101001011101101001100",
6308 => "001010010000110111101010",
6309 => "000011011111011001000101",
6310 => "111100011110110011000110",
6311 => "111001010101100011001011",
6312 => "111001011011011011001011",
6313 => "111010011001000101001011",
6314 => "111011111011011101000111",
6315 => "111110100010101010010100",
6316 => "000001101111000100100111",
6317 => "000100011101101010111011",
6318 => "000110001111001110010100",
6319 => "000111111110010001100100",
6320 => "001011000000110001000010",
6321 => "001110001101010110000100",
6322 => "001111000010010110001010",
6323 => "001110001101001011111010",
6324 => "001110010101101110011100",
6325 => "001111110000010110101010",
6326 => "010000101010100111110100",
6327 => "001110110100010010100000",
6328 => "001010101011101011010100",
6329 => "001000010001110001111010",
6330 => "001000101001101110101110",
6331 => "001000101000111101010100",
6332 => "000110110010011000100101",
6333 => "000100010011001100001010",
6334 => "000011001110000000101110",
6335 => "000100001000000011001110",
6336 => "000101000001001011011100",
6337 => "000100110101011100001101",
6338 => "000010111001010111100010",
6339 => "111101110110100010010100",
6340 => "110111101010111101111101",
6341 => "110001100100010000000000",
6342 => "101001100101000000010000",
6343 => "100010101001001101000110",
6344 => "100000111000010101001001",
6345 => "100001011001000111011101",
6346 => "100000111100001110101001",
6347 => "100000111011101011110101",
6348 => "100100000110011101100111",
6349 => "101011101010101100101110",
6350 => "110100110100110111010000",
6351 => "111011011001111010111110",
6352 => "111110010100101100000100",
6353 => "111110000111111001010011",
6354 => "111100010110010010111110",
6355 => "111011000001111100101011",
6356 => "111001100110100011011101",
6357 => "110110011000110101111000",
6358 => "110001100111111110010000",
6359 => "101101001101000010110000",
6360 => "101010110110011000100110",
6361 => "101001111001000110000100",
6362 => "101000110110010101110110",
6363 => "100111111011111101010111",
6364 => "100111100000100110000111",
6365 => "100111110000110110000101",
6366 => "101001001011001010100010",
6367 => "101011100010101111001110",
6368 => "101111000100100111101100",
6369 => "110011111011110010111000",
6370 => "111001000110000101010001",
6371 => "111110000011101001000101",
6372 => "000010011011101101100110",
6373 => "000101011110110001010000",
6374 => "000111110100011010000011",
6375 => "001001101100101001010110",
6376 => "001010011011110001101100",
6377 => "001011010110111001001100",
6378 => "001110010001111010010000",
6379 => "010001111100100110110100",
6380 => "010011100001111111101000",
6381 => "010010100011110101011000",
6382 => "010001001110000010110000",
6383 => "010001000010000000100100",
6384 => "010001011110001101001110",
6385 => "010000011000110000110000",
6386 => "001011011110100110100010",
6387 => "000100111100000011100110",
6388 => "000001110101011111011000",
6389 => "000001111101011101100011",
6390 => "000001111100001101111011",
6391 => "000010000000110010010101",
6392 => "000011101010000001001000",
6393 => "000110100100100010111010",
6394 => "001001001010001000110010",
6395 => "001001110101011111010011",
6396 => "001001111100000100101011",
6397 => "001011001111010000101010",
6398 => "001011101011110010111001",
6399 => "001010000010110001111100",
6400 => "000111111001001011100110",
6401 => "000100011011010101111110",
6402 => "111110100011011000111001",
6403 => "111000110010101011111011",
6404 => "110101000110110110000011",
6405 => "110011001000111100010100",
6406 => "110010010000011100100110",
6407 => "110000111110110011110000",
6408 => "101111000111000000010100",
6409 => "101111000001010010110110",
6410 => "110000011000000001110110",
6411 => "110000100111110000010100",
6412 => "110000101000000100001010",
6413 => "110001100111001111110010",
6414 => "110010010110010011000010",
6415 => "110010111011000111101000",
6416 => "110011110110011110110100",
6417 => "110100011000111011001110",
6418 => "110100111000101000101101",
6419 => "110101101001011111111000",
6420 => "110110100101110110111110",
6421 => "111000111000110010100011",
6422 => "111100001110111010010111",
6423 => "111110111010010000111100",
6424 => "000001000000000110101001",
6425 => "000010110100010111011100",
6426 => "000100011110001001000010",
6427 => "000110110001001100011000",
6428 => "001000110010100100010100",
6429 => "001000111110011100100011",
6430 => "000111110111110001001111",
6431 => "000110100110100010000001",
6432 => "000110000101001010111111",
6433 => "000110111110011101110100",
6434 => "001000101100010111110110",
6435 => "001010011000110000001001",
6436 => "001100000010001111011000",
6437 => "001110011110010100101000",
6438 => "010010001111111000100000",
6439 => "010101010101110010000110",
6440 => "010101101100011111111000",
6441 => "010100110011001101010000",
6442 => "010100001001110111111100",
6443 => "010010011000110101011100",
6444 => "001101110101111001010000",
6445 => "000110111010000000101011",
6446 => "000000010011111110111011",
6447 => "111100001010110010110110",
6448 => "111001111010110111101001",
6449 => "111001110101101010001000",
6450 => "111101001011110011010001",
6451 => "000010011101101000110111",
6452 => "000111000101110010101000",
6453 => "001010001111101000000000",
6454 => "001100101111010010000000",
6455 => "010000000000110110110110",
6456 => "010011110001111000101000",
6457 => "010110100011001000110110",
6458 => "010111110101000000011110",
6459 => "010110110110111000000100",
6460 => "010011110001011100001010",
6461 => "010001000001010111011100",
6462 => "001111010100111110010000",
6463 => "001101100000101000011010",
6464 => "001011110000000010100000",
6465 => "001010101010001100110010",
6466 => "001010101001101011100100",
6467 => "001011001100111111000010",
6468 => "001010000101010101101011",
6469 => "000111101100111111001100",
6470 => "000111010110111000110101",
6471 => "001001000110001101000010",
6472 => "001010000000001011010110",
6473 => "001000001100111000000101",
6474 => "000011010001100100101111",
6475 => "111100011001011001100111",
6476 => "110101100011001101001111",
6477 => "101111010100001111000110",
6478 => "101001010001011111110100",
6479 => "100100000010001000001001",
6480 => "100001011110100101111001",
6481 => "100010110000100101000010",
6482 => "100111000011110100101111",
6483 => "101101000011100000000100",
6484 => "110100001000010000110011",
6485 => "111011100101011000000001",
6486 => "000001001111001110100111",
6487 => "000010001011101111001010",
6488 => "111110011011101011010101",
6489 => "111001001001011011011111",
6490 => "110100101011001101010000",
6491 => "110001110110110100101010",
6492 => "110000110001110111000010",
6493 => "110000011011011111010000",
6494 => "110000011001110001101100",
6495 => "110000110100001110111110",
6496 => "110001000001100001100100",
6497 => "110001011110110001000000",
6498 => "110010100111110101011110",
6499 => "110010101101010000110000",
6500 => "110001010001011100110000",
6501 => "101111101011101101011100",
6502 => "101101100111100101001110",
6503 => "101011000001110011100000",
6504 => "101010100000100001100110",
6505 => "101101110101101010010100",
6506 => "110011011011100111011110",
6507 => "111000101101110111101111",
6508 => "111101010110000001100010",
6509 => "000010110011011001010101",
6510 => "001001000011100110001000",
6511 => "001101101101000110111000",
6512 => "001111100000001100011100",
6513 => "010000000101001110011110",
6514 => "010000110001000111111000",
6515 => "010000101101001111101010",
6516 => "001110111111011011000110",
6517 => "001011101100000011100010",
6518 => "000111011110100100000010",
6519 => "000011111000111011111100",
6520 => "000010000010111101010100",
6521 => "000001100101101001010111",
6522 => "000001110111010111000011",
6523 => "000010101011100110010111",
6524 => "000100010110000011100101",
6525 => "000111011010010010000011",
6526 => "001011010111000010110000",
6527 => "001110100010011010100000",
6528 => "001111110101110001101010",
6529 => "001111100011111111000000",
6530 => "001110011110110011010100",
6531 => "001100101000011111110010",
6532 => "001001111001011101001000",
6533 => "000110110001000101111111",
6534 => "000011101010010100010101",
6535 => "000001000001110100001101",
6536 => "111111000111111110000100",
6537 => "111101000111111111011001",
6538 => "111010100101010010011000",
6539 => "111000011010100111101111",
6540 => "110111100010011101101001",
6541 => "110111110000101000100101",
6542 => "110111100111000110110101",
6543 => "110110011010111010001010",
6544 => "110101001110110010110010",
6545 => "110011101101100101111100",
6546 => "110001010010110111001110",
6547 => "101111111010010100001010",
6548 => "110000000100101000101010",
6549 => "110000010001010011111110",
6550 => "110000111101110001101100",
6551 => "110010101010001011000100",
6552 => "110100010101111110000010",
6553 => "110101101111100100010101",
6554 => "110110111101011100011100",
6555 => "111000001011100001011100",
6556 => "111001110011110011111001",
6557 => "111011010100000100111110",
6558 => "111100010011010011100110",
6559 => "111101000110111111011110",
6560 => "111101011110001111111101",
6561 => "111101011010111001000110",
6562 => "111110000110110100100001",
6563 => "000000011010010010000100",
6564 => "000011100001010010110111",
6565 => "000101101011011110001110",
6566 => "000110110001100100101001",
6567 => "000111110001001011101011",
6568 => "001000100100011000000111",
6569 => "001001111001000000100100",
6570 => "001101000010011100110010",
6571 => "010000100101110001100100",
6572 => "010010011110111100101000",
6573 => "010011000111011110101110",
6574 => "010011010100010011110000",
6575 => "010010010000000101010100",
6576 => "001110100100100001000100",
6577 => "001001010000111001100111",
6578 => "000101011100001101111111",
6579 => "000011011111110001000101",
6580 => "000000010100110110000110",
6581 => "111010011110101101101110",
6582 => "110100011010100001100101",
6583 => "110001110111100010111000",
6584 => "110011110101111111111100",
6585 => "110111100010011100100000",
6586 => "111010111100010001101100",
6587 => "111111010000011010101000",
6588 => "000100011011000100110110",
6589 => "000111100111110100001000",
6590 => "000111111010110111000011",
6591 => "000111111110000101000000",
6592 => "001010000110000101000010",
6593 => "001100101111001100100110",
6594 => "001100110010010111111010",
6595 => "001011001111000010001010",
6596 => "001100001001011110100000",
6597 => "001111011101011010001100",
6598 => "010001000011001001101100",
6599 => "001111111010100111011100",
6600 => "001110111011100000100000",
6601 => "001111100000010110110110",
6602 => "001111111111110111110100",
6603 => "001110011011100101000010",
6604 => "001010111101100011001001",
6605 => "000111001010100001100110",
6606 => "000011101100011111000000",
6607 => "000000101101100101000110",
6608 => "111110101000011000111011",
6609 => "111100010100010001000111",
6610 => "111000000000101101101101",
6611 => "110010100110101011000010",
6612 => "101110100000100000011100",
6613 => "101100011010010110011110",
6614 => "101011010100110010111110",
6615 => "101010101101100000111000",
6616 => "101011101000000110011100",
6617 => "101110111110101011000100",
6618 => "110011010101111100001110",
6619 => "110111100010000100000000",
6620 => "111101010111011110101110",
6621 => "000100101110001001001110",
6622 => "001000100001001110110000",
6623 => "000110101001100100111100",
6624 => "000011001011111001100111",
6625 => "000000011001100010111011",
6626 => "111101100010011001111100",
6627 => "111100000101111011100110",
6628 => "111101001001000000010010",
6629 => "111101110101011010011110",
6630 => "111011001110000001001011",
6631 => "110110001101000000010100",
6632 => "110010011010100110010110",
6633 => "110001001001001001101000",
6634 => "110000010001101101100010",
6635 => "101111100010100010111100",
6636 => "110000001000011011110000",
6637 => "110000111101000011011010",
6638 => "110001101011011110111000",
6639 => "110011110100001010011100",
6640 => "110111011011001010100000",
6641 => "111100001001101100100011",
6642 => "000001101011111111000100",
6643 => "000110100101100000110110",
6644 => "001010001001010010101001",
6645 => "001100011001101000111100",
6646 => "001100110101010011101010",
6647 => "001011011000100110100011",
6648 => "001000101001101011110110",
6649 => "000110001111001100011011",
6650 => "000110001100000111110111",
6651 => "000111100101000111000000",
6652 => "000111010110101111110001",
6653 => "000101000111100100000011",
6654 => "000011011100011111111110",
6655 => "000100000011000101100110",
6656 => "000101001100011101100110",
6657 => "000100001110111101101110",
6658 => "000001110111110100111001",
6659 => "000000101101001010100000",
6660 => "000001011001001011110010",
6661 => "000010100011101100100001",
6662 => "000010100010110011011001",
6663 => "000001011001011110010000",
6664 => "000000110100011011101110",
6665 => "000001100010001100100001",
6666 => "000010110111111100001110",
6667 => "000100000011111000010001",
6668 => "000100101111000111000101",
6669 => "000101010011011111100100",
6670 => "000101100100010111000010",
6671 => "000100010001100000010010",
6672 => "000001011011101000001101",
6673 => "111101111000100111101010",
6674 => "111001101110110001111100",
6675 => "110101100011110011010100",
6676 => "110010000110011011110010",
6677 => "101111000000000110101000",
6678 => "101100010100100101110010",
6679 => "101011000010101110110100",
6680 => "101011100000100000101000",
6681 => "101101001001110011011010",
6682 => "101111011011001001100000",
6683 => "110001111000110100000010",
6684 => "110100001001100100100100",
6685 => "110110011101001001110010",
6686 => "111000111010100010011001",
6687 => "111010100110011000110111",
6688 => "111011010010001101110100",
6689 => "111011100101011001000000",
6690 => "111011011011111001111010",
6691 => "111011011100101111000010",
6692 => "111100100010001110001110",
6693 => "111101111101001001001110",
6694 => "111111100110010111111111",
6695 => "000010010111011100111011",
6696 => "000101001011000111110011",
6697 => "000110100010000110110010",
6698 => "000111001100111000010100",
6699 => "001000100001111110101011",
6700 => "001010011000100111010110",
6701 => "001011110010111101100101",
6702 => "001100101111101001100100",
6703 => "001101010101101011011010",
6704 => "001100111010011110001010",
6705 => "001100011001100011000110",
6706 => "001101100001101011101110",
6707 => "001111100110011000110000",
6708 => "010001011000101011011110",
6709 => "010010111110000110101000",
6710 => "010100001101001010011000",
6711 => "010100001000000101001010",
6712 => "010001011111010000101000",
6713 => "001100110101001111101110",
6714 => "001000101011010101111101",
6715 => "000101101000010000011100",
6716 => "000010010010111110000111",
6717 => "111101100011000101000111",
6718 => "110110111101110101101010",
6719 => "110001100000010000111100",
6720 => "110000111100001110010100",
6721 => "110011100011010101010010",
6722 => "110110101001000011011000",
6723 => "111010110010001100010100",
6724 => "111110110010001011110111",
6725 => "000000010110001101110010",
6726 => "000000010111001111100001",
6727 => "000001010000110101110000",
6728 => "000100011000000011111111",
6729 => "001000000111011110101010",
6730 => "001001010010111101110010",
6731 => "000111111010001000111111",
6732 => "000110111100110101101011",
6733 => "001000001000110110010111",
6734 => "001001110010100111010100",
6735 => "001000110011010010001100",
6736 => "000101101000111000110110",
6737 => "000011101001110001111010",
6738 => "000011011001111001010011",
6739 => "000010111100101000100100",
6740 => "000000100000101111110000",
6741 => "111011110110100100010100",
6742 => "110111100101101011101100",
6743 => "110101011100111110100111",
6744 => "110100000000010011010011",
6745 => "110010010001011001011010",
6746 => "101111000111010000100010",
6747 => "101010000000001011100100",
6748 => "100111001100011000001010",
6749 => "101000111100010000100000",
6750 => "101010101010001010100010",
6751 => "101010011010100000011000",
6752 => "101011100010010011101100",
6753 => "101111101011001010110000",
6754 => "110110101101111101001000",
6755 => "111111101010000011001111",
6756 => "000111000100001011001110",
6757 => "001011010000001011110100",
6758 => "001110000110010101111010",
6759 => "001111101100010000010110",
6760 => "001110000111111110110010",
6761 => "001010011111001101001001",
6762 => "000111110110110110011011",
6763 => "000110101100000011010000",
6764 => "000100011111111100100000",
6765 => "111111100010011001100011",
6766 => "111001100100101110011000",
6767 => "110101011011000110111010",
6768 => "110011001010000010001110",
6769 => "110001111011000001010110",
6770 => "110010001100001111101110",
6771 => "110100000001101000110001",
6772 => "110110111000110101100011",
6773 => "111010010110000010101111",
6774 => "111101011100111110100111",
6775 => "111111111101011010010010",
6776 => "000010101010011101110101",
6777 => "000110000011000100011010",
6778 => "001010101100111011100111",
6779 => "010000011000000100101010",
6780 => "010100101010000100000010",
6781 => "010110011101101000011000",
6782 => "010111110010011111001010",
6783 => "011001010100010111111101",
6784 => "011001000001001011010011",
6785 => "010110011000000111011000",
6786 => "010011011100101000010000",
6787 => "010001001000010001111100",
6788 => "001110000111101001101010",
6789 => "001001100101001100010010",
6790 => "000100110000000110101110",
6791 => "000001111101001001101111",
6792 => "000001100010110001010000",
6793 => "000001010010101100001100",
6794 => "000000110111110110111010",
6795 => "000010010101000111001010",
6796 => "000101011000010010101011",
6797 => "000111111111110100011100",
6798 => "001001000110101010001000",
6799 => "001000010000010010001001",
6800 => "000110101110001111111111",
6801 => "000110000010110101010010",
6802 => "000100101110110100010100",
6803 => "000001111011011100011111",
6804 => "111111101000111010010001",
6805 => "111110000100010011000111",
6806 => "111011110101010101011111",
6807 => "111001100100010001001000",
6808 => "111000010000001001100011",
6809 => "110111011011011011001010",
6810 => "110110010100001111000011",
6811 => "110100100100100111100000",
6812 => "110010011110100000000010",
6813 => "110000010011010010101000",
6814 => "101101101010100101100100",
6815 => "101010101011101111011010",
6816 => "101000010010111000111000",
6817 => "100110110010000000000111",
6818 => "100101110100000000011101",
6819 => "100101011100010011001101",
6820 => "100101101000100110010101",
6821 => "100110100011000000010111",
6822 => "101001100011100110110110",
6823 => "101111000100000011101000",
6824 => "110100100011010101010101",
6825 => "111000000110100110110000",
6826 => "111010110001100101000010",
6827 => "111101010101001111000011",
6828 => "111111000000001101000000",
6829 => "000000000010000110110010",
6830 => "000001011010000000010100",
6831 => "000010110010001101001000",
6832 => "000011001100111010100000",
6833 => "000010101010101010111111",
6834 => "000010001010101100110000",
6835 => "000010111001111110011101",
6836 => "000101101001110001110000",
6837 => "001001111100011010110000",
6838 => "001101110011000000010000",
6839 => "010000000001110001001100",
6840 => "010010011010010101110100",
6841 => "010110010010000010000110",
6842 => "011001100010000110110011",
6843 => "011010110011010000000010",
6844 => "011011001101110011101000",
6845 => "011010011010101000010110",
6846 => "010111110101110000100100",
6847 => "010101000111100100110010",
6848 => "010001111111110110001010",
6849 => "001100110000010011110110",
6850 => "000111100001101011101010",
6851 => "000101011011011101100011",
6852 => "000100111011110011101010",
6853 => "000010100001100110101100",
6854 => "111110001111100000110011",
6855 => "111011101011100111001111",
6856 => "111100110111001001001000",
6857 => "111111110011100011110101",
6858 => "000010010100110110001010",
6859 => "000100001011101011110010",
6860 => "000100111000001001010000",
6861 => "000011011000010000101110",
6862 => "000000000110001011111101",
6863 => "111101101101010110111000",
6864 => "111110111010011000001111",
6865 => "000010000111011100111101",
6866 => "000011000100010101101000",
6867 => "000001100101000101111111",
6868 => "000000111111011101011111",
6869 => "000010100000100110110000",
6870 => "000100100001000100111100",
6871 => "000100100100011000001000",
6872 => "000001101111001000011000",
6873 => "111110101001010010110110",
6874 => "111101110000010010110010",
6875 => "111100111010000011011010",
6876 => "111000111000000010111110",
6877 => "110010001010001110110000",
6878 => "101011110110110001111110",
6879 => "101000001011111011011100",
6880 => "100110010111010011000100",
6881 => "100100010001101001111111",
6882 => "100010001010101001010110",
6883 => "100001101011001110010111",
6884 => "100011000111110011011100",
6885 => "100110010110111011011011",
6886 => "101010001010100111110010",
6887 => "101011110101011100111000",
6888 => "101100010111111110000000",
6889 => "110000011001010110101110",
6890 => "110111001011101110000100",
6891 => "111011000001001101001100",
6892 => "111011011111010111110010",
6893 => "111101001100101100101101",
6894 => "000000001100001001110001",
6895 => "000000011100001010101100",
6896 => "111101111111111111000011",
6897 => "111100011011010001001110",
6898 => "111100010101011110101011",
6899 => "111011100101011101001010",
6900 => "111001011111100111111011",
6901 => "110111000000001111011101",
6902 => "110100001011111110001100",
6903 => "110000010101111001111100",
6904 => "101100110010010111111000",
6905 => "101100100000001110010100",
6906 => "101111110100011010110100",
6907 => "110100001010100011010100",
6908 => "110111110010010111110100",
6909 => "111010010010100110011110",
6910 => "111100000101101001000101",
6911 => "111110110011000110001000",
6912 => "000011101101110011011110",
6913 => "001010010011010010111010",
6914 => "010000011000010100000010",
6915 => "010100000100001111110110",
6916 => "010110110010001001011110",
6917 => "011010111001101000001011",
6918 => "011110100011001101001000",
6919 => "011110101110111100000011",
6920 => "011100100000001011111011",
6921 => "011010000111100000011011",
6922 => "010111101111110111111010",
6923 => "010100111110100100011010",
6924 => "010001110110110100111010",
6925 => "001110100101101110011000",
6926 => "001011111001101110110000",
6927 => "001010111100011010000001",
6928 => "001011110011011011111001",
6929 => "001100110111101001111000",
6930 => "001100100110010110110100",
6931 => "001011010101100001111110",
6932 => "001010111011100110000000",
6933 => "001100010101101101101010",
6934 => "001110001001010100110000",
6935 => "001110111110111111010100",
6936 => "001111001010011111000110",
6937 => "001110110000010100101010",
6938 => "001110001010010111010100",
6939 => "001110101000101011101010",
6940 => "001111001011001100110100",
6941 => "001101111101000010001100",
6942 => "001011100010010000100101",
6943 => "001000011001000011001010",
6944 => "000100001110011100101010",
6945 => "111111111001000011111000",
6946 => "111011101010001010111000",
6947 => "110110110110110000101001",
6948 => "110001100111111010110110",
6949 => "101100010110111111010110",
6950 => "100111110100010000000111",
6951 => "100101011111110101100010",
6952 => "100101110101000000011101",
6953 => "100111100110011001100010",
6954 => "101001010010110101000010",
6955 => "101010000100100100111100",
6956 => "101010001111100011111010",
6957 => "101010110000110101000100",
6958 => "101011111111011110011010",
6959 => "101101011100111111100000",
6960 => "101110110110011101111000",
6961 => "110000001110010101011000",
6962 => "110001001110111111111000",
6963 => "110010010110110110100000",
6964 => "110101010010010100101010",
6965 => "111010000110111100001010",
6966 => "111111000010001111010110",
6967 => "000010111100100111011010",
6968 => "000101011100011011001100",
6969 => "000110011000010101010010",
6970 => "000110000110010011011010",
6971 => "000100110100010000000101",
6972 => "000011001111000100111000",
6973 => "000010110010011010111000",
6974 => "000011110000010011111010",
6975 => "000101001100001101110101",
6976 => "000110100111110100010010",
6977 => "001000011000111100011110",
6978 => "001011010010011101010111",
6979 => "001111101111000111001000",
6980 => "010100010011100111101100",
6981 => "010110101111000111111010",
6982 => "010111000010111011001110",
6983 => "010110011001111101111010",
6984 => "010011110111110000000010",
6985 => "001111000010000001000010",
6986 => "001010011001001001000010",
6987 => "000111011010000110000110",
6988 => "000100111011000101001100",
6989 => "000001011010011100101001",
6990 => "111100110100111110100111",
6991 => "111010011000011110110000",
6992 => "111100101010111001100110",
6993 => "000001001011011111010100",
6994 => "000101100011110100100101",
6995 => "001001111101000000001010",
6996 => "001100110100011110011100",
6997 => "001101000100000000010000",
6998 => "001011110000100100101000",
6999 => "001010000011010110100101",
7000 => "001001101000100011011100",
7001 => "001010000001010101111011",
7002 => "000111111111111101011001",
7003 => "000100011010010100110100",
7004 => "000011000100100101000001",
7005 => "000100010010011000100011",
7006 => "000101101110111010111111",
7007 => "000101101000010011001101",
7008 => "000100101010000110001000",
7009 => "000100101010010111000010",
7010 => "000100100000111001100010",
7011 => "000010000101100100110000",
7012 => "111101010001110111010100",
7013 => "110110011110111011001000",
7014 => "101111110110111011111110",
7015 => "101100001000101011000110",
7016 => "101001111100001101111100",
7017 => "100111001000110011011011",
7018 => "100100101111100010111001",
7019 => "100100000011001110010111",
7020 => "100101010101010101010100",
7021 => "101000001101100111111110",
7022 => "101011001100111100000110",
7023 => "101100111110101110001010",
7024 => "101110000101100010001110",
7025 => "110000101010001100110110",
7026 => "110101000100011111001000",
7027 => "111000101010110001111101",
7028 => "111010110000100011110011",
7029 => "111101001100101011101101",
7030 => "111111001010110010101110",
7031 => "111110101011111101001000",
7032 => "111100100100101101101100",
7033 => "111010010101111011101000",
7034 => "111000000111100000110101",
7035 => "110101010100000000110000",
7036 => "110001010101010010011100",
7037 => "101100101010011011101100",
7038 => "101001001110100001111110",
7039 => "101000010001111111010110",
7040 => "101000100101100010101000",
7041 => "101001000011101010001010",
7042 => "101011101010111111111010",
7043 => "110001100011101010011010",
7044 => "110111100010100010100111",
7045 => "111010101111001001100010",
7046 => "111100000100110101111101",
7047 => "111101101000100101111110",
7048 => "000000010010011001010101",
7049 => "000011100111011101011100",
7050 => "000110100101001111011010",
7051 => "001000111110000000000011",
7052 => "001011110010100010000010",
7053 => "001111010101101100100000",
7054 => "010001111111100010000000",
7055 => "010010001101010001101100",
7056 => "010000000010100101011110",
7057 => "001100100011100010011110",
7058 => "001001101011100010001101",
7059 => "001000010110111101011001",
7060 => "000110111100010011101100",
7061 => "000101000011011001001100",
7062 => "000101000010000010100010",
7063 => "000111100010001100000111",
7064 => "001011000000100100101001",
7065 => "001110001000010110100000",
7066 => "010000100000011011011000",
7067 => "010011001110100011001010",
7068 => "010110100010101100010100",
7069 => "011000010101000010010100",
7070 => "011000010100011101001001",
7071 => "011000100010010010111111",
7072 => "011000110010111110100010",
7073 => "010111101100001110011010",
7074 => "010101101101111101010010",
7075 => "010100001010111101110000",
7076 => "010011001111000111011010",
7077 => "010001110101010001011000",
7078 => "001111000111000010100110",
7079 => "001011111010101111111111",
7080 => "001001000111000010001110",
7081 => "000101101000000011101100",
7082 => "000001000010001001100100",
7083 => "111101011100111110100000",
7084 => "111011110100101010100001",
7085 => "111010001011110100110001",
7086 => "110111101011011010111101",
7087 => "110101001110100010001001",
7088 => "110011001010001000000100",
7089 => "110010000010100101011000",
7090 => "110010001110011000111010",
7091 => "110010011000101100011000",
7092 => "110010000100100000001000",
7093 => "110010011111100011001000",
7094 => "110100001100110101000100",
7095 => "110110101011101100011111",
7096 => "111000110110011100001110",
7097 => "111010011011001111011001",
7098 => "111100100010100010010000",
7099 => "111110110001001100011100",
7100 => "111111110010100110001101",
7101 => "000000101110101100101101",
7102 => "000010001011110111001001",
7103 => "000010010000110111011111",
7104 => "000000100011001011110100",
7105 => "111110011000001011101100",
7106 => "111100010001010010110000",
7107 => "111010110100011001101110",
7108 => "111011001100000011010000",
7109 => "111101100110010001011111",
7110 => "000001000110000010101010",
7111 => "000100110000111000111110",
7112 => "001000010110100111100100",
7113 => "001011011111010101100010",
7114 => "001101011100001000001000",
7115 => "001110000000100011000010",
7116 => "001101010101110000100100",
7117 => "001011101001010001010001",
7118 => "001001111110000001101001",
7119 => "001001001100101001110111",
7120 => "001000001110001011011100",
7121 => "000101100101111111000011",
7122 => "000010100011111011010010",
7123 => "000001100100001101100000",
7124 => "000010001111110100101101",
7125 => "000010000010100001100010",
7126 => "111111110000101110010100",
7127 => "111100010001101100100010",
7128 => "111001010011000111011000",
7129 => "111000001010001100010001",
7130 => "111000011011001110010110",
7131 => "111000111100100000111001",
7132 => "111001101001110001110001",
7133 => "111010011101101000110010",
7134 => "111010101111000011001100",
7135 => "111011000011110110011101",
7136 => "111101010100110000100011",
7137 => "000001111010001110110011",
7138 => "000101111000011110111011",
7139 => "000110100100011110111110",
7140 => "000101111101010010111100",
7141 => "000110111011110010001100",
7142 => "001000010101000011001100",
7143 => "000111111010011011011111",
7144 => "000101001110100011000100",
7145 => "000000111001010001110010",
7146 => "111100111011100101011110",
7147 => "111010000101011100111110",
7148 => "110101101101110001100110",
7149 => "101110111011100100010100",
7150 => "101001000010000001010110",
7151 => "100110111101100011010100",
7152 => "101001000010000110111110",
7153 => "101101100110100100001110",
7154 => "110010001110110110000010",
7155 => "110101111110011010011110",
7156 => "111001011101011011100101",
7157 => "111100111100100000101100",
7158 => "111111110111100001001001",
7159 => "000000101101010011100001",
7160 => "111101100110010101001101",
7161 => "110111110111011111001000",
7162 => "110101000101100101101000",
7163 => "110111111011010010101000",
7164 => "111011110110101010101101",
7165 => "111110000110010101010011",
7166 => "000010001010111100111111",
7167 => "000111110000101001000010",
7168 => "001001001101101110101010",
7169 => "000101110101011101001110",
7170 => "000001011011000110011101",
7171 => "111101010100000000001010",
7172 => "111000100101110101111101",
7173 => "110010110110101001101000",
7174 => "101101100110110111010010",
7175 => "101010100001000000100100",
7176 => "101000100110111100011000",
7177 => "100111111110111101101110",
7178 => "101011001111011111001010",
7179 => "110001000111100101101010",
7180 => "110101010010000100111000",
7181 => "110110111110111011000100",
7182 => "111000010101100111101101",
7183 => "111010101100100000011011",
7184 => "111101011000011100011000",
7185 => "111110110011100010111101",
7186 => "000000000000000101111011",
7187 => "000010111101001111011011",
7188 => "000101110111000011101101",
7189 => "000110111100011111110101",
7190 => "001000000011100010010010",
7191 => "001001000101000110011010",
7192 => "000111001000011010111100",
7193 => "000010101101011100111011",
7194 => "111111000111110111001010",
7195 => "111101110101101100100110",
7196 => "111110001011011000011100",
7197 => "111110100101100111001111",
7198 => "111110101010000000010101",
7199 => "000000011110101100110010",
7200 => "000100111001000001101111",
7201 => "001001001111001010111111",
7202 => "001011011111010111011110",
7203 => "001100000101100111010110",
7204 => "001100001111011011100000",
7205 => "001100111011011101100000",
7206 => "001101000011110001000100",
7207 => "001010110000110001001111",
7208 => "000111101010001000011000",
7209 => "000110001001101001011010",
7210 => "000101011000000010011101",
7211 => "000100101111000110010010",
7212 => "000101000001110010101110",
7213 => "000101010010001110010111",
7214 => "000100110100101110111000",
7215 => "000100101011010011001110",
7216 => "000100001111101110011001",
7217 => "000010010001001010111101",
7218 => "111111011110011110111111",
7219 => "111100101001011000100101",
7220 => "111010010000010001010000",
7221 => "111001011000111001101001",
7222 => "111001100101100010101010",
7223 => "111001101111011100101110",
7224 => "111010101000111101101000",
7225 => "111100011110010100000010",
7226 => "111110000010000010011001",
7227 => "111111001100000111110101",
7228 => "000000000101100100100000",
7229 => "000000111010011111101100",
7230 => "000010110100111001000110",
7231 => "000101010100011000111011",
7232 => "000110011101111110010001",
7233 => "000110101000000010111111",
7234 => "000111001101000011101010",
7235 => "001000100000111000110100",
7236 => "001010101100010111110011",
7237 => "001101000110110001011000",
7238 => "001110001110000000000110",
7239 => "001101111000100011000000",
7240 => "001100111000001110000010",
7241 => "001011000110011111001010",
7242 => "001000101101010110001001",
7243 => "000110110110101010001101",
7244 => "000110010111000001001001",
7245 => "000111011000101000001011",
7246 => "001001100011001001100010",
7247 => "001100001011100000011100",
7248 => "001111011101000101111010",
7249 => "010011001100001011111010",
7250 => "010101110100000011101010",
7251 => "010111011111111111010110",
7252 => "011001100001001100011101",
7253 => "011010010001100110010011",
7254 => "011000101001101001101101",
7255 => "010110101100010001001000",
7256 => "010100110000000111011100",
7257 => "010000111110101010100110",
7258 => "001011001111011010111100",
7259 => "000101001111110010000110",
7260 => "000001000010001001110000",
7261 => "111110000111101111111010",
7262 => "111000101011110000011000",
7263 => "110000001111111011101110",
7264 => "101010010010000111111010",
7265 => "101001111110010001101010",
7266 => "101100010101101100011000",
7267 => "101110000101111110010110",
7268 => "101111010101001001010000",
7269 => "110000111001101000001100",
7270 => "110010000001000001000110",
7271 => "110001111001010011111110",
7272 => "110010010110001011101100",
7273 => "110101100010100000100110",
7274 => "111001000100000001111011",
7275 => "111001000001011001111001",
7276 => "110111101100011101000011",
7277 => "111001101110110000010001",
7278 => "111110001000000000000111",
7279 => "000001000110011010011011",
7280 => "000000011101010111011101",
7281 => "111100011011001011101110",
7282 => "111000100010000100111011",
7283 => "110101100010001010010110",
7284 => "101111000111001111000100",
7285 => "100110011110111100100001",
7286 => "100001111100010000111001",
7287 => "100001110011101010010100",
7288 => "100010101100000011010011",
7289 => "100011011101001110101101",
7290 => "100100100110101000001111",
7291 => "101000010100101011100010",
7292 => "101111111110011000100100",
7293 => "111001110011001100001110",
7294 => "000011011110010101100101",
7295 => "001001110000000101000001",
7296 => "001010010001110010001011",
7297 => "001000101001001111011011",
7298 => "001001000001011111111010",
7299 => "001001101101001110110010",
7300 => "001000101000100010110110",
7301 => "000111101011100000000011",
7302 => "001000011111101100011010",
7303 => "001001101010101111011101",
7304 => "001000111001000101101010",
7305 => "000101101101111000100111",
7306 => "000001110001101010101000",
7307 => "111111000110111011000001",
7308 => "111110000000010110110011",
7309 => "111100111100000010011001",
7310 => "111011100101010011110111",
7311 => "111011001011011100111110",
7312 => "111011110010001000100100",
7313 => "111101000110000110000101",
7314 => "111111100101011111011010",
7315 => "000010101101010101011110",
7316 => "000101010001011010010100",
7317 => "000110101010011101101000",
7318 => "000110111011010001010010",
7319 => "000111010110011001010101",
7320 => "001000111000100110000010",
7321 => "001010110010001110100000",
7322 => "001100101101011010100000",
7323 => "001110110011001111000110",
7324 => "010000010001110111111000",
7325 => "010000010110011010101110",
7326 => "001110100011100110101000",
7327 => "001011000101001110011010",
7328 => "000111000010000100011000",
7329 => "000010011001100010011001",
7330 => "111100110100111011010110",
7331 => "111000101000011000110110",
7332 => "111000000100011110110000",
7333 => "111001101011010111101111",
7334 => "111011000010101101010010",
7335 => "111100011010001000010101",
7336 => "111111100111000001010100",
7337 => "000100100101101000001010",
7338 => "001000010100000100001101",
7339 => "001000111001010100010010",
7340 => "001000100101110000000011",
7341 => "001000111110100101111100",
7342 => "000111011010011001111010",
7343 => "000010101010000101100100",
7344 => "111101110011001001110011",
7345 => "111010100110000011101000",
7346 => "111000000011011100011101",
7347 => "110110011001011011000010",
7348 => "110110001001110101010101",
7349 => "110110010001100100101100",
7350 => "110110001110011010010110",
7351 => "110110001110111100010100",
7352 => "110110000010000010010010",
7353 => "110101011101100110110010",
7354 => "110100001111100000101010",
7355 => "110001111110000011000110",
7356 => "101111110101000011000110",
7357 => "101111011100110110101010",
7358 => "110000000100011100100000",
7359 => "101111110110110011101110",
7360 => "101111001000101101101100",
7361 => "101111100101101110011000",
7362 => "110001001011111110000100",
7363 => "110010100101111001000100",
7364 => "110011101000111101010110",
7365 => "110100111001101010100110",
7366 => "110110100010000011100010",
7367 => "111000110111010111110001",
7368 => "111011101101101101100000",
7369 => "111101110100100010000101",
7370 => "111110111011010000001010",
7371 => "000000001100011011101100",
7372 => "000010000000100111001100",
7373 => "000011101100101100101111",
7374 => "000101001001101011100010",
7375 => "000110110110010110111100",
7376 => "001000101010110100010100",
7377 => "001010001111010010010011",
7378 => "001011110110000110110010",
7379 => "001110001001111110010110",
7380 => "010010010010011000100100",
7381 => "011000010010010101110100",
7382 => "011100101111110001010101",
7383 => "011101001010001100011111",
7384 => "011100001011010110011111",
7385 => "011011111000110101111101",
7386 => "011011000010010001000111",
7387 => "011001111011111100101000",
7388 => "011001110101101011001101",
7389 => "011010010000101100111001",
7390 => "011010100110100010111101",
7391 => "011010000100000010011111",
7392 => "011000100110101011001011",
7393 => "011000000011001001110011",
7394 => "010111100110101100111010",
7395 => "010100010110010010011110",
7396 => "001111101011000110000110",
7397 => "001100100110101001101110",
7398 => "001001010111100000001000",
7399 => "000010011010010101101110",
7400 => "111000010001001011110011",
7401 => "101111010000010100001000",
7402 => "101011001111010001110010",
7403 => "101100101001100101100110",
7404 => "110001000000000111111000",
7405 => "110101011000001101110110",
7406 => "111000010101100110000101",
7407 => "111010011101000000010101",
7408 => "111101010100100111101011",
7409 => "000001010000101110011100",
7410 => "000100100110111000001100",
7411 => "000101110110010001001100",
7412 => "000100010011101000011101",
7413 => "000000001101100010100110",
7414 => "111100000010110101010111",
7415 => "111000001101000111111011",
7416 => "110000011110010110011100",
7417 => "100110010000000110111001",
7418 => "100001101000111101111111",
7419 => "100010111000001111110111",
7420 => "100011011001100101110111",
7421 => "100010011011000101010111",
7422 => "100010100101100101110111",
7423 => "100011100110100101011110",
7424 => "100100010010000100110101",
7425 => "100101010001001101110010",
7426 => "101000110011000001110010",
7427 => "101110011110001100101110",
7428 => "110010011101010011011110",
7429 => "110100010100000100100100",
7430 => "110110011101110010110110",
7431 => "111000010000011100101100",
7432 => "111000110010101001100111",
7433 => "111001010010110110001010",
7434 => "111010110000001011000101",
7435 => "111110010010110111010111",
7436 => "000011011011000000011000",
7437 => "000110111001011100111000",
7438 => "000111110000000100010011",
7439 => "000111011100110011000100",
7440 => "000101100011110111001100",
7441 => "000001000000011001110000",
7442 => "111010010101111011111010",
7443 => "110011101010111100011110",
7444 => "110000011010110100101110",
7445 => "110001110101101110111000",
7446 => "110100101000010011001011",
7447 => "110110011001111011100110",
7448 => "111001001000110101011110",
7449 => "111110000001000000011100",
7450 => "000011011111010100101111",
7451 => "001001001101000110101000",
7452 => "001111001111101001100010",
7453 => "010011101111110100010110",
7454 => "010101101100001000010110",
7455 => "010101111111111110101100",
7456 => "010101010100100110100100",
7457 => "010100000001101101011010",
7458 => "010010011100111100101110",
7459 => "010000011111001101000000",
7460 => "001110101001111010110100",
7461 => "001101111110110100010000",
7462 => "001110100000110101111110",
7463 => "001111001011100000011010",
7464 => "001110101111001100010110",
7465 => "001101010100011110001110",
7466 => "001100100101101101010000",
7467 => "001101011101001101110110",
7468 => "001111000110101101100110",
7469 => "001111111011111111110110",
7470 => "001110101011011101011100",
7471 => "001100000001100100001110",
7472 => "001010010101011100000100",
7473 => "001010100001100101001011",
7474 => "001011001101000000011110",
7475 => "001011000001111110111001",
7476 => "001010011101000001001011",
7477 => "001010110110111110110011",
7478 => "001011111100110011111101",
7479 => "001011011010110101110011",
7480 => "001000010010111111111000",
7481 => "000100001100101000001111",
7482 => "000000101101100000111111",
7483 => "111101110101110101100001",
7484 => "111010110011011101001100",
7485 => "110111001011101101100110",
7486 => "110011010010011011010010",
7487 => "101111101000110100101110",
7488 => "101100100001111000101110",
7489 => "101001110011111111000100",
7490 => "100111000101101011010111",
7491 => "100100111000010111101110",
7492 => "100100011000001011111101",
7493 => "100101101010010000100001",
7494 => "100111100100011101111100",
7495 => "101000101010010000010100",
7496 => "101000011101011100110010",
7497 => "101000001110010110110110",
7498 => "101000100101011000010000",
7499 => "101000100101110011010010",
7500 => "101000011101000101011010",
7501 => "101000111010111100000010",
7502 => "101001100000011111101100",
7503 => "101010101011111011100110",
7504 => "101101100010111001110000",
7505 => "110001001100111101010100",
7506 => "110100011001101000001011",
7507 => "110111010001011010100000",
7508 => "111010000011111110111110",
7509 => "111100011110110000100101",
7510 => "111110011101010000110010",
7511 => "000000010110100011111010",
7512 => "000010010001000010110001",
7513 => "000100000000100000010001",
7514 => "000101010100110101001101",
7515 => "000101110110001111001110",
7516 => "000110110110010111010010",
7517 => "001010100100100111010100",
7518 => "001111101001101100010010",
7519 => "010011000101010010110100",
7520 => "010101100001000001110000",
7521 => "011000100001011110100101",
7522 => "011011011111100100101110",
7523 => "011101100101000010100000",
7524 => "011110011011110010100110",
7525 => "011110010010000111111011",
7526 => "011101101011110101110011",
7527 => "011100101110010111110101",
7528 => "011011110011111100001011",
7529 => "011011001010010111100011",
7530 => "011010011110100100001000",
7531 => "011001111000100001101100",
7532 => "011000010000110000111001",
7533 => "010101000111100010101110",
7534 => "010010101111111101111000",
7535 => "001111110010010000010110",
7536 => "001000100011000010010000",
7537 => "000000111111011001110010",
7538 => "111111001011110000110010",
7539 => "000001011001011111011100",
7540 => "000011010100000100001001",
7541 => "000100100010110110001010",
7542 => "000110110001011011010001",
7543 => "001001101010100100111000",
7544 => "001010101011110000010100",
7545 => "001001111011001011011100",
7546 => "001010000011001111001011",
7547 => "001010010011011111110010",
7548 => "000111001001110101011101",
7549 => "000000000000101001010001",
7550 => "111000101010010100111000",
7551 => "110100000011111011000010",
7552 => "101111000110111001010000",
7553 => "100111010011010011110111",
7554 => "100001101100010010111010",
7555 => "100001011101010011101011",
7556 => "100010100001111100101100",
7557 => "100010100110111100111111",
7558 => "100010110100100011011101",
7559 => "100011101101000000100101",
7560 => "100110111111000000111111",
7561 => "101110000000100011010110",
7562 => "110110100011101000010111",
7563 => "111110001000110010111000",
7564 => "000011111001111101110000",
7565 => "000111001010100110100111",
7566 => "001000011100000000001100",
7567 => "001001100000010010001110",
7568 => "001001111011011111011101",
7569 => "000111001000111010010011",
7570 => "000001001100000101110011",
7571 => "111011001001110010111111",
7572 => "110110011110000101110000",
7573 => "110001111111111101011110",
7574 => "101101010000110111111010",
7575 => "101010000011100011001110",
7576 => "101010010010001111011000",
7577 => "101100110011011011000100",
7578 => "101111001001100100111010",
7579 => "110001101000010011011100",
7580 => "110101011010110010010100",
7581 => "111001010100001011010010",
7582 => "111011011011111100000011",
7583 => "111011100010000111011111",
7584 => "111011011110001111111000",
7585 => "111101000000101011001001",
7586 => "111111000101011010010110",
7587 => "000001001111011111000110",
7588 => "000101111011111001101100",
7589 => "001100101010000111011110",
7590 => "010001001100111000001010",
7591 => "010010100001010011110100",
7592 => "010010110001010001100010",
7593 => "010010001101001001000000",
7594 => "001111010101110001001000",
7595 => "001010011100100100101101",
7596 => "000101111001110100110100",
7597 => "000010110111000101101000",
7598 => "000000001110001101100001",
7599 => "111101111110010110111010",
7600 => "111110000000011111101000",
7601 => "000000111000110010011000",
7602 => "000100100101101011110110",
7603 => "000111001111010111111010",
7604 => "001010001010101100100110",
7605 => "001111101110000010100100",
7606 => "010110001101100101011000",
7607 => "011001101111111101110000",
7608 => "011001111010111001011101",
7609 => "011001000011111000000101",
7610 => "011000011011111110011011",
7611 => "010111011011111111010010",
7612 => "010100110001100100101010",
7613 => "010000110011101100000000",
7614 => "001101100000100011111010",
7615 => "001011010111000011010010",
7616 => "001001011001000001101111",
7617 => "000111001111111100000110",
7618 => "000100110101000110100001",
7619 => "000010001001011011110000",
7620 => "111111110111011100000000",
7621 => "111110110001001110011101",
7622 => "111110110100000001111111",
7623 => "111101111111100100111110",
7624 => "111010011110101001100000",
7625 => "110110000110101011010100",
7626 => "110010110111010000001000",
7627 => "101111010111001111110000",
7628 => "101011010000010111101010",
7629 => "101000110101000000001110",
7630 => "101001000011110010111010",
7631 => "101010110001100100011010",
7632 => "101100000100110010010010",
7633 => "101100011011000000111000",
7634 => "101101101010101111111010",
7635 => "110000011101011111101100",
7636 => "110010110101000101011010",
7637 => "110011010111010011010000",
7638 => "110010001000100110001000",
7639 => "110000100010110100110000",
7640 => "101111111101101010101000",
7641 => "101110101110100010100110",
7642 => "101011011110011000101010",
7643 => "101000111000011100101110",
7644 => "101000101111000001101010",
7645 => "101001101001010001000000",
7646 => "101011000111011101000000",
7647 => "101110000100110100100010",
7648 => "110011000011000100001100",
7649 => "111001101101111101110110",
7650 => "000000101110101101001000",
7651 => "000110010001010100101011",
7652 => "001000111010110111001001",
7653 => "001001001000011111100000",
7654 => "001001011110110011000001",
7655 => "001010101101111000010100",
7656 => "001011000100111101010111",
7657 => "001010100110010101011110",
7658 => "001010111101000000111000",
7659 => "001101001101010111100100",
7660 => "010001101011100011101100",
7661 => "010110011011110011011000",
7662 => "011001001100110101110011",
7663 => "011010111001110000001111",
7664 => "011100001100100011011011",
7665 => "011100001100001001011101",
7666 => "011011100101000110000010",
7667 => "011001001111010111101010",
7668 => "010010010000010100011100",
7669 => "001001101101010010100111",
7670 => "000101010101100011110110",
7671 => "000011110110010110100000",
7672 => "111111110011111111101111",
7673 => "111000000011111100011001",
7674 => "110000111001110100101010",
7675 => "101110100010001101000000",
7676 => "110000010010111010100000",
7677 => "110100000010000111110100",
7678 => "111001010010101110010111",
7679 => "111101101100101010110111",
7680 => "111110001111101000001111",
7681 => "111100000000100100010111",
7682 => "111001011110101111111111",
7683 => "110111101111111101101010",
7684 => "110110100110100001110100",
7685 => "110011100001111100110010",
7686 => "101101101010101101010100",
7687 => "101001101001111011010010",
7688 => "101011010010101000100110",
7689 => "101111111010001001000100",
7690 => "110011010100000110010000",
7691 => "110101101111101100010110",
7692 => "111010000111001110101001",
7693 => "000001001110010000001010",
7694 => "001000111000011110111011",
7695 => "001101011100010110110010",
7696 => "001100100111001100011100",
7697 => "001001001011111100010010",
7698 => "001000001100000010111100",
7699 => "001010000111000111110101",
7700 => "001011111001101001001110",
7701 => "001011011111000101101110",
7702 => "001001001111001110101001",
7703 => "000111101100101010000110",
7704 => "000111110010101000101010",
7705 => "000110100101011000111110",
7706 => "000001110111011000011000",
7707 => "111011010101110111101111",
7708 => "110110101101011101101001",
7709 => "110101100110000111110000",
7710 => "110101001100001110101110",
7711 => "110011101011110000100010",
7712 => "110100100010101110001110",
7713 => "111001100111110010111111",
7714 => "111111000001000011100001",
7715 => "000001001110011111011100",
7716 => "000001011111111111000101",
7717 => "000011101111110101110100",
7718 => "001001101000111111111111",
7719 => "001111101111101000010010",
7720 => "010001011110000101100010",
7721 => "001110101111111100100100",
7722 => "001011000111111101110001",
7723 => "001000100110010101010101",
7724 => "000110010110001111101010",
7725 => "000011100111001001100100",
7726 => "000000000101111100000000",
7727 => "111011001100100000101101",
7728 => "110101110001111110101010",
7729 => "110001011010100111001010",
7730 => "101110011010101100100100",
7731 => "101101010111000010000010",
7732 => "101110111011111111101100",
7733 => "110010011100001111100100",
7734 => "110111000100010100111110",
7735 => "111100001111011101011001",
7736 => "000000111111100101001101",
7737 => "000100110110001000101100",
7738 => "000111101101101101011001",
7739 => "001001010000101100010001",
7740 => "001001000111101111010101",
7741 => "001000000001101011101111",
7742 => "001000100011111100111000",
7743 => "001011011110111111110001",
7744 => "001101000011101001001100",
7745 => "001011011000010111100000",
7746 => "001010011110011100010101",
7747 => "001100111001011100110110",
7748 => "001111000010010100000010",
7749 => "001101100010011010011110",
7750 => "001001110110011101011101",
7751 => "000110001011111011011100",
7752 => "000010100101011011001110",
7753 => "111110100010100001100100",
7754 => "111001111010000110101111",
7755 => "110101010010110001100001",
7756 => "110010001001011010010110",
7757 => "110001010101010110100010",
7758 => "110011001010010111100010",
7759 => "110111100101011101001000",
7760 => "111100101111001010111110",
7761 => "000000010101001101010000",
7762 => "000010001100011011100111",
7763 => "000011001000001000100110",
7764 => "000010110011110011010011",
7765 => "111111111010011010101010",
7766 => "111010101110010100110101",
7767 => "110110000010011110010010",
7768 => "110010111001111001000110",
7769 => "101111101111000001101110",
7770 => "101101011011101011000000",
7771 => "101110101111111111100100",
7772 => "110010111110111001110100",
7773 => "110110111000000101001110",
7774 => "111000111101000000100010",
7775 => "111010001111110011100000",
7776 => "111100000100011010011001",
7777 => "111101111001110101010000",
7778 => "111101111101100111000101",
7779 => "111100000011001000001001",
7780 => "111010001011110011011101",
7781 => "111001100111111011100010",
7782 => "111001110100000000101101",
7783 => "111010111101111010110110",
7784 => "111110001001000001111011",
7785 => "000010101100011111010111",
7786 => "000110111010011100110011",
7787 => "001010011101000000001111",
7788 => "001110001100101001100100",
7789 => "010001111111111111000100",
7790 => "010100100000110001011010",
7791 => "010101111000101110001000",
7792 => "010111010011100100001110",
7793 => "011000000100100011101101",
7794 => "010111100011000101101100",
7795 => "010111000101000001010000",
7796 => "010111000111001110011010",
7797 => "010110111001110010010110",
7798 => "010110010001110000111100",
7799 => "010100100001001001011100",
7800 => "010000111001111101000010",
7801 => "001101001101000110001000",
7802 => "001011101011001110101000",
7803 => "001011000111110101010111",
7804 => "001000100011101110100101",
7805 => "000011111010111110000100",
7806 => "111111101010100101100110",
7807 => "111101001110011101000111",
7808 => "111011110001010100011010",
7809 => "111000011110100010111011",
7810 => "110001111000011001011110",
7811 => "101011001110100100100110",
7812 => "100111110110111000111001",
7813 => "100110110000001001001101",
7814 => "100110010101101010100011",
7815 => "100110010100111011111001",
7816 => "100101101100110010000011",
7817 => "100100011111110011001011",
7818 => "100100010110000101010001",
7819 => "100100111101111001110011",
7820 => "100100111001000101111111",
7821 => "100100110111001101010101",
7822 => "100101101110100010111101",
7823 => "100110001000110001010001",
7824 => "100110101011110111000111",
7825 => "101010100101011010111100",
7826 => "110001010011010111101000",
7827 => "110110110010111101100110",
7828 => "111010000101100101000001",
7829 => "111101011001111101100011",
7830 => "000001111100001111001001",
7831 => "000110011100011010000100",
7832 => "001000011011011111100110",
7833 => "000111000010011001111100",
7834 => "000100111100100100000011",
7835 => "000101101110010110010001",
7836 => "001001010001010000101011",
7837 => "001011110111110000101100",
7838 => "001011010110110010100001",
7839 => "001001100101111111000110",
7840 => "001000111001100010101010",
7841 => "001000110101001101111000",
7842 => "000111111010111110110010",
7843 => "000110011011100100000010",
7844 => "000101101110011010011101",
7845 => "000110111110101110011001",
7846 => "001011000000001001100110",
7847 => "010000000111110101000110",
7848 => "010011010101000001110000",
7849 => "010101101011000100110110",
7850 => "011001011110000101111000",
7851 => "011100111000011111110001",
7852 => "011110000110010101000111",
7853 => "011101100100110100111010",
7854 => "011011101100000110111111",
7855 => "011010001010010001001000",
7856 => "011001110110100110011101",
7857 => "010111110100101001001110",
7858 => "010010011101010110100110",
7859 => "001100000001000100100000",
7860 => "000111000100000000000000",
7861 => "000011111100001100111110",
7862 => "000000011100101100100101",
7863 => "111011010010000110110110",
7864 => "110101110011001100011010",
7865 => "110000110001000011010100",
7866 => "101100111100100011100110",
7867 => "101100001101100000101010",
7868 => "101110001110110010010000",
7869 => "110001010110111010010010",
7870 => "110101101000111001110101",
7871 => "111011100000000100111111",
7872 => "000010001100011101111010",
7873 => "001000011001111100001110",
7874 => "001101110011011001001000",
7875 => "010001111101101011000010",
7876 => "010010010001101001010100",
7877 => "001110010110010101100100",
7878 => "001010010110110011000000",
7879 => "000111111100010000101010",
7880 => "000100001111111101110010",
7881 => "111101111010101110100111",
7882 => "110111001110010001110111",
7883 => "110011011010011101111000",
7884 => "110010110000101010100100",
7885 => "110010011011111101010100",
7886 => "110001010110000011110010",
7887 => "110000101010000110111100",
7888 => "110000110111011100001110",
7889 => "110001101101001111010000",
7890 => "110001111110000111000110",
7891 => "110000101110101101110010",
7892 => "101111011000100101011000",
7893 => "101110110001011010001100",
7894 => "101110111000111111001000",
7895 => "110001110001111001110010",
7896 => "110111000000111111101010",
7897 => "111010001110101001100111",
7898 => "111011001101000100000010",
7899 => "111101010011100010000011",
7900 => "111111100100000000111101",
7901 => "111110110111001100001111",
7902 => "111011101101010001101111",
7903 => "111000110100001000001001",
7904 => "110111001110010111011001",
7905 => "110101001010110111110011",
7906 => "110001101110110110011110",
7907 => "101111011010100001000000",
7908 => "101111001100000100110010",
7909 => "101110101010111111000100",
7910 => "101101100100000110001010",
7911 => "101110001100010101000000",
7912 => "110001111111111011011010",
7913 => "111000100100101100010011",
7914 => "111111110101011011001000",
7915 => "000110000101001010110000",
7916 => "001011000010010001110101",
7917 => "001110010011000110101110",
7918 => "001111111010111100010100",
7919 => "010000011000010011010000",
7920 => "001111110101000101010010",
7921 => "001111001001111100101000",
7922 => "001110010100110101010010",
7923 => "001101000010000101110100",
7924 => "001101010011110000111010",
7925 => "001110111010111100111110",
7926 => "010000000000101111111000",
7927 => "010011000011010100001000",
7928 => "011000001010111110000101",
7929 => "011010001110110110000111",
7930 => "011000110101000011000101",
7931 => "010111101100110010011110",
7932 => "010111011110110100000100",
7933 => "010111000101000111000010",
7934 => "010110011110001111111000",
7935 => "010110100001001101001110",
7936 => "010110001110000101010110",
7937 => "010010111011010100000000",
7938 => "001110101001000111001110",
7939 => "001100111000001110100110",
7940 => "001010110011101100001101",
7941 => "000110011010010010010010",
7942 => "000011011001111111010011",
7943 => "000010101000111111011110",
7944 => "000001110101101001000111",
7945 => "000001000011101110100011",
7946 => "111110001011011110000111",
7947 => "110100110100111001010011",
7948 => "101000011111101001000010",
7949 => "100001111111011001110000",
7950 => "100001101111011100100010",
7951 => "100001110101110101100000",
7952 => "100001001011101100011110",
7953 => "100001011011110110101111",
7954 => "100010001110000111001100",
7955 => "100011000000011011101011",
7956 => "100011010111010101010110",
7957 => "100011011010000110001111",
7958 => "100100000011101001111101",
7959 => "100100101011111000101011",
7960 => "100101100111100011101111",
7961 => "101001010001110001111100",
7962 => "101110110101000100100000",
7963 => "110010110111100010000100",
7964 => "110100001000000001000111",
7965 => "110011101111110111010010",
7966 => "110100101100010100011011",
7967 => "111000011101101110101000",
7968 => "111100000011111111111100",
7969 => "111100100101100001011000",
7970 => "111010101111110010011101",
7971 => "111000010110111000001100",
7972 => "110110110111010000010111",
7973 => "110110110100001100110000",
7974 => "110111011000010100011010",
7975 => "110111101100110000000010",
7976 => "110111111100101001011010",
7977 => "111001010010111000111101",
7978 => "111100101110110000110011",
7979 => "000000111101111001101011",
7980 => "000011010010011100010100",
7981 => "000011100110000001010010",
7982 => "000101010110101111011010",
7983 => "001010100001001000111000",
7984 => "010000010110001011110110",
7985 => "010100101110100100100010",
7986 => "011001001100010100110011",
7987 => "011101011000100001111110",
7988 => "011110110111011111010111",
7989 => "011110101111101001100111",
7990 => "011110110010110101000010",
7991 => "011101011110001000010101",
7992 => "011010001111000110111111",
7993 => "010110111000011000000100",
7994 => "010011100100100011000010",
7995 => "001111001000100010111000",
7996 => "001001101100101001001100",
7997 => "000101001111100100010010",
7998 => "000100000001011111101001",
7999 => "000101110000010100001100",
8000 => "000111111111101000100100",
8001 => "001001001110001100010001",
8002 => "001001101101101000111110",
8003 => "001010011101100011101111",
8004 => "001011001011101101111010",
8005 => "001010101000110000101000",
8006 => "001010000000100011001011",
8007 => "001010111001001001000010",
8008 => "001011111110001001001000",
8009 => "001100101101000101001110",
8010 => "001101101001000101100010",
8011 => "001101011011110011111110",
8012 => "001011110110110100010100",
8013 => "001001110101000011100110",
8014 => "000110110000110110001010",
8015 => "000011010110000011111000",
8016 => "000000110010000000110011",
8017 => "111101100110000000110111",
8018 => "111000010010100010001111",
8019 => "110001101100001110100000",
8020 => "101100110101100110010000",
8021 => "101100010110101000111000",
8022 => "101101101011100001111100",
8023 => "101100111110010101011010",
8024 => "101100000111100000001100",
8025 => "101110010010100111111010",
8026 => "110010010111101110100000",
8027 => "110101111110010010010010",
8028 => "111000100011000111011101",
8029 => "111001111111100111100001",
8030 => "111001110000000010110011",
8031 => "111000110010101100101010",
8032 => "111000100001010110111111",
8033 => "110111000100100001000100",
8034 => "110010110111110101001000",
8035 => "101110110001011110010110",
8036 => "101100110001101001110010",
8037 => "101010111100111110100000",
8038 => "101000000000100101011100",
8039 => "100101100110010110011101",
8040 => "100101011100111111110011",
8041 => "100110101010000110001101",
8042 => "100111101101110101111111",
8043 => "101001000011111110110100",
8044 => "101010111100011101001110",
8045 => "101101000001101100111010",
8046 => "101111110000101110101010",
8047 => "110010111000101010110000",
8048 => "110110001010000110011100",
8049 => "111010001101010010011000",
8050 => "111110010100010100000010",
8051 => "000010001000111100000000",
8052 => "000111000100010111101000",
8053 => "001100011111001111100110",
8054 => "001111110110010110010110",
8055 => "010000111000011011101010",
8056 => "010001110110011110010100",
8057 => "010011101110011011111010",
8058 => "010100111111110100001010",
8059 => "010101011111011110110100",
8060 => "010110100101100101100110",
8061 => "010111101011001001000010",
8062 => "011000001111001010100010",
8063 => "011001011100110110101111",
8064 => "011010101111000000100010",
8065 => "011010100111111101000111",
8066 => "011001101100000111010111",
8067 => "011000111100100001010100",
8068 => "011000010100000111100101",
8069 => "010111101100000110010100",
8070 => "010111101011010101101000",
8071 => "011000000111100100010011",
8072 => "010111110100010011010100",
8073 => "010110111111101010110100",
8074 => "010110011111100110001000",
8075 => "010110000110110111011000",
8076 => "010101111001010011101010",
8077 => "010100100101100011011000",
8078 => "001111100111100000110010",
8079 => "000111100101100101011011",
8080 => "111111001000100100110000",
8081 => "111000001001111101011101",
8082 => "110011000110110111110100",
8083 => "101101000110000011101100",
8084 => "100101010101101110010101",
8085 => "100001000101011010001011",
8086 => "100001011001101011011110",
8087 => "100001100010101110011111",
8088 => "100001001010000001100011",
8089 => "100010000001001100110111",
8090 => "100010101110111001100100",
8091 => "100011000001000011000111",
8092 => "100011110100100011011111",
8093 => "100100110000111110000111",
8094 => "100110110111010100011101",
8095 => "101011101111000000001110",
8096 => "110001100100010001100000",
8097 => "110101011100011100001011",
8098 => "110111111100011000011100",
8099 => "111011110110110111111111",
8100 => "000000111110011110100111",
8101 => "000010111001111100111000",
8102 => "111111100010101100011000",
8103 => "111011000010010010100001",
8104 => "111000010110011011010000",
8105 => "110100101011110011111000",
8106 => "101111000100000101110100",
8107 => "101010101110010011111000",
8108 => "101000101100000001001010",
8109 => "101000000110111100000010",
8110 => "101010000111000111101110",
8111 => "110000000001010111110000",
8112 => "111000000110101100100001",
8113 => "111101110111010110101000",
8114 => "000000000110000101100101",
8115 => "000011100001000111001101",
8116 => "001001011001001001000111",
8117 => "001100010001100101110100",
8118 => "001011000000000111011010",
8119 => "001010110100010100000101",
8120 => "001101111101110110001100",
8121 => "010001110101011001101110",
8122 => "010100001101100111011100",
8123 => "010101101010010000100100",
8124 => "010111001001110000111110",
8125 => "010111010001101101010010",
8126 => "010100011011111101000000",
8127 => "001111100011100001110000",
8128 => "001010000011010010101100",
8129 => "000101010101011100001101",
8130 => "000011000110000110001101",
8131 => "000010001000111110101011",
8132 => "000000001111001100000110",
8133 => "111110011110001000100110",
8134 => "111101110100111111110110",
8135 => "111101111101011110101001",
8136 => "000000010001111010000001",
8137 => "000011110010111111011111",
8138 => "000101000100011011000011",
8139 => "000101110100011010000100",
8140 => "001000110010111100110100",
8141 => "001011001001000110110000",
8142 => "001010101110100000001110",
8143 => "001001100010101110011101",
8144 => "001001011000101110010110",
8145 => "001010100001011011111000",
8146 => "001011110110101000000111",
8147 => "001100001011100111110010",
8148 => "001100000011110010001100",
8149 => "001100001011100110011000",
8150 => "001011110110111111001100",
8151 => "001001101101101110001101",
8152 => "000110000110011110101110",
8153 => "000100010001010100011111",
8154 => "000100111110010101101110",
8155 => "000100100110000111000011",
8156 => "000010010100110110101110",
8157 => "000001000001000101101010",
8158 => "000001101100110011001111",
8159 => "000011000011011101000101",
8160 => "000011011001011110100000",
8161 => "000010101101111110110110",
8162 => "000010011001111100001011",
8163 => "000010010111010101011110",
8164 => "000010000010011101110100",
8165 => "000001011101100000110011",
8166 => "111111101001100110001011",
8167 => "111100100001010101100101",
8168 => "111001101010010000010101",
8169 => "110111111010100101001000",
8170 => "110110111000011010110000",
8171 => "110100101010010100010010",
8172 => "110000010110000101011000",
8173 => "101100111001100100000000",
8174 => "101100001101101101001100",
8175 => "101011111010010110001110",
8176 => "101010010010111111111100",
8177 => "101000110011100011101110",
8178 => "101001101011000011101100",
8179 => "101101000101101011111110",
8180 => "110000111011100001000110",
8181 => "110100010110000111010111",
8182 => "111000011001101110111000",
8183 => "111100111010101001000001",
8184 => "000000011111011001011011",
8185 => "000010010110111011010001",
8186 => "000010100011010011011011",
8187 => "000001010000100111100100",
8188 => "111110111001001010101011",
8189 => "111101000000101011110011",
8190 => "111100110110010001000010",
8191 => "111101101010011101111100",
8192 => "111111001110100100110100",
8193 => "000010011000010110110111",
8194 => "000110100010100100110001",
8195 => "001010101011010011010110",
8196 => "001110101010000100101000",
8197 => "010001111011010010010100",
8198 => "010011101100010110000110",
8199 => "010100001100011010101100",
8200 => "010100011000010110101010",
8201 => "010101001100011011010110",
8202 => "010110111100000010110100",
8203 => "011000011010110011001100",
8204 => "011000011011101101110001",
8205 => "011000000001011000111101",
8206 => "011000000011001101111001",
8207 => "010111011110101110110110",
8208 => "010110011001110110101100",
8209 => "010101110010111001110110",
8210 => "010101101010101101000100",
8211 => "010101010001011010111110",
8212 => "010001101100000011111000",
8213 => "001001100101110000110100",
8214 => "000000100010101100100000",
8215 => "110110111011010000110100",
8216 => "101011000100001100001110",
8217 => "100010100011001111011101",
8218 => "100001010100100101111111",
8219 => "100010001000011100010001",
8220 => "100001011111111110100011",
8221 => "100001010101011110111111",
8222 => "100010010011000101111111",
8223 => "100011001000001001100001",
8224 => "100100000001101100000111",
8225 => "100111000111110000111100",
8226 => "101011011011100011101010",
8227 => "101100111101010111000010",
8228 => "101100111101001101110000",
8229 => "101110101111011110010000",
8230 => "110000001010000001010100",
8231 => "110000010111000000011010",
8232 => "110010111001011000110110",
8233 => "111000000000111100101000",
8234 => "111100001001111100110011",
8235 => "111101010001011011101110",
8236 => "111100111100011010101001",
8237 => "111101010101111001011100",
8238 => "111100101001010011001011",
8239 => "111000100110000001010011",
8240 => "110011110001000111110110",
8241 => "110001011101111110000010",
8242 => "110001111010101100010100",
8243 => "110011111111100001010000",
8244 => "110110001100111100110111",
8245 => "110111101111001101101111",
8246 => "111001100011000100010100",
8247 => "111101000101100100011110",
8248 => "000010111110000111000011",
8249 => "001010001011101111111100",
8250 => "010000000011110001000110",
8251 => "010011000101011010101110",
8252 => "010101100111000110001100",
8253 => "011010001111111010111011",
8254 => "011110000111001100010011",
8255 => "011100011000000001111111",
8256 => "010110010000100100101110",
8257 => "010000110100001101001010",
8258 => "001101010010000001010110",
8259 => "001001001101001010101000",
8260 => "000100000100011010010011",
8261 => "000000011100000001110010",
8262 => "111111010101110111110010",
8263 => "111110110011100110111101",
8264 => "111110000101111000011011",
8265 => "111110011001100100111100",
8266 => "111111110110010001101000",
8267 => "000001110000100000100110",
8268 => "000011011111101110110000",
8269 => "000011110110001100110100",
8270 => "000010001111011011000001",
8271 => "111111110111111010100111",
8272 => "111110010111110101001110",
8273 => "111110000011000011110001",
8274 => "111101111001000001011001",
8275 => "111101010100110010010001",
8276 => "111100110001101001001001",
8277 => "111100010010101011110011",
8278 => "111011011100010000100000",
8279 => "111010001011101101101011",
8280 => "111000100011111011010011",
8281 => "110110110110101010011000",
8282 => "110101111101010110010111",
8283 => "110101111000110010111010",
8284 => "110101100011001100110100",
8285 => "110101001011010111001000",
8286 => "110101101111101100100100",
8287 => "110110010111111100010000",
8288 => "110101111000110111010111",
8289 => "110101010010100000111100",
8290 => "110110011000110010110100",
8291 => "111001010111110110011110",
8292 => "111100100000111101010111",
8293 => "111110011001100111110001",
8294 => "111111100011111010011101",
8295 => "000001000010101001010011",
8296 => "000011001100000001101010",
8297 => "000101010110001110001011",
8298 => "000101111101000101010000",
8299 => "000101001101011100000110",
8300 => "000101100001101101100000",
8301 => "000111100011111101100000",
8302 => "001001101011001000110000",
8303 => "001010100111000101110110",
8304 => "001010000001100000000110",
8305 => "001000010001110110101000",
8306 => "000110010111001001011100",
8307 => "000101000100001000000100",
8308 => "000100001100111011110110",
8309 => "000010111001100001101011",
8310 => "000001011010010011110111",
8311 => "000001000101010000110111",
8312 => "000001110110111100011010",
8313 => "000010001101101001110100",
8314 => "000001010000111110001101",
8315 => "000000000010010101001001",
8316 => "000000001100100100001110",
8317 => "000001010110001111100001",
8318 => "000010000101010110000011",
8319 => "000010010011111101001111",
8320 => "000010011010011000011011",
8321 => "000011001010000100000011",
8322 => "000100100000110000011101",
8323 => "000100001100010000000010",
8324 => "000010001101000010111011",
8325 => "000001100110100000100100",
8326 => "000011001010111010110110",
8327 => "000110000001110011111111",
8328 => "001001000111100100011000",
8329 => "001010110000001111101101",
8330 => "001011011011011101110100",
8331 => "001100101111101000110100",
8332 => "001110111010111010111010",
8333 => "010010100000000100001100",
8334 => "010110101010001111100110",
8335 => "011000111001000101011011",
8336 => "011001010001100011011110",
8337 => "011001001100110000100011",
8338 => "011000101100000010001101",
8339 => "010111101000001011101010",
8340 => "010110011110101011011000",
8341 => "010101110001000011101000",
8342 => "010100000010101100001110",
8343 => "001111001110110100010000",
8344 => "001001010000010011110100",
8345 => "000100001111010000110101",
8346 => "111110010111100000101101",
8347 => "110110111100110011011011",
8348 => "101111011111111001101000",
8349 => "101001000101111011110100",
8350 => "100101010111100100101111",
8351 => "100101000011101010100000",
8352 => "100110101011000101001010",
8353 => "101000100011101100111010",
8354 => "101001111101010100010110",
8355 => "101011110001111100101000",
8356 => "101111010001111011001100",
8357 => "110011101110100001011010",
8358 => "110111000011010001101110",
8359 => "110110100110010100001111",
8360 => "110010100111111011111100",
8361 => "110000011001001011000110",
8362 => "110001101111101110001100",
8363 => "110010100001011110000110",
8364 => "110001101111111111100110",
8365 => "110001100100111100000000",
8366 => "110001011001111001000110",
8367 => "101111100011110101111100",
8368 => "101011110110111111010010",
8369 => "101000000010101001100100",
8370 => "100110011100100100111111",
8371 => "100110111001101111110010",
8372 => "101000010010010111101010",
8373 => "101011100010111110010010",
8374 => "110001100001001000001010",
8375 => "111000101111111111101101",
8376 => "111111000101010100111000",
8377 => "000100000010011001101100",
8378 => "001000011111001100100010",
8379 => "001100100101101101111010",
8380 => "010000001001100001100110",
8381 => "010011000010001000100000",
8382 => "010100010010011101101110",
8383 => "010011101010101011000100",
8384 => "010010101100110011001100",
8385 => "010011100000010100110010",
8386 => "010110111110001110100010",
8387 => "011010010111010011100010",
8388 => "011010011001100001000001",
8389 => "011001000011101101010101",
8390 => "011001011000001111110010",
8391 => "011001000111011100110101",
8392 => "010100011001111011010100",
8393 => "001011011110010100001100",
8394 => "000010111100100011010010",
8395 => "111110110101011000011100",
8396 => "111101111111011010111100",
8397 => "111110010101100000110100",
8398 => "000000111110111000001100",
8399 => "000101100010111100101110",
8400 => "001001001000101010101100",
8401 => "001011001101000000001101",
8402 => "001100111011001101111000",
8403 => "001110110011110000110100",
8404 => "010001010101111000010010",
8405 => "010011101101000110110110",
8406 => "010011010100001000010000",
8407 => "001111011011101110111100",
8408 => "001001110011010010000100",
8409 => "000011100110010110101100",
8410 => "111101011011111000110010",
8411 => "111000001101010001001110",
8412 => "110011101110000001101100",
8413 => "101111100000000010101010",
8414 => "101100001010011101111100",
8415 => "101001011010100010010100",
8416 => "100110000100001111101010",
8417 => "100010101110100010111011",
8418 => "100001000000110101101101",
8419 => "100001001110000110000001",
8420 => "100010100101111010001001",
8421 => "100100100111010000101011",
8422 => "100111100001110000100101",
8423 => "101011010001111000100000",
8424 => "101110101101100110101100",
8425 => "110001000111000110001000",
8426 => "110010101111110100100100",
8427 => "110011111001111010101110",
8428 => "110101100110110011001000",
8429 => "111000101101011100000111",
8430 => "111011010000111111111000",
8431 => "111011011110100000110010",
8432 => "111011110010010110111000",
8433 => "111110100111011001010100",
8434 => "000001110001101001101101",
8435 => "000010100100100010010100",
8436 => "000001110111001101011011",
8437 => "000001010100000100000000",
8438 => "000000011000001111011000",
8439 => "111101111001110100010000",
8440 => "111010101010011011011010",
8441 => "111000000111001100011101",
8442 => "110110000101011011001010",
8443 => "110100101110011010001110",
8444 => "110101110010010001111011",
8445 => "111001011000000101110101",
8446 => "111110000000110101000011",
8447 => "000011011101010011011000",
8448 => "001000111000101101110110",
8449 => "001100001001001010100000",
8450 => "001101001000111101011000",
8451 => "001101001001001101110010",
8452 => "001100010100010111010010",
8453 => "001011011100010011110101",
8454 => "001011110111001101110110",
8455 => "001100111010011100101110",
8456 => "001101101000001101110110",
8457 => "001111001111001000010100",
8458 => "010010101010100000011000",
8459 => "010110010000111000000010",
8460 => "010111111001011111101110",
8461 => "010111011010100100010110",
8462 => "010110100010101111100000",
8463 => "010110101010011100010010",
8464 => "010110111101011101000100",
8465 => "010101110110110000110010",
8466 => "010011011000011110110010",
8467 => "010000111110001111100000",
8468 => "010000000011110011001000",
8469 => "010000110110001101111010",
8470 => "010010001101000110001010",
8471 => "010011011100101101000100",
8472 => "010100110001010101111110",
8473 => "010101110000010011110000",
8474 => "010101001111101010110010",
8475 => "010010000101101100110110",
8476 => "001011110101010010100110",
8477 => "000011011111010111001011",
8478 => "111010111101101111011100",
8479 => "110011110010010111011100",
8480 => "101110010110001000010100",
8481 => "101010001001000110010110",
8482 => "100111100001011101110101",
8483 => "100111101010011100100111",
8484 => "101010010101100001010010",
8485 => "101110000111001001001110",
8486 => "110010010101011110011110",
8487 => "110111001111101110110000",
8488 => "111100100010001011110011",
8489 => "000000101001110100100011",
8490 => "000001111110111001110010",
8491 => "111111110110010011011011",
8492 => "111011001011100001111101",
8493 => "110110111010100000000110",
8494 => "110100001101111001001001",
8495 => "110000001000111000111010",
8496 => "101001100011001010001100",
8497 => "100100000100110010011101",
8498 => "100010100101010010111011",
8499 => "100011110011101010000110",
8500 => "100100101111101101011101",
8501 => "100100101110000100011110",
8502 => "100101001010100101000001",
8503 => "100110000001000110110111",
8504 => "100111000011000011010000",
8505 => "101000010100110110000100",
8506 => "101000001111001001100100",
8507 => "101001000010100001000110",
8508 => "101110111101010001011000",
8509 => "110101111011010100011111",
8510 => "111010010100010110000110",
8511 => "000001001001111110001100",
8512 => "001010101010001100010110",
8513 => "010001000111010101111000",
8514 => "010101000001111011110110",
8515 => "011001000011111011110101",
8516 => "011100001110010000110001",
8517 => "011110000101011001001001",
8518 => "011110100001011110110111",
8519 => "011011110110010010110011",
8520 => "010101110011110010100000",
8521 => "001111001111101110100000",
8522 => "001010111010011110111001",
8523 => "001000001001000110011010",
8524 => "000101011101101100100001",
8525 => "000011110010101000101100",
8526 => "000100010000110001000101",
8527 => "000111001101110011100001",
8528 => "001011111100101001110000",
8529 => "001111001101100001011100",
8530 => "001110111010001010101110",
8531 => "001101100011000101011000",
8532 => "001101111101101011011000",
8533 => "001111010110011110001110",
8534 => "001111101011101101101000",
8535 => "001111101100110110101000",
8536 => "010001010011010010001010",
8537 => "010011000101010010100100",
8538 => "010010110000000010011010",
8539 => "010001001010101100100110",
8540 => "001111110000000101110110",
8541 => "001110101011111001111100",
8542 => "001101111001110100100000",
8543 => "001011110100011111100001",
8544 => "000110001010010101101110",
8545 => "111101110001010110110011",
8546 => "110101111001100011101011",
8547 => "101111001001100010000000",
8548 => "100111111101100110011101",
8549 => "100010001111011000100101",
8550 => "100000110010001010010011",
8551 => "100001010111011001111001",
8552 => "100001010011110010000101",
8553 => "100001010100001000000001",
8554 => "100001101011100110100011",
8555 => "100011000010000101001001",
8556 => "100111001011111110010011",
8557 => "101101001111011010001100",
8558 => "110010110001101100100100",
8559 => "110111001000110111000000",
8560 => "111010011100110001100111",
8561 => "111100011100010000111111",
8562 => "111100001100000111010111",
8563 => "111001100101000110101010",
8564 => "110110101101100100010101",
8565 => "110101000111110111010001",
8566 => "110100100001110111111111",
8567 => "110100010100001000001000",
8568 => "110011001110111010111110",
8569 => "110001011001010000001000",
8570 => "110001010111110010011110",
8571 => "110011000111001110100010",
8572 => "110011110010110011000100",
8573 => "110011110010101010110100",
8574 => "110101011011111010111100",
8575 => "111000010110010100111101",
8576 => "111011001011011001001111",
8577 => "111101111100111111110000",
8578 => "000000011011111111011101",
8579 => "000001101000110000000010",
8580 => "000001101101111001011011",
8581 => "000010001010000110100111",
8582 => "000011011010101010010111",
8583 => "000100001011111110111000",
8584 => "000011111010001010101111",
8585 => "000011110110011000110100",
8586 => "000100100010010000100100",
8587 => "000100111110111111000101",
8588 => "000101001000000010011001",
8589 => "000110000001000111010010",
8590 => "001000000011101010001000",
8591 => "001010111001011000111110",
8592 => "001101110000100110011000",
8593 => "001111010111001001000000",
8594 => "001111010110001110101000",
8595 => "001111010011111110001010",
8596 => "010000100001101000010010",
8597 => "010001110001001110000110",
8598 => "010001010101101100010110",
8599 => "001111111001100000001000",
8600 => "001111101110100111000110",
8601 => "010001101111011011001010",
8602 => "010100001000001100101100",
8603 => "010100110111100101011000",
8604 => "010100100110000100111000",
8605 => "010101000000011010110100",
8606 => "010110001100011000000100",
8607 => "010110101000100101001010",
8608 => "010100100110000010001110",
8609 => "010000100010010011001010",
8610 => "001100101100011001011100",
8611 => "001001000010110011110000",
8612 => "000100001111111010110001",
8613 => "111111011011111100011000",
8614 => "111100100101110010101111",
8615 => "111100001110011111100100",
8616 => "111101111000010110001001",
8617 => "000000101100001001000100",
8618 => "000011111010110100110000",
8619 => "000110101110111110000011",
8620 => "001000101010100100000110",
8621 => "001010000101111011000100",
8622 => "001010000111111010011000",
8623 => "000111111111111111111101",
8624 => "000110000000011010001101",
8625 => "000101110000100101001110",
8626 => "000110000111101000111110",
8627 => "000101000000001110011000",
8628 => "111111110010111110111100",
8629 => "110111100100110010010010",
8630 => "110000111000000001111000",
8631 => "101011001011001010100000",
8632 => "100100100010111110110101",
8633 => "100000111110011111000011",
8634 => "100001110100001101001010",
8635 => "100010101111101111001111",
8636 => "100010111100110000001101",
8637 => "100011101001010011011111",
8638 => "100011101111011001111001",
8639 => "100100110111111001010111",
8640 => "101001101111000101011000",
8641 => "101111011101010111100100",
8642 => "110011000110101011101010",
8643 => "110111000101011101101001",
8644 => "111100001101110101101110",
8645 => "111111011000100101010000",
8646 => "000000000110011010010000",
8647 => "000000101110110001111010",
8648 => "000011000001010101100111",
8649 => "000111010100100011001000",
8650 => "001011001011101011000101",
8651 => "001011110101010111010001",
8652 => "001010100010000111001101",
8653 => "001001100100010101001110",
8654 => "001000111010000111001101",
8655 => "000111100000110011100000",
8656 => "000011111111111100101010",
8657 => "111110100001110111000001",
8658 => "111010100100001010010000",
8659 => "111011101000011101010010",
8660 => "000001001011000010100001",
8661 => "000110101010101101100001",
8662 => "001001011110100000000101",
8663 => "001100111101001100101110",
8664 => "010011100110101110111110",
8665 => "011001100101010000000101",
8666 => "011011100001000000010111",
8667 => "011011000100101010010011",
8668 => "011010101000011110000001",
8669 => "011010010001011011011001",
8670 => "011000110011101001100011",
8671 => "010101110110000110001000",
8672 => "010010001010010010101100",
8673 => "001101111010000100001100",
8674 => "001000110001111101001000",
8675 => "000011001111101110110001",
8676 => "111110000100100001110011",
8677 => "111010011110101111011011",
8678 => "111001011110110000100110",
8679 => "111001101111001011110010",
8680 => "111001000100100100111001",
8681 => "110111001000001110101110",
8682 => "110100001011101011100010",
8683 => "110000010111100100011100",
8684 => "101100110101000111110010",
8685 => "101010011100010001110010",
8686 => "101000110111001000001110",
8687 => "101000011010110101011100",
8688 => "101001100101000100101000",
8689 => "101011000110010010011010",
8690 => "101100000011011111111010",
8691 => "101101001111111000111100",
8692 => "101111010000000111000100",
8693 => "110001111011010001001000",
8694 => "110101000111000000101100",
8695 => "111000010000001101101111",
8696 => "111010011110110010011100",
8697 => "111011000111110101011111",
8698 => "111010010010101100010111",
8699 => "111000100010011100111011",
8700 => "110101101101011001110010",
8701 => "110010010100011100101000",
8702 => "110000100010101111111100",
8703 => "110000111011101000000100",
8704 => "110001101010100011101010",
8705 => "110010100000000101000000",
8706 => "110101001111000000011110",
8707 => "111010100001101001011110",
8708 => "000001000010101101110100",
8709 => "000110111101100100001100",
8710 => "001011011111001100000011",
8711 => "001110111100111010110000",
8712 => "010001001110001000001010",
8713 => "010001000000011001100000",
8714 => "001101101100001101001110",
8715 => "001000100000100011001100",
8716 => "000011000001000001110100",
8717 => "111110001000001011001110",
8718 => "111011000000101001010110",
8719 => "111010100011101001010110",
8720 => "111100000000000011111101",
8721 => "111110001101111001011000",
8722 => "000001010110101010011000",
8723 => "000100110101110010100010",
8724 => "000110001011101011011111",
8725 => "000100101110101000101001",
8726 => "000010111111110100111111",
8727 => "000010010100010011001000",
8728 => "000010000011100111100011",
8729 => "000010010010101010011010",
8730 => "000010110001001100110111",
8731 => "000010101111111001110000",
8732 => "000010111001101000101011",
8733 => "000011101100010101100011",
8734 => "000100010101100001000000",
8735 => "000100001110010000101110",
8736 => "000011001101100011000100",
8737 => "000010000011000010011111",
8738 => "000001001011010001011101",
8739 => "111110101010001001010100",
8740 => "111001010110100010111111",
8741 => "110011010111001101001010",
8742 => "101110110001111011010100",
8743 => "101100001010011010110100",
8744 => "101011001000100111100010",
8745 => "101010110111110110000000",
8746 => "101100001110001000111110",
8747 => "110000101011100011011110",
8748 => "110111000001111111101100",
8749 => "111101000110010000001010",
8750 => "000010110101011111010100",
8751 => "001000111001010101010000",
8752 => "001110011110111001010100",
8753 => "010010011101000111110000",
8754 => "010101001110111000011010",
8755 => "010111011000101100000000",
8756 => "010111111111100110101010",
8757 => "010110110101100000111110",
8758 => "010101010110000000000110",
8759 => "010100011001100100110010",
8760 => "010011011111010110111010",
8761 => "010001101011000110101100",
8762 => "001111100011010000101100",
8763 => "001110001011010011001110",
8764 => "001010101101001011000110",
8765 => "000010100100001001101001",
8766 => "111010100001011100001101",
8767 => "110111101111011000011010",
8768 => "111000000110100110101001",
8769 => "110111010110101010010010",
8770 => "110011111011100011000010",
8771 => "101111100111100010100110",
8772 => "101110001111100000011110",
8773 => "101111110010100011111010",
8774 => "110000111011001111110100",
8775 => "110010010110101010101000",
8776 => "110110110000000011101110",
8777 => "111100011101100001010111",
8778 => "111111011111001111000011",
8779 => "111111000101011011011010",
8780 => "111110111101011000011110",
8781 => "000001000100111001010110",
8782 => "000001111100011001100100",
8783 => "000000000111110001110011",
8784 => "111110111101001111011111",
8785 => "111111001000010001111100",
8786 => "111110100101010111101010",
8787 => "111101001010001011000111",
8788 => "111011101101100111101100",
8789 => "111011100110001101111111",
8790 => "111110011001101101010110",
8791 => "000011111001011110111011",
8792 => "001001111101001000100111",
8793 => "001101100011010001010000",
8794 => "001101101100000011001010",
8795 => "001101100010111111111100",
8796 => "001111100011011010001100",
8797 => "010001100000011101000110",
8798 => "010000010111101001001100",
8799 => "001100010111111101000000",
8800 => "001001001011110000111011",
8801 => "001001010110011011000001",
8802 => "001010001011111010000010",
8803 => "001000001110000101100100",
8804 => "000100010010011011001100",
8805 => "000000111001110110010110",
8806 => "111110111111101000000111",
8807 => "111101110110000001000011",
8808 => "111100101001000001101001",
8809 => "111011101101001000101011",
8810 => "111010111101000011001100",
8811 => "111001100110011010000111",
8812 => "110111111111111110111110",
8813 => "110110101101110001110101",
8814 => "110101111000000101000100",
8815 => "110110010110000000000101",
8816 => "111000011010100101101100",
8817 => "111010101000111111101000",
8818 => "111011100001000011101111",
8819 => "111011001111001100010110",
8820 => "111010110001001010101011",
8821 => "111001100101000010101101",
8822 => "110110111010101010011100",
8823 => "110011110100110011111110",
8824 => "110000110110010001011110",
8825 => "101101110001000100111100",
8826 => "101011101100100011010100",
8827 => "101010110100011011001000",
8828 => "101001111001101110001000",
8829 => "101001110111111110000100",
8830 => "101100101010010000011000",
8831 => "110001100100010110100010",
8832 => "110110011000111001000110",
8833 => "111010010001011101000100",
8834 => "111101011101101010100010",
8835 => "111111011101010111011110",
8836 => "111111110001111011111000",
8837 => "111111011100100110011111",
8838 => "111111110100001001100110",
8839 => "000001101011111100010100",
8840 => "000101001111110110011010",
8841 => "001001100001000100010010",
8842 => "001101100011111001100110",
8843 => "010001100001011110011100",
8844 => "010101011100001010110110",
8845 => "011000110010010100100001",
8846 => "011010101110011001011101",
8847 => "011010101100100101010101",
8848 => "011001011101011011100001",
8849 => "010111111100000010100100",
8850 => "010101101001000100110100",
8851 => "010001110111001000011010",
8852 => "001101001001010110111010",
8853 => "001000110111111001000111",
8854 => "000110001011111010110011",
8855 => "000101101100111001111010",
8856 => "000111001010000001001010",
8857 => "001001000001111000011100",
8858 => "001010011001100011110110",
8859 => "001100000110000111100000",
8860 => "001110011000011101011100",
8861 => "010000000100100000100110",
8862 => "010000000001000001010000",
8863 => "001110100001000101100100",
8864 => "001101101100001000011010",
8865 => "001110000000010010101010",
8866 => "001100110100100111010100",
8867 => "001001010110010011000011",
8868 => "000100111101110010001011",
8869 => "111111100010110011001011",
8870 => "111000101101011001100011",
8871 => "110000011100010111100110",
8872 => "100111011110000011011000",
8873 => "100001100010011110111111",
8874 => "100000101110110111100000",
8875 => "100001101111100000010000",
8876 => "100010000011010101101000",
8877 => "100010010011101110000100",
8878 => "100010101010000010101111",
8879 => "100011010101010001101001",
8880 => "100101111000100000000111",
8881 => "101010110110010110000100",
8882 => "110000110001111110100000",
8883 => "110110101111101011111100",
8884 => "111101000001110100110001",
8885 => "000010010000010011100111",
8886 => "000100110011010000101111",
8887 => "000110001111010000010010",
8888 => "000111111000111111011001",
8889 => "001000111001100010110110",
8890 => "001001110000110101000001",
8891 => "001011000101010011011010",
8892 => "001011001100011110010110",
8893 => "001000110011000000000001",
8894 => "000100011001011011110101",
8895 => "111111001111110001000001",
8896 => "111010100110011010111011",
8897 => "110111101111110000001000",
8898 => "110111101011100000101100",
8899 => "111001011100000011111001",
8900 => "111011000100101000010100",
8901 => "111100000111101110001001",
8902 => "111100110001000001110001",
8903 => "111101111100111110101110",
8904 => "000000110000010110010010",
8905 => "000010111110101010001100",
8906 => "000010100010001010100100",
8907 => "000001000100010000111110",
8908 => "111111100100001001110010",
8909 => "111110011001101011101111",
8910 => "111111100110100111010101",
8911 => "000011000111100101100011",
8912 => "000111001100100011011010",
8913 => "001011010010001000011011",
8914 => "001110011111001111101010",
8915 => "001111101100001101000100",
8916 => "001110110011000110101010",
8917 => "001101000100000100101110",
8918 => "001100100100010011111010",
8919 => "001100110001110110100010",
8920 => "001100000000000010100110",
8921 => "001011111001110100100011",
8922 => "001101011110000011001010",
8923 => "001110011011010100100000",
8924 => "001101110011110000100000",
8925 => "001100011001011011110100",
8926 => "001011100011110010000110",
8927 => "001100111000110011001000",
8928 => "001111110000100010111010",
8929 => "010010010000010011000110",
8930 => "010010110000001100110110",
8931 => "001111111111001101100100",
8932 => "001011110101001111100000",
8933 => "001001010100001010010101",
8934 => "000111101101100111101101",
8935 => "000101010011010101101010",
8936 => "000010001100110111110100",
8937 => "111111100000110110011110",
8938 => "111110101110101101101010",
8939 => "111110101011001101110111",
8940 => "111100011010101111011010",
8941 => "111000101010000010101011",
8942 => "110101110111101101001010",
8943 => "110100110110010101000000",
8944 => "110101100000111010110000",
8945 => "110110010010101000111000",
8946 => "110101110000010010110110",
8947 => "110101000010000110010111",
8948 => "110100100010110111110110",
8949 => "110011000011010011100110",
8950 => "110000110001000010110110",
8951 => "101111001101000001100010",
8952 => "101111010110101010100010",
8953 => "110000011101000111111110",
8954 => "110000100010100110011000",
8955 => "101111001000001111011110",
8956 => "101101000001001101010010",
8957 => "101010100111000011001100",
8958 => "101000011101011101001110",
8959 => "100110110110110100111110",
8960 => "100101101011011111011111",
8961 => "100101100010011100100101",
8962 => "100110001111111010111111",
8963 => "100110101001001100101101",
8964 => "100111000001111110111100",
8965 => "100111100011101010100101",
8966 => "100111001100101111101110",
8967 => "101000000101101010011000",
8968 => "101110000010111100010100",
8969 => "110111101100111000111111",
8970 => "000001000000110101000101",
8971 => "001001100010011101011001",
8972 => "010001010101000000101000",
8973 => "010101111010101001100100",
8974 => "010110011010110101001100",
8975 => "010100111100111100100110",
8976 => "010011101100111100001000",
8977 => "010010110110101111100010",
8978 => "010000101110100010101110",
8979 => "001101001011001001001100",
8980 => "001011001110001111100011",
8981 => "001100110010111110110000",
8982 => "010000001111101101111100",
8983 => "010011010111111101111100",
8984 => "010110000000001100111110",
8985 => "011000110010111101100101",
8986 => "011011000101100101100011",
8987 => "011011101011000100000101",
8988 => "011010000101000000010100",
8989 => "010101110011100011010010",
8990 => "001111101010110111100000",
8991 => "001010100110111100110011",
8992 => "001000100101000101000111",
8993 => "001001011000100111111000",
8994 => "001011101010011001111100",
8995 => "001110001010110100111010",
8996 => "010001010000011011100000",
8997 => "010100001101111010100000",
8998 => "010100101101010011010010",
8999 => "010011000000011100011100",
9000 => "001111101100000110010010",
9001 => "001001101101011001100010",
9002 => "000010000101111110101111",
9003 => "111000100001001010011100",
9004 => "101011111100010110101100",
9005 => "100010011010000111011011",
9006 => "100000100111011010000001",
9007 => "100001011010101011011111",
9008 => "100001000100000110010111",
9009 => "100001000101001110110101",
9010 => "100001000111101110011111",
9011 => "100001101000010011010000",
9012 => "100101011011101101000100",
9013 => "101100010010001001110010",
9014 => "110011100010110100110100",
9015 => "111001100011001010011101",
9016 => "111101111100010101110000",
9017 => "000001100011110110111000",
9018 => "000100011110100011111011",
9019 => "000101010100100001011010",
9020 => "000100101100001110001010",
9021 => "000100111100111101111001",
9022 => "000101110100011111100111",
9023 => "000100111101000000101001",
9024 => "000001111001110100011110",
9025 => "111110000001100101100011",
9026 => "111010010111101101011110",
9027 => "110111001001011101011000",
9028 => "110100010100011111101110",
9029 => "110010101010001111000110",
9030 => "110010101101000011101000",
9031 => "110011010111000001001110",
9032 => "110100011010010111001010",
9033 => "110111001110000000100010",
9034 => "111011010000111000010100",
9035 => "111110100101010001000011",
9036 => "000000100010001011010010",
9037 => "000001010011111101100100",
9038 => "000001010001010100000011",
9039 => "000000110101111011010000",
9040 => "000000000001100110000010",
9041 => "111111010110110000001010",
9042 => "111111111011111011010000",
9043 => "000000100100011001011011",
9044 => "111101110101001101100100",
9045 => "110111110010011100011010",
9046 => "110011010100010111111110",
9047 => "110010010000111010110010",
9048 => "110001001100000101101110",
9049 => "101111010001110000100110",
9050 => "101111011011101100100000",
9051 => "110010001101011100110000",
9052 => "110101101000100111001000",
9053 => "111000001001011010000001",
9054 => "111010000101101100001111",
9055 => "111101110001001000010111",
9056 => "000011110100110100110000",
9057 => "001001101111101111010101",
9058 => "001101111010100101101010",
9059 => "010000111011001101100000",
9060 => "010011010011111010000010",
9061 => "010101000101000101111000",
9062 => "010110010011110100111110",
9063 => "010111100001111010011110",
9064 => "011001000110011000110011",
9065 => "011010001001100110111000",
9066 => "011010000101011001011101",
9067 => "011001101111010101111011",
9068 => "011000111111011001000001",
9069 => "010110111010101111101110",
9070 => "010101000000001000000110",
9071 => "010100011000000000110000",
9072 => "010010001100011110101010",
9073 => "001101010010000100000100",
9074 => "001001010010101110111100",
9075 => "000111101100100011001010",
9076 => "000101110100010100100000",
9077 => "000010001011001111010001",
9078 => "111101101001011011100000",
9079 => "111010010111000111101010",
9080 => "111010011100100110001011",
9081 => "111101010000101101101101",
9082 => "000000000100111110111111",
9083 => "000000111100000110010110",
9084 => "111111011001000110010101",
9085 => "111100001000100011011110",
9086 => "110111100000010011011001",
9087 => "110001110001010001101000",
9088 => "101101000011101111111000",
9089 => "101010111110111110000100",
9090 => "101010100101001110010110",
9091 => "101010101000001111101100",
9092 => "101010010011111110100000",
9093 => "101001010011000010010110",
9094 => "101000101010101000010100",
9095 => "101001010011101100101000",
9096 => "101010111100010111010100",
9097 => "101101000001001001101110",
9098 => "101110110111011101100100",
9099 => "110000011101000010110110",
9100 => "110010010110010001011010",
9101 => "110100010010111010010101",
9102 => "110101100100000011010010",
9103 => "110110010111100000001111",
9104 => "111000010110001010111000",
9105 => "111100110011101001101101",
9106 => "000010001101010111010101",
9107 => "000101111100111000010000",
9108 => "000111111000010011010000",
9109 => "001001011011011100010011",
9110 => "001011000010110010110010",
9111 => "001011110101101110010100",
9112 => "001011100100001100000100",
9113 => "001100000101011010101010",
9114 => "001110110010110111011010",
9115 => "010010001001000111101100",
9116 => "010100001010010000101110",
9117 => "010101001000001101011010",
9118 => "010110010111111000011000",
9119 => "011000010011100101011101",
9120 => "011010001110011001101001",
9121 => "011011001010100101011011",
9122 => "011010111001111100111101",
9123 => "011010100000000110111011",
9124 => "011010101001000010111001",
9125 => "011010010101111111000101",
9126 => "011001100101010110111001",
9127 => "011001000001101111101101",
9128 => "010110010100101001111110",
9129 => "001111111111100000000000",
9130 => "001001101101101100010111",
9131 => "000101100100011100100110",
9132 => "000000011011111011000000",
9133 => "111001001101110000110011",
9134 => "110010110110011100111100",
9135 => "101101110001001110110100",
9136 => "100111101110001011110011",
9137 => "100010010110101101101011",
9138 => "100001001001000010100101",
9139 => "100010010000011010001011",
9140 => "100010010100010001110111",
9141 => "100010000111000000000100",
9142 => "100010101111010000100100",
9143 => "100011111100110111101011",
9144 => "100110101011001001000101",
9145 => "101010111100000110101010",
9146 => "101111001011011100011110",
9147 => "110011001001010101111100",
9148 => "110111011100010011100110",
9149 => "111011110001011101010101",
9150 => "111111101110001001111110",
9151 => "000011100111000001001001",
9152 => "000111011000001000001100",
9153 => "001001110101000001101011",
9154 => "001010100001110111010001",
9155 => "001001100111001001000011",
9156 => "000101011011100000111000",
9157 => "111101110010100101111000",
9158 => "110110111010011011001100",
9159 => "110011111010110111001000",
9160 => "110011001111001010011110",
9161 => "110011001111111110010010",
9162 => "110101100111011010101100",
9163 => "111011111010000101010110",
9164 => "000011110100110111100000",
9165 => "001010000010110001001010",
9166 => "001111000001001110011110",
9167 => "010100011101101001001010",
9168 => "011000111100100011001101",
9169 => "011010100101111101000111",
9170 => "011010010010100110001001",
9171 => "011001100011001011010011",
9172 => "011000110010110100111001",
9173 => "010111100101110011000100",
9174 => "010100010010000101110000",
9175 => "001101110100110010011100",
9176 => "000101110110001111101100",
9177 => "111110010011111010101010",
9178 => "110111110010111011111101",
9179 => "110010000101001101111000",
9180 => "101011111011000010100000",
9181 => "100110000000010010100110",
9182 => "100011110010101010101011",
9183 => "100101000011000001101101",
9184 => "100110100110101110011100",
9185 => "101000110111011100010100",
9186 => "101100110000000111111000",
9187 => "110001010100010101010000",
9188 => "110110100110001010110000",
9189 => "111010110110100010111111",
9190 => "111011100001011110000001",
9191 => "111011010010001011010110",
9192 => "111101101001111001100001",
9193 => "000000100101100000110110",
9194 => "000000101110101011000010",
9195 => "111110110111011110011000",
9196 => "111110010011010001010100",
9197 => "111111110000000111100010",
9198 => "000000110000011101111011",
9199 => "000000101011101010100110",
9200 => "000001110010011001001100",
9201 => "000101000011110010110100",
9202 => "001000011100100001000000",
9203 => "001001000110010111010000",
9204 => "000110110011011101110001",
9205 => "000011111010010011100111",
9206 => "000001110011110101010010",
9207 => "000000011111100000010011",
9208 => "111111111000000011101001",
9209 => "111111001111101000111000",
9210 => "111110001100010010000000",
9211 => "111101110001101100100100",
9212 => "111110110110100000111100",
9213 => "000000011001010111101111",
9214 => "000000011101100011000100",
9215 => "111111011110101011001100",
9216 => "000000101001100101101101",
9217 => "000100110011011101000100",
9218 => "001000101111001010000111",
9219 => "001010001111000011010110",
9220 => "001010011101001101111001",
9221 => "001010111000101101100101",
9222 => "001010111110000111100001",
9223 => "001001101000111100100110",
9224 => "000111011101110001000111",
9225 => "000101100100100100010011",
9226 => "000011110100100111001011",
9227 => "000001011001011001111101",
9228 => "111110000011100101111010",
9229 => "111010011101010100111000",
9230 => "110111001110111101000011",
9231 => "110100101001011101000101",
9232 => "110100000100000010001101",
9233 => "110110110001100100111001",
9234 => "111011000010001010000110",
9235 => "111110000011111110100101",
9236 => "111111010011100001010110",
9237 => "111110101101011000100100",
9238 => "111011011010011101000110",
9239 => "110110011000000111101000",
9240 => "110011000000101000001000",
9241 => "110011101101111000000000",
9242 => "110111110001001011101111",
9243 => "111101001010110110001011",
9244 => "000011000111010111010000",
9245 => "001001101100100000001100",
9246 => "010000000110010101000010",
9247 => "010101001001110011110110",
9248 => "011000111100111101010001",
9249 => "011011010111010010100111",
9250 => "011011011000010101001001",
9251 => "011010000000011111001001",
9252 => "011001001111110011011001",
9253 => "011000101001010100101101",
9254 => "010111101011011110010110",
9255 => "010111100100010010110000",
9256 => "010111101100011110011010",
9257 => "010110000010101000111110",
9258 => "010011100101100010010110",
9259 => "010010100101110101111010",
9260 => "010010000000010110101110",
9261 => "001111001000001010101010",
9262 => "001000111111101101111110",
9263 => "111111110000001101010100",
9264 => "110100110000110010011100",
9265 => "101011000111001111000110",
9266 => "100100101101111011001011",
9267 => "100001100101100100001101",
9268 => "100001011100000110001011",
9269 => "100010101000101011101111",
9270 => "100011100001111010100011",
9271 => "100101001010011000111111",
9272 => "101000010011111010001000",
9273 => "101011111001101111011000",
9274 => "110000001010001111000010",
9275 => "110101111000000000100101",
9276 => "111011010110001001110000",
9277 => "111101111011010100001111",
9278 => "111101100001110000001101",
9279 => "111100010001000100001111",
9280 => "111010110110100001010011",
9281 => "111000001011101010000110",
9282 => "110100100111011000110101",
9283 => "110001101011111011110100",
9284 => "101111010010101110101010",
9285 => "101100110101101001001000",
9286 => "101011001001100011110000",
9287 => "101010011110011111010100",
9288 => "101001110101111101010010",
9289 => "101010010001000101111010",
9290 => "101101110100100111100010",
9291 => "110011001100110111011000",
9292 => "110111101100000111100111",
9293 => "111011010010100000011001",
9294 => "111111000111011001101111",
9295 => "000011001011010000011011",
9296 => "000110100100101000001000",
9297 => "001000111010011110010000",
9298 => "001011101010101111001110",
9299 => "001111110000010010010000",
9300 => "010100001101000010100100",
9301 => "011000101111001010010011",
9302 => "011100011100000011000011",
9303 => "011101010100000100111011",
9304 => "011100100001001110101100",
9305 => "011100010110100001110011",
9306 => "011100011110100011100011",
9307 => "011011101110101000110101",
9308 => "011000010111011100010011",
9309 => "010001100001011110110010",
9310 => "001001110001101111011110",
9311 => "000010110010010011100110",
9312 => "111011011110110000111100",
9313 => "110100110110010111010010",
9314 => "110001110110100011001000",
9315 => "110011011101010110001110",
9316 => "110110100111010101101011",
9317 => "110110110111100010001011",
9318 => "110101000110000011010101",
9319 => "110101111000111101100000",
9320 => "111001001011101111010001",
9321 => "111011111101000100100010",
9322 => "111101111110010000011111",
9323 => "000000000111010101100110",
9324 => "000001111011100000010010",
9325 => "000010000011110100001111",
9326 => "111111110011100001100000",
9327 => "111100101101101001011010",
9328 => "111010111010011010011010",
9329 => "111010101100101011101000",
9330 => "111010101101001101010010",
9331 => "111001101000000111000001",
9332 => "111000010100010111000011",
9333 => "110111111101011000001000",
9334 => "110110111000110101111010",
9335 => "110100001000111000110100",
9336 => "110001111011100111101010",
9337 => "110001110001010100011010",
9338 => "110011100001010011111100",
9339 => "110110011000000010001110",
9340 => "111000010001100101011000",
9341 => "111000100001100011110110",
9342 => "111000111110000010110101",
9343 => "111010101011111111011101",
9344 => "111101000001001010000000",
9345 => "111110100100101011111100",
9346 => "111110010010011101110110",
9347 => "111101000111101100010111",
9348 => "111100101110000011011111",
9349 => "111100111010101011101001",
9350 => "111100011011000111111101",
9351 => "111010100011101010011101",
9352 => "111000100010100110110000",
9353 => "111000110010011101110111",
9354 => "111011011101110011001101",
9355 => "111110010011110110001100",
9356 => "000000000101111000001000",
9357 => "000001000111000001001000",
9358 => "000001011000011011010110",
9359 => "000000101110101101000111",
9360 => "111111111010110101001111",
9361 => "000000001100111101110111",
9362 => "000010000000100000101101",
9363 => "000101000110101001010110",
9364 => "001000101010101011011101",
9365 => "001010111100110011101000",
9366 => "001011001000011111101110",
9367 => "001010000010011001011101",
9368 => "001000010010111000011111",
9369 => "000110101111111010011010",
9370 => "000110101111001000000011",
9371 => "001000000100101000001001",
9372 => "001001111100000001001001",
9373 => "001100101110011001010110",
9374 => "010000001100011001111110",
9375 => "010010101111111101011000",
9376 => "010100100101001111101100",
9377 => "010111110000001101010110",
9378 => "011011010011000110010011",
9379 => "011011110011101101010001",
9380 => "011010000000101010011011",
9381 => "011001000110101111100101",
9382 => "011000110011001110101111",
9383 => "010111111100000101110000",
9384 => "010111000101001011001110",
9385 => "010110010110101001101100",
9386 => "010110000001011010011010",
9387 => "010101111101100000101010",
9388 => "010101001000101001000000",
9389 => "010100100001100001001000",
9390 => "010100001101111110010000",
9391 => "010000101101110001011110",
9392 => "001001001011010011100101",
9393 => "000000011011000100011100",
9394 => "111000000011110111011100",
9395 => "110001001100001100001010",
9396 => "101100011100100010011110",
9397 => "101000110001100011001000",
9398 => "100110010001010000101111",
9399 => "100101101110000110000110",
9400 => "100110001010001011100011",
9401 => "100111010010111110101001",
9402 => "101010100011101110110110",
9403 => "101111110111010111011010",
9404 => "110101010000000110011100",
9405 => "111001111100001101111100",
9406 => "111101110000010001111101",
9407 => "111110011101100111001110",
9408 => "111011011001000101000010",
9409 => "110111100101111111111110",
9410 => "110100000011011000101100",
9411 => "110000010100001101100000",
9412 => "101111000001111000111100",
9413 => "110000100111110111111000",
9414 => "110001010011111010110100",
9415 => "101111001100010011000000",
9416 => "101010110100100011110010",
9417 => "100110010001010110100101",
9418 => "100100011000101101010111",
9419 => "100100110101011011111101",
9420 => "100101110111000110001011",
9421 => "100111000000110010011110",
9422 => "100111011011110011000101",
9423 => "101000100101001100010100",
9424 => "101101101100000100110100",
9425 => "110101011100111111001000",
9426 => "111100101011111001011101",
9427 => "000011110000001101101010",
9428 => "001100011111110110100010",
9429 => "010110001001111010101100",
9430 => "011100100001010001110011",
9431 => "011101111001101001101111",
9432 => "011101111000001111010101",
9433 => "011101111100000011011101",
9434 => "011101001001011000101111",
9435 => "011100001000111110010011",
9436 => "011001011110100011100111",
9437 => "010100010011101110010010",
9438 => "001111101100001001110110",
9439 => "001100001001111000011010",
9440 => "001000110101000011000000",
9441 => "000110110010100001101000",
9442 => "000101001110110100111110",
9443 => "000100001001111111110010",
9444 => "000101101000101010000001",
9445 => "001000110000110100111000",
9446 => "001011111100010100011011",
9447 => "001110011010011100011100",
9448 => "001110001110110000100000",
9449 => "001011001011000010110100",
9450 => "000110101110100010111010",
9451 => "000010100101111000000000",
9452 => "000000110110001001011101",
9453 => "111111111101101001010010",
9454 => "111100010100111100011011",
9455 => "110110111101101101010000",
9456 => "110011110000100110110010",
9457 => "110100000111100101100000",
9458 => "110101010111010101100010",
9459 => "110100101100010001110101",
9460 => "110100010101011100111000",
9461 => "110101110110000100111010",
9462 => "110101001011000100100111",
9463 => "110000101011101010110100",
9464 => "101011101000011010010100",
9465 => "101000100000000011100000",
9466 => "100111111000010001000011",
9467 => "101000110011100111101110",
9468 => "101010010011001000011010",
9469 => "101100110111101101110100",
9470 => "110000001001000011111100",
9471 => "110011011110010110110010",
9472 => "110111100110100011010011",
9473 => "111100011101000110111101",
9474 => "000001011011011000111100",
9475 => "000110001000011010001001",
9476 => "001001001110000010000011",
9477 => "001001011011001101000110",
9478 => "000110100110011100110110",
9479 => "000010001100110111110010",
9480 => "111110111010100101100011",
9481 => "111101011101000010010110",
9482 => "111011111111001010001010",
9483 => "111001001101000010010001",
9484 => "110101111100000010001000",
9485 => "110100001111001011011100",
9486 => "110100000000111111010101",
9487 => "110010101011010011110010",
9488 => "101111111001011111110010",
9489 => "101110100000111100001010",
9490 => "110000010001010001110110",
9491 => "110100000011101010001111",
9492 => "111000010101101001001100",
9493 => "111101010001111111011100",
9494 => "000010110101001001110001",
9495 => "000111011100101000100000",
9496 => "001010001110010100101100",
9497 => "001011000001011011010111",
9498 => "001010001011111001110010",
9499 => "001000111010011110010001",
9500 => "000111100110011111010010",
9501 => "000110001111001110011001",
9502 => "000101000001001001101010",
9503 => "000011011110011100010011",
9504 => "000010100110011011001110",
9505 => "000011110001110100111000",
9506 => "000101110110011001000100",
9507 => "000111111010010001010010",
9508 => "001001110101100110000010",
9509 => "001011001100110011110010",
9510 => "001100110001100111110100",
9511 => "001101111101000110011100",
9512 => "001101011111110101010110",
9513 => "001101100001000001111010",
9514 => "001111010001101010011110",
9515 => "010010000011010000011010",
9516 => "010110001101101000101010",
9517 => "011001111010110000111111",
9518 => "011010011110011101000011",
9519 => "011001001010100110111010",
9520 => "011000001010010110000001",
9521 => "010111101010101000100010",
9522 => "010110011100110101001010",
9523 => "010011010011010101000100",
9524 => "001110110101111111110110",
9525 => "001001010100011110010000",
9526 => "000010011010101000011011",
9527 => "111100010101110000000010",
9528 => "111001010101110010100101",
9529 => "111001010110000100111100",
9530 => "111011000010101111001100",
9531 => "111100100100100101010011",
9532 => "111101111101111100110000",
9533 => "000000100111110101101010",
9534 => "000011101101000101101001",
9535 => "000101001001010010011011",
9536 => "000011100101111111110111",
9537 => "111111101101010110101100",
9538 => "111100001010011100001001",
9539 => "111001111000111010101011",
9540 => "111000000110000101100110",
9541 => "110110110011110110010001",
9542 => "110101111011011111011101",
9543 => "110100110010100110111101",
9544 => "110001010010001001110000",
9545 => "101010001000010100011110",
9546 => "100100000011000110101001",
9547 => "100011001000100101001110",
9548 => "100100010001010010100101",
9549 => "100100101011100100110001",
9550 => "100101000100101010100010",
9551 => "100101110100000000111111",
9552 => "100110101000101011011111",
9553 => "100110111111011100011111",
9554 => "101000101110111000000010",
9555 => "101110101111001100110000",
9556 => "110101111011011101111000",
9557 => "111010011010001101101100",
9558 => "111110010100000101101100",
9559 => "000010110001001011110110",
9560 => "000101011101100101111100",
9561 => "000110001011011001110011",
9562 => "000110010010110101000011",
9563 => "000110110000100100100100",
9564 => "001000010111101001010010",
9565 => "001010110110101011111000",
9566 => "001100110000100100000000",
9567 => "001101011100110010011000",
9568 => "001101101011011011000110",
9569 => "001101010111000111111110",
9570 => "001100000100000000100000",
9571 => "001010111100001100010001",
9572 => "001010010000011010111011",
9573 => "001001100100000001001011",
9574 => "001010110100100100010011",
9575 => "001111000001110010011000",
9576 => "010011101011110010101110",
9577 => "010110011100111100110000",
9578 => "010111100001111010111110",
9579 => "011000110010100101011111",
9580 => "011010100010110001011011",
9581 => "011010111101101111011101",
9582 => "011010000010110111100111",
9583 => "011001001100110100001111",
9584 => "011000110000111111110001",
9585 => "010111110001011110110010",
9586 => "010011001111010011100100",
9587 => "001010011101101111011111",
9588 => "000001111011101111011110",
9589 => "111100000010011100000000",
9590 => "110110101110110010000010",
9591 => "110000011011111110011110",
9592 => "101001101101110100001000",
9593 => "100101100010001000110111",
9594 => "100101001001111110000101",
9595 => "100101000101100011101011",
9596 => "100100001101011000110111",
9597 => "100101000001011010011000",
9598 => "100110111010101011011100",
9599 => "100111110011010111001001",
9600 => "100111100101110110101011",
9601 => "100111011101100010101111",
9602 => "101001001111101100100110",
9603 => "101100110100001011011100",
9604 => "110000001010111000100100",
9605 => "110011011011000111100000",
9606 => "110111100111101100011011",
9607 => "111011110101101110001000",
9608 => "111110110110111000101111",
9609 => "000000110111100000101110",
9610 => "000010111001100010001000",
9611 => "000101111000011111101111",
9612 => "001001011100110000010010",
9613 => "001011000100101000101000",
9614 => "001000100110000010100010",
9615 => "000011010101011000101101",
9616 => "111101110110110010100000",
9617 => "111001010001001111110010",
9618 => "110101110100010111101000",
9619 => "110011000000000001111110",
9620 => "110001000101000110001100",
9621 => "110001101011100010110100",
9622 => "110100111101111010000111",
9623 => "111010010101110100010010",
9624 => "000000110110000000011001",
9625 => "000101110111001111110011",
9626 => "001001110011000010000000",
9627 => "001111011110011110101110",
9628 => "010100111111111000010100",
9629 => "010111010101011011110100",
9630 => "010111100011111000101110",
9631 => "010110111001000111110100",
9632 => "010100111101000111000000",
9633 => "010001100010111100010010",
9634 => "001101101101111000101100",
9635 => "001011101001010011100011",
9636 => "001011101010001101101000",
9637 => "001100001100101100111110",
9638 => "001100010100011001111100",
9639 => "001011000111101110100001",
9640 => "001000011001011010011000",
9641 => "000101001010011101011111",
9642 => "000010000001101011101111",
9643 => "000000000110010111001110",
9644 => "000000000110101110100010",
9645 => "000000011111001111011000",
9646 => "000000101110111101101011",
9647 => "000001111011111101000111",
9648 => "000011010100010101000101",
9649 => "000011011101011101101111",
9650 => "000010111010101110111110",
9651 => "000010110000101000101001",
9652 => "000010010000001100101100",
9653 => "000000000010001000110011",
9654 => "111100110110011001100000",
9655 => "111001110011111000010000",
9656 => "110101111000000010100010",
9657 => "110000100100001010011010",
9658 => "101011111100000010000000",
9659 => "101010010111110001110100",
9660 => "101100001010110011011000",
9661 => "101111010001001000011100",
9662 => "110001110111011001001100",
9663 => "110100101111100101110101",
9664 => "111001011101001110100100",
9665 => "111111011100001111111110",
9666 => "000100001011110001101001",
9667 => "000110010010000001010000",
9668 => "000111000010000011101010",
9669 => "001000000111101001000010",
9670 => "001001011101110001100011",
9671 => "001001101011111010110101",
9672 => "001000010010100010001111",
9673 => "000110101101110110110011",
9674 => "000101001001010001011011",
9675 => "000001101010111000101001",
9676 => "111100011000001111111010",
9677 => "110110111100000001010011",
9678 => "110010100011100010101100",
9679 => "110000110001010101100110",
9680 => "110000111110101101101100",
9681 => "110000111000101100001010",
9682 => "110001011001111110010100",
9683 => "110011110000110110110110",
9684 => "110110000101000001100001",
9685 => "110111110111101000011110",
9686 => "111010100001011001000000",
9687 => "111101011001011000000000",
9688 => "111110111011010010011101",
9689 => "111111011010001100111110",
9690 => "000000101010101111001100",
9691 => "000011011110101111100111",
9692 => "000110000101001001110001",
9693 => "000110110001010011100101",
9694 => "000110100011001010000101",
9695 => "000110100000110000110001",
9696 => "000100110100101100001111",
9697 => "111111101100000010001010",
9698 => "111000111100111010000010",
9699 => "110011001000010111110100",
9700 => "101110101101010100000100",
9701 => "101101000001101000110100",
9702 => "101111101010111111101100",
9703 => "110100101011011010001010",
9704 => "111001110011111010000011",
9705 => "000000001001001111001110",
9706 => "001000000011001101110100",
9707 => "010000001111000100000010",
9708 => "011000011110010110111101",
9709 => "011110101100011010110101",
9710 => "011111101011100000000101",
9711 => "011101100000101000100111",
9712 => "011011111100111010110000",
9713 => "011010110110101111011001",
9714 => "011010000000111010110101",
9715 => "011000110111010101011100",
9716 => "010100111100000011111010",
9717 => "001111011101101011100110",
9718 => "001011001011100011100110",
9719 => "000111001011001101101010",
9720 => "000011001111000101101011",
9721 => "111111111101110010110011",
9722 => "111011110001011011001111",
9723 => "110110100000001111100000",
9724 => "110001100110110111100110",
9725 => "101101111000011110010000",
9726 => "101011101010000110110110",
9727 => "101000111001110110010000",
9728 => "100100011011000001001100",
9729 => "100001111100011110010010",
9730 => "100011000110110100110100",
9731 => "100100010101010000111111",
9732 => "100100110010110110111011",
9733 => "100111110100101101100001",
9734 => "101110001111110100111110",
9735 => "110100100111101010101000",
9736 => "111000001011000110100111",
9737 => "111001110111110101100110",
9738 => "111011011000010011100010",
9739 => "111100101010000001101100",
9740 => "111100111000011110110111",
9741 => "111011100101011001110101",
9742 => "111010000111110010111010",
9743 => "111010001110111011100001",
9744 => "111010110111000000100000",
9745 => "111010010001000111001100",
9746 => "111000101100110000000110",
9747 => "110111110010110100011001",
9748 => "111001110010111101100101",
9749 => "111110000111010000011101",
9750 => "000000110100101011100100",
9751 => "000001000011001101110101",
9752 => "000001011011000101100000",
9753 => "000011001000101100001011",
9754 => "000110000011111011001101",
9755 => "001001001010011000001111",
9756 => "001010011100001110001101",
9757 => "001001111111011111011101",
9758 => "001001100000110010101010",
9759 => "001001101001110010010111",
9760 => "001010101110010010010010",
9761 => "001100011110000100100100",
9762 => "001110100010101000001110",
9763 => "010010110101000010100110",
9764 => "011001110101011111010001",
9765 => "011111001011111011101111",
9766 => "011111101101010011110001",
9767 => "011101110110011000100000",
9768 => "011100111010001101011100",
9769 => "011100010100000110011001",
9770 => "011000110110100001001101",
9771 => "010001110001000111001100",
9772 => "001010101111011011011000",
9773 => "000110111000101111010001",
9774 => "000101011110011100001011",
9775 => "000100101100100111110110",
9776 => "000011110111100011011100",
9777 => "000011101100100010010101",
9778 => "000101000010010100111010",
9779 => "000110100110001010100010",
9780 => "000110011000011000100011",
9781 => "000100011001011001101100",
9782 => "000001100010000111110100",
9783 => "111101011001011000101000",
9784 => "110110010000000011011101",
9785 => "101100011010011010101000",
9786 => "100100010111010101010101",
9787 => "100001010011011000101011",
9788 => "100001001101001011101110",
9789 => "100001010001100001111000",
9790 => "100001101100111110010001",
9791 => "100100101001111011101111",
9792 => "101010011001011000111110",
9793 => "101111010111111001111010",
9794 => "110001110111001111111110",
9795 => "110100100100110100010100",
9796 => "110111111011111101011010",
9797 => "111001011111010101101100",
9798 => "111001110110111001111000",
9799 => "111010111101110101000000",
9800 => "111011100100100110011110",
9801 => "111010001110101000010001",
9802 => "111001000111011111101110",
9803 => "111010001101100011010011",
9804 => "111010101100100111110101",
9805 => "110111101000111111011110",
9806 => "110011010111010000011000",
9807 => "110000111001111011100010",
9808 => "101111001100001101101000",
9809 => "101100101110000011000010",
9810 => "101011000110001110000010",
9811 => "101011110010101011101010",
9812 => "101101101100101011000100",
9813 => "110000011001001010110000",
9814 => "110100111011000101101000",
9815 => "111010100000000000100100",
9816 => "111111011100000110000011",
9817 => "000011110010011001000010",
9818 => "000111111010010010011100",
9819 => "001011000111111111001100",
9820 => "001100101111010010001100",
9821 => "001101000110111101110100",
9822 => "001101000001011110111100",
9823 => "001100111101000100011010",
9824 => "001101100110010001110100",
9825 => "001110001010000001111110",
9826 => "001100000101101111101110",
9827 => "001000011010100100101110",
9828 => "000110100011010100101010",
9829 => "000101110101100110111111",
9830 => "000100001100100001010100",
9831 => "000010101001101001001111",
9832 => "000011010110110101010110",
9833 => "000111000011010111001110",
9834 => "001011111011110011101010",
9835 => "010000010001110001010000",
9836 => "010101000010111000011010",
9837 => "011010000101111001101011",
9838 => "011101010110011111000111",
9839 => "011110010011000001010010",
9840 => "011101100100001110101111",
9841 => "011100100010001100100101",
9842 => "011100001010011101000101",
9843 => "011011010101011010001111",
9844 => "011001111111111001100110",
9845 => "011001000111001100110001",
9846 => "011000001110110011101101",
9847 => "010111011011011111101010",
9848 => "010101100010010000101100",
9849 => "010000000011000011010000",
9850 => "001000110101011011011100",
9851 => "000010111010001010100000",
9852 => "111101101110010111101010",
9853 => "111001011100100001110000",
9854 => "110111000110000011111110",
9855 => "110101101001001101111000",
9856 => "110100000101010110011000",
9857 => "110010100101100011101110",
9858 => "110001110011101110011000",
9859 => "110010000000110100011110",
9860 => "110010100011000001001110",
9861 => "110011100011001011110100",
9862 => "110101101001000011101010",
9863 => "110111011111111111110010",
9864 => "110110100010101101000101",
9865 => "110001011000010011101110",
9866 => "101001111010100100101000",
9867 => "100100100100000010100101",
9868 => "100011010111001110000101",
9869 => "100100010000110011000001",
9870 => "100101000001101101100101",
9871 => "100101101010100111101101",
9872 => "100110101110000101111001",
9873 => "100111100111000101111010",
9874 => "100111110000010110010111",
9875 => "100111101010000100101101",
9876 => "101000100100110101000100",
9877 => "101011011110010101110010",
9878 => "101110111100010011101000",
9879 => "110001001101011111000100",
9880 => "110100010001001111000010",
9881 => "111001100101101110010100",
9882 => "111110100010110100001101",
9883 => "000010010001101100101110",
9884 => "000111010000110011101101",
9885 => "001110110000100011101100",
9886 => "010111001110001101101110",
9887 => "011101000111010111010110",
9888 => "011110110000011010110110",
9889 => "011110000001101011111001",
9890 => "011100001001110101111101",
9891 => "011001111100101111011111",
9892 => "011000111111110011001101",
9893 => "011000011001001101101000",
9894 => "010111101110111111100110",
9895 => "011001001100000011101001",
9896 => "011011011001110011100110",
9897 => "011011011000110110001101",
9898 => "011010011101101111111000",
9899 => "011010001001011011111011",
9900 => "011001101100100000010111",
9901 => "011001011010100001001101",
9902 => "011001011001011111101111",
9903 => "011000110111101111100101",
9904 => "011000100010100000110111",
9905 => "010111111110000101101100",
9906 => "010100100010101010001000",
9907 => "001110110101111001011000",
9908 => "001010001110000100010110",
9909 => "000110111110010001110110",
9910 => "000011010100101001101110",
9911 => "111111000010000101001010",
9912 => "111010111000111001111001",
9913 => "110111011010101001001001",
9914 => "110100001100110010010100",
9915 => "110000100000111100110010",
9916 => "101101000011000100011000",
9917 => "101011001110100000111010",
9918 => "101011010011110010010110",
9919 => "101011110000000000110100",
9920 => "101010101001010100111010",
9921 => "101000001010001010010100",
9922 => "100101010011010010000111",
9923 => "100010011001001000101101",
9924 => "100000101110111101111000",
9925 => "100000110111001001110110",
9926 => "100001101011001111111001",
9927 => "100100010110011101110101",
9928 => "101010000100101111110010",
9929 => "110000011011000100111110",
9930 => "110101011101010100100101",
9931 => "111001100011100011011110",
9932 => "111101001001100111010101",
9933 => "000000001010010110100000",
9934 => "000001100110110011111000",
9935 => "000000011010111101010001",
9936 => "111100011011101001100110",
9937 => "110110011011000100010100",
9938 => "110001000011010011001110",
9939 => "101110010000111100000000",
9940 => "101100111001011010001110",
9941 => "101100010100100000011110",
9942 => "101101101000000001001100",
9943 => "110001001000110000100010",
9944 => "110101101110111011001011",
9945 => "111000111101111001000101",
9946 => "111001111100110001010010",
9947 => "111010100110111000100011",
9948 => "111011100001110011011110",
9949 => "111100001010011101101001",
9950 => "111101000011001111111100",
9951 => "111101101101110110111001",
9952 => "111101110001010011011110",
9953 => "111110011100110000111100",
9954 => "111111110000110001110100",
9955 => "000000001101110111101111",
9956 => "111110101000001010101100",
9957 => "111011000000001101111101",
9958 => "110111000001001100001111",
9959 => "110100001010111000100100",
9960 => "110010101111010001001110",
9961 => "110010110101001100111100",
9962 => "110100001000110110000010",
9963 => "110110011001010111010111",
9964 => "111001111110111001011010",
9965 => "111110100111110010111000",
9966 => "000011000111000001111110",
9967 => "000110011101010011000100",
9968 => "001001010010001000101010",
9969 => "001101010000111100110100",
9970 => "010010000110110010010000",
9971 => "010101111010000010001100",
9972 => "010111110110000000100110",
9973 => "011000001011010111010011",
9974 => "011000000101111111001111",
9975 => "011000100010111011101001",
9976 => "011000100011110101000101",
9977 => "010111011110010111011000",
9978 => "010110001100100000101100",
9979 => "010101011000001010101000",
9980 => "010101010001111101000010",
9981 => "010101101000100101010010",
9982 => "010101011101110011001000",
9983 => "010100101011000011100010",
9984 => "010100010100011000111110",
9985 => "010100111101001011100100",
9986 => "010101011010001001101010",
9987 => "010100101100110101000010",
9988 => "010100000110110111110010",
9989 => "010100000001110010101000",
9990 => "010010111100001010001100",
9991 => "010001000000101010001100",
9992 => "001111001011111100010110",
9993 => "001101010100101111000110",
9994 => "001011010101011011000110",
9995 => "001000110011010001111010",
9996 => "000101010101000011101110",
9997 => "000000011111100101010100",
9998 => "111001111110111000111100",
9999 => "110100100101110111000001",
10000 => "110001001101000111101000",
10001 => "101011000011001111000100",
10002 => "100011011100011010110101",
10003 => "100001100010000111011101",
10004 => "100011011101110111101101",
10005 => "100011100110011111100111",
10006 => "100011011110001100101101",
10007 => "100100110011111100111110",
10008 => "100101110011111111111011",
10009 => "100110011011011011010110",
10010 => "100111000100100011100001",
10011 => "100110100100111000100100",
10012 => "100110111100000110100100",
10013 => "101101001111111001001110",
10014 => "111000100110001101111110",
10015 => "000001110101011101101000",
10016 => "000110111000111000011100",
10017 => "001010101010111001010011",
10018 => "001100011100011110000110",
10019 => "001010011011001101110110",
10020 => "000110100010000100000000",
10021 => "000100001010101101000001",
10022 => "000101101001111111000000",
10023 => "001010001010101101000001",
10024 => "001110111100101111001100",
10025 => "010010110011001010000110",
10026 => "010100110101100001000110",
10027 => "010100100110100111101110",
10028 => "010100000011011101011100",
10029 => "010100011111010011110110",
10030 => "010101000010100010010010",
10031 => "010100110111001111111010",
10032 => "010100010000101110011110",
10033 => "010100111001110010110100",
10034 => "010110110101110000011110",
10035 => "010111100001000101100110",
10036 => "010111000000101101010000",
10037 => "010111010100001110110000",
10038 => "010111101001001001001100",
10039 => "010110111100110000001110",
10040 => "010101011001000101101100",
10041 => "010010001110001010001110",
10042 => "001101000100001011001110",
10043 => "000101111011000100100100",
10044 => "111100010001101110000011",
10045 => "110001111100010100010110",
10046 => "101010111011000001000010",
10047 => "101000101111100100100000",
10048 => "101001011100110001111110",
10049 => "101011001101011010000010",
10050 => "101101110010010110000000",
10051 => "110000011001001011110010",
10052 => "110010000000110101010010",
10053 => "110011010011000001111100",
10054 => "110100101100111010001100",
10055 => "110101011001011000001101",
10056 => "110101000101011101011000",
10057 => "110011110000001100011100",
10058 => "110001001000010001011100",
10059 => "101101010111100001011100",
10060 => "101000110011001110011010",
10061 => "100100011111011110100111",
10062 => "100010000011000011010011",
10063 => "100001100110101001010100",
10064 => "100010100111101001001011",
10065 => "100101010100100101101101",
10066 => "101001011000100010101100",
10067 => "101110000010000110000110",
10068 => "110011001100110110110010",
10069 => "111000100001111000110100",
10070 => "111101010011101111111110",
10071 => "000001111000001010001101",
10072 => "000110011101101111110100",
10073 => "001001010101011010010110",
10074 => "001001000111011000011000",
10075 => "000111100001100000101100",
10076 => "000110101000101100010101",
10077 => "000110000010010110100001",
10078 => "000100111101111100001010",
10079 => "000100000000001111010010",
10080 => "000011111000111000000100",
10081 => "000100110011010100001101",
10082 => "000101111110111001000100",
10083 => "000110000100100000111100",
10084 => "000100100101001011010101",
10085 => "000010001110000001100010",
10086 => "111111111011101010001000",
10087 => "111101111101010001100011",
10088 => "111011110111000010101110",
10089 => "111001111101010101010010",
10090 => "111001001100011010111001",
10091 => "111001100111001011010000",
10092 => "111010110110100010000111",
10093 => "111100010111101110000011",
10094 => "111100111100000110110100",
10095 => "111100100010001111110000",
10096 => "111100110000101011010100",
10097 => "111110001111110110000010",
10098 => "000000001101001001100101",
10099 => "000001011100110111111000",
10100 => "000001000010111000011101",
10101 => "111111011100111100000001",
10102 => "111101101111100100010100",
10103 => "111011111101000011010101",
10104 => "111010000011110111011111",
10105 => "111000011100010000101000",
10106 => "110111000011010111011100",
10107 => "110110000110000110111010",
10108 => "110110000011100011001110",
10109 => "110110101011101100000001",
10110 => "110111010101100110011011",
10111 => "110111101001000001110111",
10112 => "110111110101111101000000",
10113 => "111000101111101111010000",
10114 => "111010011011101001001110",
10115 => "111100001101111110101011",
10116 => "111110000111100010001011",
10117 => "000000100111101011001101",
10118 => "000011111011101110110000",
10119 => "001000001100110111110001",
10120 => "001101000010110000110000",
10121 => "010001010111110101001110",
10122 => "010100101110011011110100",
10123 => "010111011010000111100100",
10124 => "011001001010001101111010",
10125 => "011001101010010100110111",
10126 => "011001011101000101101001",
10127 => "011000010010001110101100",
10128 => "010101000101101101010010",
10129 => "010000110111011010101110",
10130 => "001101100110110011010100",
10131 => "001010111001110010000001",
10132 => "000111010100011010110110",
10133 => "000010111110001011100100",
10134 => "111110110010100001000000",
10135 => "111011010000111010000000",
10136 => "111000100001101110001110",
10137 => "110110110101010101110100",
10138 => "110110000110110010011011",
10139 => "110101011001101010110001",
10140 => "110100000101000100111001",
10141 => "110010011100111101111110",
10142 => "110001100111110010111000",
10143 => "110011011001010011111000",
10144 => "110111011110011111000001",
10145 => "111010110100100110100100",
10146 => "111100010000110011010010",
10147 => "111100101001000111000100",
10148 => "111100011110011010101110",
10149 => "111101111011111000011010",
10150 => "000010100110100100000101",
10151 => "000111111000101110000000",
10152 => "001011101010111101001101",
10153 => "001110101001000101101100",
10154 => "010000100100001111000000",
10155 => "010000001001101101100010",
10156 => "001100101011111110010010",
10157 => "000110111101010011100110",
10158 => "000010011101111000001001",
10159 => "000010101101001100110011",
10160 => "000110101100011000101111",
10161 => "001001101110111011001010",
10162 => "001001001000001000000101",
10163 => "000111111000110011110110",
10164 => "001010001000000101110101",
10165 => "001110111000010111110110",
10166 => "010010101101001010010000",
10167 => "010100011010111011101010",
10168 => "010100001100001111001100",
10169 => "010001111011011001100110",
10170 => "001101111001011001000100",
10171 => "001000011011011000000000",
10172 => "000000101001010001100110",
10173 => "110110011001011101000000",
10174 => "101101110100111000110110",
10175 => "101011100000011100010000",
10176 => "101101111011010100101100",
10177 => "110001000000111000010000",
10178 => "110011101001100010100100",
10179 => "110101101000111110101010",
10180 => "110110101101101000101110",
10181 => "110111011111110001110000",
10182 => "110111100101000111111101",
10183 => "110110010111111000110000",
10184 => "110101101111011000101100",
10185 => "110111001010110111010000",
10186 => "111001001011100000010010",
10187 => "111010000001001001001110",
10188 => "111001001100100001110111",
10189 => "110110101111011001001001",
10190 => "110100000001101010010010",
10191 => "110010110001001101101100",
10192 => "110010001101111001011010",
10193 => "110000101111110000110110",
10194 => "101110010111011001011100",
10195 => "101011010111010110001100",
10196 => "100111111100100001010000",
10197 => "100101001010010010001011",
10198 => "100100000011110111100011",
10199 => "100101100000110010011111",
10200 => "101010001010100011001010",
10201 => "110001100000001010111010",
10202 => "111010010100011001111000",
10203 => "000010111011101110010101",
10204 => "001001001110110111001110",
10205 => "001100110101000010111110",
10206 => "001111001101111011010000",
10207 => "010001000101100010001010",
10208 => "010010000011100001000000",
10209 => "010010000100100110000100",
10210 => "010001000001001110111010",
10211 => "001110001010111110101100",
10212 => "001001011101100101101011",
10213 => "000100010001110111000110",
10214 => "111111101011110001100010",
10215 => "111011101100001001011000",
10216 => "111001001011001100111010",
10217 => "111001101001100001111011",
10218 => "111101000110100001110101",
10219 => "000010000100000000100110",
10220 => "000110111011110101100000",
10221 => "001011001111001001100100",
10222 => "001111100110111001111010",
10223 => "010011100111000100000000",
10224 => "010101011100001001111110",
10225 => "010100100010111101100000",
10226 => "010010000110000001101100",
10227 => "001111010011000010000100",
10228 => "001100011001100111100100",
10229 => "001000101001100110101000",
10230 => "000011111001011100000001",
10231 => "111111010011011011100011",
10232 => "111011001110100010000111",
10233 => "110111001010110101010011",
10234 => "110011110011111010011110",
10235 => "110001111000010011100110",
10236 => "110000110010011110101110",
10237 => "110000001011011101100110",
10238 => "110000010010000001010000",
10239 => "110000111000111010000000",
10240 => "110001011101001111110000",
10241 => "110001100001011011001000",
10242 => "110001010111010101001110",
10243 => "110001100111101010111110",
10244 => "110001101000011001110000",
10245 => "110000110001001101011110",
10246 => "110000011100110011011100",
10247 => "110001111100010000001100",
10248 => "110100101111001110010010",
10249 => "111000001011001100100010",
10250 => "111011110100000110010011",
10251 => "111110110011000111111001",
10252 => "000000011111000000111011",
10253 => "000001010000101011001001",
10254 => "000001111011110100101101",
10255 => "000010010110100111010011",
10256 => "000010000101111101111010",
10257 => "000001110001001001001010",
10258 => "000001101111010111110001",
10259 => "000001100000100100011100",
10260 => "000000110001000110001010",
10261 => "111111011100010011100001",
10262 => "111110001100010110011011",
10263 => "111101111100100111001111",
10264 => "111101101101110000101111",
10265 => "111100011001100110101110",
10266 => "111011100100111010011011",
10267 => "111100100111011010001111",
10268 => "111110001111011110001010",
10269 => "111111010101001110100010",
10270 => "000000110110011101011010",
10271 => "000011100100100101001010",
10272 => "000110011011001000010000",
10273 => "001000100000101000110001",
10274 => "001010000110101111100100",
10275 => "001010101101100111110011",
10276 => "001000111010101000100101",
10277 => "000100100000101010001101",
10278 => "111111110011011100011100",
10279 => "111110000101010000001001",
10280 => "111111011111110011000111",
10281 => "000001011100010011011000",
10282 => "000011110110000000110001",
10283 => "001000001101010101001100",
10284 => "001100110000010110011000",
10285 => "001110101000110100100010",
10286 => "001110101011000111001010",
10287 => "010000011011111111010110",
10288 => "010101101011000111000100",
10289 => "011011100001110001000011",
10290 => "011101110101000011111100",
10291 => "011100101001010110101001",
10292 => "011011001011000110110001",
10293 => "011010011010011100010001",
10294 => "011001011000011111100001",
10295 => "011000011000111000101111",
10296 => "010111110011011111110000",
10297 => "010111000111011010111000",
10298 => "010110110100010111111110",
10299 => "010101111000101110100110",
10300 => "010000101110011000111110",
10301 => "000111101111111011111110",
10302 => "111111110000110111011101",
10303 => "111011010001010100010001",
10304 => "111001110101000001000010",
10305 => "111001011101101010100100",
10306 => "110111101111010110000000",
10307 => "110101100110011100100100",
10308 => "110101001100010010110101",
10309 => "110100110110001011011010",
10310 => "110010101100101100010110",
10311 => "110000011010101110101100",
10312 => "110000001010100010110110",
10313 => "110010010011100000001010",
10314 => "110101111000010111111111",
10315 => "111001000110000101101111",
10316 => "111010101101111011011100",
10317 => "111011110011101101100010",
10318 => "111101100100111110110101",
10319 => "111110010000100010001001",
10320 => "111100101101011111001101",
10321 => "111011001000110010000111",
10322 => "111001101000001000000110",
10323 => "110101101111111101011111",
10324 => "101111110111111101110110",
10325 => "101001110101111011011010",
10326 => "100101001100001000111101",
10327 => "100011011111110100100011",
10328 => "100011110111110011101011",
10329 => "100101010101011011111001",
10330 => "101001001100110111101110",
10331 => "101101110111011001110110",
10332 => "110000010110010011000100",
10333 => "110010000010100011110100",
10334 => "110100011000111100001000",
10335 => "110110000010110011100000",
10336 => "110111010100001111000001",
10337 => "111010000101111101011011",
10338 => "111110100111110100001011",
10339 => "000011110010111110000000",
10340 => "001000011000110000100010",
10341 => "001011011010000001011110",
10342 => "001100011100000111110010",
10343 => "001011111010100010101001",
10344 => "001010111100010110010011",
10345 => "001010111000101010110010",
10346 => "001100011011001110000110",
10347 => "001110000110110010101100",
10348 => "001101110110001000100000",
10349 => "001100011101010100110010",
10350 => "001100001111100000001100",
10351 => "001101011111100001011100",
10352 => "001111000111111001101110",
10353 => "010000011101111011000010",
10354 => "010010011110001010011010",
10355 => "010110100011111111101100",
10356 => "011010110010100000100111",
10357 => "011100001011110110011001",
10358 => "011011101110101010101110",
10359 => "011010100000000101110010",
10360 => "010111000111000010010010",
10361 => "010001111011011000111100",
10362 => "001100001101110101001110",
10363 => "000101011000010000011010",
10364 => "111101101000111011110111",
10365 => "110110101100001111100100",
10366 => "110001010001111100011000",
10367 => "101101001101011001001000",
10368 => "101001111110100010011000",
10369 => "100111010011101100010001",
10370 => "100110011100111101000111",
10371 => "101000110100001011010010",
10372 => "101101001111000100000100",
10373 => "110001010011000100011110",
10374 => "110100011000101011010101",
10375 => "110111011110000100101011",
10376 => "111010111100101010010111",
10377 => "111101111000000110101111",
10378 => "111110100111000000100011",
10379 => "111100000001001010010011",
10380 => "110111000111101101101111",
10381 => "110010101011000101010110",
10382 => "110000011000100011111110",
10383 => "101111110000100000100110",
10384 => "101111011101101001100110",
10385 => "101111001010100101110000",
10386 => "101111111101101111101110",
10387 => "110010100010000011011000",
10388 => "110110000110100110111011",
10389 => "111001110111100010010011",
10390 => "111101111000000000101011",
10391 => "000010001001000101111010",
10392 => "000101100100111010111110",
10393 => "000111001110000101111110",
10394 => "000111101001110001001010",
10395 => "000111100111011110000101",
10396 => "000111010100000001001100",
10397 => "000110111010111001000010",
10398 => "000110011010001011110000",
10399 => "000110001111101100011110",
10400 => "000111000110110000100011",
10401 => "001000011101010001101010",
10402 => "001001011000100111010010",
10403 => "001001011010111110101010",
10404 => "001000001110100010111011",
10405 => "000110011111110101001100",
10406 => "000101110000111101000100",
10407 => "000110001010110001010001",
10408 => "000110011110001000000110",
10409 => "000110000101000101101001",
10410 => "000101100010010100101011",
10411 => "000101101010001010001101",
10412 => "000101111010010110010101",
10413 => "000011110000111101101010",
10414 => "111101101100100001001100",
10415 => "110110010000000111100101",
10416 => "110001110011011000100010",
10417 => "110001010000011010000100",
10418 => "110010010100000100000110",
10419 => "110100011011010011111110",
10420 => "110111101101000000000110",
10421 => "111010100001000111111000",
10422 => "111101001011011110011010",
10423 => "000001001011010000011100",
10424 => "000101011010110000011100",
10425 => "001000011100100000001000",
10426 => "001001101011111000101011",
10427 => "001000110111111011111010",
10428 => "000110111110011101000001",
10429 => "000100110010100000101001",
10430 => "000001111110001010010110",
10431 => "111110011000011101010111",
10432 => "111011000110000101010110",
10433 => "111010110100110011000100",
10434 => "111111000000000110000110",
10435 => "000100110101100000000000",
10436 => "001001001011010000110000",
10437 => "001011111010100100100111",
10438 => "001101101111101000000110",
10439 => "001111010110011100000010",
10440 => "010001011111010011011000",
10441 => "010011000111110111101000",
10442 => "010010111100111111111000",
10443 => "010001100011001111101100",
10444 => "001111110111000000011000",
10445 => "001110100101101000101100",
10446 => "001101011111010101101000",
10447 => "001010111010000111000000",
10448 => "000110111110101101011011",
10449 => "000011101110000000111111",
10450 => "000001011101010110011101",
10451 => "111111001101110110011011",
10452 => "111100111101000000110111",
10453 => "111011100000101101010101",
10454 => "111010111100111011110010",
10455 => "111010011000111110010011",
10456 => "111001111100010101101011",
10457 => "111010100100010000001101",
10458 => "111100000110110110111111",
10459 => "111101001111001100110001",
10460 => "111100101000111110100100",
10461 => "111001110101111111010101",
10462 => "110101010011101110011110",
10463 => "110000010011010101110000",
10464 => "101100001110101010000000",
10465 => "101001100100100100011100",
10466 => "101000001110110010000010",
10467 => "101000010110110010011010",
10468 => "101010010000011101011000",
10469 => "101101000001111101000010",
10470 => "101110011100100101011110",
10471 => "101110100100010111100110",
10472 => "101111011111110010001000",
10473 => "110001010100101000100000",
10474 => "110011110101100000101010",
10475 => "110111110101101101101000",
10476 => "111100010111000101001100",
10477 => "111111110111100100101001",
10478 => "000010100001110101000010",
10479 => "000101000100100101000110",
10480 => "000111011010101101011000",
10481 => "001000111101000000111010",
10482 => "001010010010110001111011",
10483 => "001100111100011110000000",
10484 => "010000001010101100001000",
10485 => "010001011101001011001110",
10486 => "010000100101000111010100",
10487 => "001111001100011110110110",
10488 => "001101101101110101110110",
10489 => "001100010111100111001110",
10490 => "001100000101100111100110",
10491 => "001100011111000010010100",
10492 => "001100001001000110001110",
10493 => "001010100110000001001011",
10494 => "001000100101111101011110",
10495 => "000110010100111000011011",
10496 => "000011001100110010010000",
10497 => "000000000110110000001110",
10498 => "111101111110000100001010",
10499 => "111100001110000001011101",
10500 => "111010110100101000001000",
10501 => "111001001011000011100101",
10502 => "110110001010110111101110",
10503 => "110010111001101100001000",
10504 => "110000111010101000101100",
10505 => "110000100111011101000000",
10506 => "110001100001111010100110",
10507 => "110010100010001111000110",
10508 => "110011011011000101111100",
10509 => "110100101000000011000011",
10510 => "110110001100000100001010",
10511 => "111000000010110101110001",
10512 => "111001100101010101111010",
10513 => "111001111001100000110110",
10514 => "111000100111001010010000",
10515 => "110110010001011101110010",
10516 => "110011101101100111111000",
10517 => "110000100110101001111000",
10518 => "101100110010100110001110",
10519 => "101001100011010011000010",
10520 => "100111101000101011111111",
10521 => "100111001000100000100110",
10522 => "101000100101010111111100",
10523 => "101011111011101111110110",
10524 => "110001001000110000100110",
10525 => "111000111110110111110111",
10526 => "000010100011011011001100",
10527 => "001100010110100100110100",
10528 => "010110001110101010010110",
10529 => "011101010000000101010111",
10530 => "011110101011000001110111",
10531 => "011101111111000001110111",
10532 => "011110001111011101001101",
10533 => "011110011010000001010100",
10534 => "011101100010110011010100",
10535 => "011010110110111001001110",
10536 => "010111011010011011101110",
10537 => "010101101000111000101100",
10538 => "010100110110100011110010",
10539 => "010100010000011011111000",
10540 => "010100111111000111010010",
10541 => "010110011110100101011010",
10542 => "010111000110000101111100",
10543 => "010110111110100100010100",
10544 => "010111011101011000011100",
10545 => "011000001110100111010011",
10546 => "010111101001111001110110",
10547 => "010101100111101100011010",
10548 => "010010011110011100110100",
10549 => "001110010000101101110000",
10550 => "001010000101001000010110",
10551 => "000110000000100011111010",
10552 => "000000010100010101010101",
10553 => "111000110111111110001100",
10554 => "110001100111011011010010",
10555 => "101100001010000111011110",
10556 => "101000101101111001100010",
10557 => "100101111000010000111111",
10558 => "100010101111000010010001",
10559 => "100000110111010000000101",
10560 => "100000111111100111101101",
10561 => "100001111001110101011111",
10562 => "100011000100001100110001",
10563 => "100011111011110001001011",
10564 => "100101000001001110100101",
10565 => "101000000101110001000010",
10566 => "101100011110011101100100",
10567 => "110001000111000110111100",
10568 => "110101100111001111110110",
10569 => "111000000011011101101001",
10570 => "111000100001000010110011",
10571 => "111001101101010010001011",
10572 => "111100111001011011101101",
10573 => "000000110001110111100101",
10574 => "000010011100111000111100",
10575 => "000001001101011010100101",
10576 => "111111100101010001111111",
10577 => "111111001011010010010100",
10578 => "111111010000010011100001",
10579 => "111110010001010100110010",
10580 => "111100001011010000000000",
10581 => "111010110011001010000010",
10582 => "111011000000010000101000",
10583 => "111100011100011100100011",
10584 => "111110100101100010110000",
10585 => "000000010011110001001110",
10586 => "000001101101101110000111",
10587 => "000101001011000111001011",
10588 => "001011110001011101010000",
10589 => "010010111110011011010000",
10590 => "010111111101001010101110",
10591 => "011010100001001111010011",
10592 => "011011101110100011101011",
10593 => "011011110011101111011100",
10594 => "011001110110101110000111",
10595 => "010110001110010111000010",
10596 => "010011001101010100000000",
10597 => "010010000111000101011000",
10598 => "010010000010110010111110",
10599 => "010000001110001011111010",
10600 => "001011001001001101110011",
10601 => "000101010001111101000100",
10602 => "000000010101001001111101",
10603 => "111100011000010110010011",
10604 => "111011000001110000011100",
10605 => "111100000110010101011100",
10606 => "111101101001001110100111",
10607 => "111111001101010101100101",
10608 => "000000110001100000011010",
10609 => "000001111101000010000010",
10610 => "000010010101001101101011",
10611 => "000010100111000110010000",
10612 => "000100000100010001001000",
10613 => "000101100100001011101100",
10614 => "000101000110011111111010",
10615 => "000010011111011110001101",
10616 => "111110110000011010101010",
10617 => "111011001100001001011111",
10618 => "111000011000111000011111",
10619 => "110110011101000010010011",
10620 => "110101101100010110000100",
10621 => "110110010000110100010000",
10622 => "110111110110011110000001",
10623 => "111001101000001001101010",
10624 => "111011001101100000000101",
10625 => "111100111110000100111111",
10626 => "111110111010010110000000",
10627 => "000000011110101101001001",
10628 => "000001010010110000100111",
10629 => "000001101000101101000110",
10630 => "000001000000001100001010",
10631 => "111110000100011010111100",
10632 => "111001010111011101010101",
10633 => "110100011101110000100110",
10634 => "110000100101000000110000",
10635 => "101110101010000000011100",
10636 => "101101111000101000001100",
10637 => "101100100001110101000110",
10638 => "101010001011000000011010",
10639 => "101000100100110001110100",
10640 => "101001101111101000101000",
10641 => "101100000100100001010000",
10642 => "101101000111000111001100",
10643 => "101101001101111001110000",
10644 => "101101000011010110100000",
10645 => "101101010111101010110000",
10646 => "101110100110111000010010",
10647 => "101111100100111111001110",
10648 => "101111111111010101011010",
10649 => "110000110100011010001100",
10650 => "110010101001111111000110",
10651 => "110100111010001001110110",
10652 => "110110000011100001110110",
10653 => "110110010101110111000111",
10654 => "110111101000001001110100",
10655 => "111010001111110111010100",
10656 => "111100111110101100000110",
10657 => "111111011100010011100000",
10658 => "000010100001001010010001",
10659 => "000110001000110011001101",
10660 => "001001100010011110111001",
10661 => "001100110100011100110100",
10662 => "001111110001011111000010",
10663 => "010010000111111001110110",
10664 => "010100111100010111011110",
10665 => "011001011010010010010001",
10666 => "011101110001100010011110",
10667 => "011110101011111011011111",
10668 => "011101001110100101100101",
10669 => "011100011111101111001101",
10670 => "011100000000111111001001",
10671 => "011011010101011011110001",
10672 => "011010101010111111100111",
10673 => "011001000110110000111101",
10674 => "010111110100100110110100",
10675 => "011000000011111101111111",
10676 => "011000010111101010110111",
10677 => "011000001000111110100111",
10678 => "010111110100010000111000",
10679 => "010111000111010000000110",
10680 => "010110101001011011110000",
10681 => "010110110001001001011000",
10682 => "010110010111001100101010",
10683 => "010110010111110010111100",
10684 => "010110001000011101110100",
10685 => "010000010010011010111000",
10686 => "000101001000100110000001",
10687 => "111001001010010000001001",
10688 => "101100011000001110010110",
10689 => "100010101001000001000001",
10690 => "100000111001101100101011",
10691 => "100001111011000110010010",
10692 => "100001001111010001001100",
10693 => "100001100001100000001111",
10694 => "100010111101010100111101",
10695 => "100011011111011010111111",
10696 => "100100010100000110111001",
10697 => "100111101110011101110011",
10698 => "101101000111000111100010",
10699 => "110010010100001111011100",
10700 => "110110111001000101101011",
10701 => "111010100001011001110000",
10702 => "111011111010111111111010",
10703 => "111011101100000110110001",
10704 => "111011100111011110111011",
10705 => "111010100110110100111000",
10706 => "110110110001111110011100",
10707 => "110010010001101011101110",
10708 => "101111110000101000010100",
10709 => "101110101001011110110110",
10710 => "101101111010011001111110",
10711 => "101101010101011111101000",
10712 => "101100101111011000000100",
10713 => "101100001000101111111110",
10714 => "101100100110000111001100",
10715 => "101111011010110011100000",
10716 => "110011101001101100110000",
10717 => "111000010001001101111111",
10718 => "111100110111011111101011",
10719 => "111111110101001000110001",
10720 => "000010001010101001100110",
10721 => "000101100010000100111100",
10722 => "000111100111000101001011",
10723 => "000111001111000111011000",
10724 => "000110100101111000011111",
10725 => "001000000000010100011101",
10726 => "001011010000101010101001",
10727 => "001101000100110001010000",
10728 => "001100011000011001101100",
10729 => "001010110111101100101011",
10730 => "001000010001010111000000",
10731 => "000100000101011011111000",
10732 => "111111110111110010110111",
10733 => "111101100101110000011001",
10734 => "111101100101101100011110",
10735 => "111110101001101011101011",
10736 => "000000010001100111010001",
10737 => "000010011011110101011110",
10738 => "000100010000111101101000",
10739 => "000101010001000101111111",
10740 => "000110010101110001111100",
10741 => "001000111010110101101101",
10742 => "001100111000111010101010",
10743 => "010000001010100110110110",
10744 => "010000110111101100110000",
10745 => "001111101111111100001010",
10746 => "001110110010011111011110",
10747 => "001101011100110101001010",
10748 => "001011001010111110001010",
10749 => "001001111000011101111000",
10750 => "001010000010101001101100",
10751 => "001010100100101010010000",
10752 => "001011000001010001111000",
10753 => "001011000111001101000010",
10754 => "001010101101010100001110",
10755 => "001001001100001110001000",
10756 => "000110111010100100100110",
10757 => "000101010100010001001101",
10758 => "000100100011001011000111",
10759 => "000100011001101000101001",
10760 => "000011101111010110111000",
10761 => "000001100100101001111001",
10762 => "000000000010101000101110",
10763 => "000000101001000010010011",
10764 => "000010100101001000111001",
10765 => "000100011110110010010111",
10766 => "000100001010111111101000",
10767 => "000001011111011000001101",
10768 => "111101110000101001001001",
10769 => "111000110101101001011010",
10770 => "110011010001111111101000",
10771 => "101110010100011001100010",
10772 => "101001110010011100010010",
10773 => "100101111100110010111001",
10774 => "100100100110110110010001",
10775 => "100101110100000100011110",
10776 => "100110111101100001010111",
10777 => "100111011101000111000011",
10778 => "101001010010100001001010",
10779 => "101101000010001001101000",
10780 => "110000111111100010010110",
10781 => "110011001111111010000100",
10782 => "110100001111100101000000",
10783 => "110101011010101010000011",
10784 => "110110011100100111100111",
10785 => "110110111101110000100011",
10786 => "110111100011010001111110",
10787 => "111001000011001111100001",
10788 => "111011001111101110000111",
10789 => "111100011001001001011000",
10790 => "111100011010001100010111",
10791 => "111100010000000110110000",
10792 => "111100001011011011111011",
10793 => "111101011111110011000100",
10794 => "000000011101010111100010",
10795 => "000011111100001000011100",
10796 => "001000000010011100000100",
10797 => "001100110101000011010110",
10798 => "010001110110111010000000",
10799 => "010110010110101100110110",
10800 => "011001011010011010110010",
10801 => "011011010000001000100011",
10802 => "011100100100101100110101",
10803 => "011101011001110010001111",
10804 => "011101000010011111010101",
10805 => "011011110101100111100111",
10806 => "011011000110110111000101",
10807 => "011010011011001110101001",
10808 => "011001011110111000001000",
10809 => "011000110000111111101000",
10810 => "010111111101010111101110",
10811 => "010111100100010000010010",
10812 => "010111011100010100011110",
10813 => "010110111110110001010100",
10814 => "010111000000010011100110",
10815 => "010101110011101011000010",
10816 => "010001010010011010011000",
10817 => "001011110000100110110011",
10818 => "000111000100110011001100",
10819 => "000010010011111001111000",
10820 => "111101110000101111101011",
10821 => "111010000001100001001011",
10822 => "110101100111101010110001",
10823 => "110000101100110100101110",
10824 => "101101110011101001101000",
10825 => "101100100010001101110100",
10826 => "101010000001011000011110",
10827 => "100101100001010101101011",
10828 => "100001110010110011111010",
10829 => "100001100001110110010011",
10830 => "100010010010001010001001",
10831 => "100010101001111001011111",
10832 => "100110110111100100111001",
10833 => "101110110100101000001110",
10834 => "110101011101000110100110",
10835 => "111000111101011110101100",
10836 => "111010000000101000001001",
10837 => "111001110010101011101000",
10838 => "111001001001010000001100",
10839 => "110111001001011101011110",
10840 => "110011010101100010111000",
10841 => "101111100100001010001100",
10842 => "101101110101110111011100",
10843 => "101101011110111110001000",
10844 => "101101001111001011100010",
10845 => "101110000100010101111000",
10846 => "110001101000111110101010",
10847 => "111000101100100011110101",
10848 => "000001100011100101010101",
10849 => "001001011010000010001111",
10850 => "001111001111001010111100",
10851 => "010010011111101100000000",
10852 => "010011011000101011010010",
10853 => "010011000101101001000110",
10854 => "010001100111001010000010",
10855 => "001111011111110100001000",
10856 => "001101100100000110111010",
10857 => "001011010010001100111101",
10858 => "001000010100101001111110",
10859 => "000100100111110101110111",
10860 => "000000100100001001011101",
10861 => "111100111101100101111111",
10862 => "111010101111011110100010",
10863 => "111011000111100111110110",
10864 => "111101001101001011111111",
10865 => "111110111100000101111011",
10866 => "000000010110101111001000",
10867 => "000001110111010100111011",
10868 => "000010011111100000001000",
10869 => "000001100001010011101000",
10870 => "000000000110111001100110",
10871 => "111111011001101001111010",
10872 => "111110101111110001111001",
10873 => "111101111001010001101010",
10874 => "111100111011001011011101",
10875 => "111011010010011000010100",
10876 => "111000111001011110011110",
10877 => "110110001001110111100000",
10878 => "110100100111100010100100",
10879 => "110101001101100110110101",
10880 => "110110010100000110110000",
10881 => "110110110000001001001011",
10882 => "110110010111010111100000",
10883 => "110101001101010001011010",
10884 => "110100000010011110001010",
10885 => "110011011100000110010100",
10886 => "110011110101001011110010",
10887 => "110100110110100011111100",
10888 => "110101111111101110110110",
10889 => "110111110110000010100100",
10890 => "111010010100101000110110",
10891 => "111101100010101001110000",
10892 => "000001100001101000000100",
10893 => "000100101100000010101001",
10894 => "000111001101110000111111",
10895 => "001010100000110001101111",
10896 => "001101111001100111110000",
10897 => "001111110101100011100010",
10898 => "001111110110101000110110",
10899 => "001111000101011111101000",
10900 => "001110010101000110101100",
10901 => "001101011011001101001010",
10902 => "001100100110101100111000",
10903 => "001011100011101001110110",
10904 => "001010010101111101011000",
10905 => "001001111000100100000110",
10906 => "001010000000110010010110",
10907 => "001010000001111111101010",
10908 => "001001001111010011111001",
10909 => "000111000111111111011011",
10910 => "000011110111110100010011",
10911 => "000000010001100111001000",
10912 => "111101111001001101101110",
10913 => "111101010111010001000001",
10914 => "111101110100001100001110",
10915 => "111110101111111001011110",
10916 => "000000100011010010101100",
10917 => "000011011010000001100100",
10918 => "000100111110110010110101",
10919 => "000010001001001110111010",
10920 => "111011011100111101010111",
10921 => "110100001100010010111101",
10922 => "101110110101010000101110",
10923 => "101011011010011100101000",
10924 => "101001111011010000001000",
10925 => "101011110011110011100000",
10926 => "101111111101100010100010",
10927 => "110100001010010011010100",
10928 => "111000100001000001010010",
10929 => "111101000010100011100010",
10930 => "000010000100010001001111",
10931 => "000111110110000101110000",
10932 => "001101100000010111001000",
10933 => "010011101011100101100110",
10934 => "011001101110101010011101",
10935 => "011100101110111101100111",
10936 => "011100011101000111101101",
10937 => "011011000011110100010101",
10938 => "011010000101110111101001",
10939 => "011001011110000111011010",
10940 => "011000110101101010100111",
10941 => "011000011111000001001001",
10942 => "010111011010110010110110",
10943 => "010100001101001100011100",
10944 => "001110110101001001000000",
10945 => "001000100001001000001100",
10946 => "000011001111011011110100",
10947 => "111111100001110100100011",
10948 => "111100010010110100111101",
10949 => "111001101100110011011010",
10950 => "111001011101111000010101",
10951 => "111011100011010000001110",
10952 => "111101101000101001100011",
10953 => "111111011111111111101110",
10954 => "000010000101011110001110",
10955 => "000100100000011111110000",
10956 => "000111000101000010011101",
10957 => "001010101100100111111111",
10958 => "001101011110000010111100",
10959 => "001100110001100100101010",
10960 => "001001001111111101010110",
10961 => "000101101010011100110000",
10962 => "000001100111110010010111",
10963 => "111011011001100110010100",
10964 => "110011001110001001011010",
10965 => "101001100010101101000010",
10966 => "100010010100011010111111",
10967 => "100001001101111011001101",
10968 => "100001110110111000101011",
10969 => "100001001011100001101110",
10970 => "100001100110111010010011",
10971 => "100010110001011101010101",
10972 => "100011101000110010000011",
10973 => "100100110000100011100001",
10974 => "100101010110011010010011",
10975 => "100110010111100111000011",
10976 => "101010010111010001000110",
10977 => "101111100110111000011010",
10978 => "110010011000011010000100",
10979 => "110011111011111000001110",
10980 => "110111000011000100110100",
10981 => "111010100011010111110110",
10982 => "111101101001000101110010",
10983 => "000001011010010010110001",
10984 => "000110001111011001001010",
10985 => "001100110001110010111110",
10986 => "010100100011000001000110",
10987 => "011010011111110001010010",
10988 => "011011111101001000001000",
10989 => "011001110011100100010000",
10990 => "010111000111111101111100",
10991 => "010100000111011101110100",
10992 => "001111010111010111101110",
10993 => "001001110010101101110101",
10994 => "000100111001001111100101",
10995 => "000001011011110000001011",
10996 => "111111100001011011110110",
10997 => "111110101010000000111110",
10998 => "111110001011001010010110",
10999 => "111110010100100001010100",
11000 => "000001000011000010101111",
11001 => "000110011010011101111011",
11002 => "001100100101011100110110",
11003 => "010010110110101000100010",
11004 => "010111010110100001111000",
11005 => "011000100000001100000011",
11006 => "010110110001001100000110",
11007 => "010010111010100011101000",
11008 => "001110100001010111001110",
11009 => "001001110110111011100000",
11010 => "000100101011000101010001",
11011 => "111111111100100010010101",
11012 => "111010100100101111011001",
11013 => "110100000101000010100100",
11014 => "101110101001011001000010",
11015 => "101011000000111000110110",
11016 => "101000010110011110010110",
11017 => "100110010110000110110000",
11018 => "100101101011101010001001",
11019 => "100101110001001011010001",
11020 => "100100101001000000000101",
11021 => "100011011101100101100011",
11022 => "100100000011110100100110",
11023 => "100100110010100001101011",
11024 => "100101001101100110111011",
11025 => "100111011011010100110010",
11026 => "101011000111000001111110",
11027 => "101110011101000010110100",
11028 => "110001101110100111000110",
11029 => "110101011101001011000101",
11030 => "111000101001000000000010",
11031 => "111010010101010111111001",
11032 => "111010111101001110100100",
11033 => "111011110011001001110000",
11034 => "111101010000110101011110",
11035 => "111110011010011111110000",
11036 => "111110010111010000110100",
11037 => "111101010100001110110000",
11038 => "111100011100011010100100",
11039 => "111100111000100011110111",
11040 => "111110100001110001000100",
11041 => "000000001100010010000001",
11042 => "000010010000010111101100",
11043 => "000110010111000001111010",
11044 => "001011100111001111000111",
11045 => "001111100111110000010110",
11046 => "010001011100011111010010",
11047 => "010001101011110010010000",
11048 => "010001010110100111111100",
11049 => "010000010011011111110010",
11050 => "001110010011110000101110",
11051 => "001100010111100111000100",
11052 => "001011101100001111110100",
11053 => "001100111000000100111100",
11054 => "001110110100111000001110",
11055 => "001111111111100000100100",
11056 => "010000101111101001001000",
11057 => "010001110101001101001100",
11058 => "010010110001100111100010",
11059 => "010011001011100011011100",
11060 => "010011011100010110011100",
11061 => "010011110110110100101010",
11062 => "010100100101011011110010",
11063 => "010101010101010101111100",
11064 => "010101010111110100111110",
11065 => "010101000110101010110000",
11066 => "010100111100101011000000",
11067 => "010101001000100100111000",
11068 => "010110011000010110000000",
11069 => "010111010101011001010010",
11070 => "010110110110010111011000",
11071 => "010110001101110010111010",
11072 => "010100000111111010111000",
11073 => "001101100000000011000010",
11074 => "000100000001111101000010",
11075 => "111011101101100111111110",
11076 => "110101000100000011110000",
11077 => "110000000000100101101010",
11078 => "101101001110101101000000",
11079 => "101011001000110000010000",
11080 => "101001110000110011011100",
11081 => "101011100010101110101100",
11082 => "110000001111100100011110",
11083 => "110110010000001011100011",
11084 => "111101000100111011100000",
11085 => "000100100010010100001110",
11086 => "001011100000010111010110",
11087 => "010000110111011000110000",
11088 => "010100101011101000110000",
11089 => "010100111111011010010110",
11090 => "010000001100100010111110",
11091 => "001001110100100011010101",
11092 => "000100101111011111000100",
11093 => "000000010100111110001001",
11094 => "111100010110100110011000",
11095 => "111000111101101011010001",
11096 => "110101110101010001010100",
11097 => "110001111011001011000110",
11098 => "101100011011011111011100",
11099 => "100111101001110100100101",
11100 => "100110001010100011000110",
11101 => "100101010111010000100011",
11102 => "100010100011001110000011",
11103 => "100001001010011110001000",
11104 => "100010111000010111110011",
11105 => "100100000011101111111001",
11106 => "100100100100111001100001",
11107 => "100101101110111110111011",
11108 => "100101110011110010011001",
11109 => "100110100000001100011100",
11110 => "101010111111001000000100",
11111 => "110001001111001011101110",
11112 => "110110000000000001010001",
11113 => "111001101101001110101011",
11114 => "111101110011011000100100",
11115 => "000001011101100101111000",
11116 => "000100000001111111110001",
11117 => "000101111100100110010111",
11118 => "000111000000000100011001",
11119 => "000111001001100101000010",
11120 => "000101110101111101000110",
11121 => "000011110101111100001011",
11122 => "000011111001100101110110",
11123 => "000101101111110110010111",
11124 => "001000101011111010000111",
11125 => "001100111100110101011100",
11126 => "001111100001001101110110",
11127 => "001110111100100111110010",
11128 => "001101100011101100011110",
11129 => "001100110000101110111100",
11130 => "001011110001000010100110",
11131 => "001000110001110000000110",
11132 => "000100110011100000010110",
11133 => "000010101001101101100001",
11134 => "000010101110111011101000",
11135 => "000100010101001110101111",
11136 => "000101011110110110010100",
11137 => "000101001011011001000101",
11138 => "000101111111001111111000",
11139 => "001000111101110011011110",
11140 => "001100111010111111100110",
11141 => "010000101110001001101000",
11142 => "010010110100000011101110",
11143 => "010010100000000010101110",
11144 => "001111110010011110001100",
11145 => "001011001001011100011001",
11146 => "000100110100110100111011",
11147 => "111101001011010100001011",
11148 => "110110100100011111001110",
11149 => "110010000100001100111100",
11150 => "101110111110011100000110",
11151 => "101100011101011000001000",
11152 => "101001110001101100010110",
11153 => "101000101111011011111110",
11154 => "101001111111001100001000",
11155 => "101100100001101011101100",
11156 => "101111110111010101101010",
11157 => "110001100011100001001110",
11158 => "110001101111001110111000",
11159 => "110001101101001111010000",
11160 => "110000011001100000101110",
11161 => "101110001110011101000000",
11162 => "101011011011001010001100",
11163 => "101001011001100110010100",
11164 => "101001011110111000000000",
11165 => "101010100010011001011100",
11166 => "101101100100010010011110",
11167 => "110001111111000001000110",
11168 => "110101101001001101100101",
11169 => "110111111111110111000111",
11170 => "111000010010100000001111",
11171 => "111000010011111010111001",
11172 => "111001011011111011101011",
11173 => "111011010010111110001110",
11174 => "111101101110100010010001",
11175 => "111111001011001110001011",
11176 => "000000110000000111101000",
11177 => "000011101011001011101110",
11178 => "000101101000000101110100",
11179 => "000101100111001000110101",
11180 => "000100100101111011000101",
11181 => "000100001011001001000011",
11182 => "000100100010110000010100",
11183 => "000100100000000100001100",
11184 => "000100010010011000001101",
11185 => "000100101000010111101110",
11186 => "000101011001000111001000",
11187 => "000101110100100110000000",
11188 => "000110011001100010011001",
11189 => "000111110111101111000010",
11190 => "001001001111000001000101",
11191 => "001001110100111010111100",
11192 => "001010010110111011111000",
11193 => "001011111001110000101011",
11194 => "001101011110010010010100",
11195 => "001110010010111111101010",
11196 => "010000000000101111101010",
11197 => "010010001100011100100010",
11198 => "010100001010100101011010",
11199 => "010101110111000101000110",
11200 => "010110010100111000010000",
11201 => "010110011001101001110110",
11202 => "010101110010101110011100",
11203 => "010010111101111000001110",
11204 => "001101111101111011100100",
11205 => "001000001010010100011010",
11206 => "000011101010001011110100",
11207 => "000000010001110011000100",
11208 => "111101000111100101000110",
11209 => "111010011011110111100001",
11210 => "111000100100000000000101",
11211 => "111000010100100100011100",
11212 => "111001100110111001011010",
11213 => "111011111110010101010100",
11214 => "111111010011001001001000",
11215 => "000100001000101110110001",
11216 => "001001111010010110111100",
11217 => "001110001110010011011010",
11218 => "010010100001011001101010",
11219 => "010110100111110100100010",
11220 => "010111000011010000010000",
11221 => "010101101111100011101100",
11222 => "010100100111011111110100",
11223 => "010010110010001001100010",
11224 => "001111100101101111010010",
11225 => "001011000111110000001100",
11226 => "000110011111111000000010",
11227 => "111111110011011101010000",
11228 => "110110111010111010000011",
11229 => "101111001101110001011000",
11230 => "101001000100011001101110",
11231 => "100100111011111101000101",
11232 => "100011101010000011101001",
11233 => "100100110110001100001000",
11234 => "100111011000100000110011",
11235 => "101001100101111011111010",
11236 => "101100100100110000101110",
11237 => "110001101011000111010110",
11238 => "110111101011110001110111",
11239 => "111100111000010101011000",
11240 => "000000011110111010010111",
11241 => "000001011011010000010010",
11242 => "111101110111101110101011",
11243 => "111000010101010001111111",
11244 => "110100000010111100110101",
11245 => "110000001100001101100100",
11246 => "101101101110010110111110",
11247 => "101110011000101100101110",
11248 => "110000100000111011111110",
11249 => "110000001111000100000000",
11250 => "101101010000010100101100",
11251 => "101011111000010101000100",
11252 => "101101010011100001011100",
11253 => "110000100111101001101110",
11254 => "110100011101010100100001",
11255 => "110111100111010100101111",
11256 => "111100011101010010101001",
11257 => "000010101010000110011110",
11258 => "000111111111001001010111",
11259 => "001100100100011100011100",
11260 => "010000001110000101110110",
11261 => "010100101001101101010110",
11262 => "011010010111111001000111",
11263 => "011110010011001001001001",
11264 => "011110101111101011001111",
11265 => "011101000100111100101111",
11266 => "011100000100100101010101",
11267 => "011011010000100011111001",
11268 => "011000111010100110101011",
11269 => "010101010110001000011010",
11270 => "001111110111001111010010",
11271 => "001001100010001000011000",
11272 => "000101001000011011110011",
11273 => "000010111010101001110011",
11274 => "000001011000010011011000",
11275 => "111111000100010101000111",
11276 => "111101000001001101000001",
11277 => "111101000000011000010111",
11278 => "111110011101011010111011",
11279 => "000000010001110011001101",
11280 => "000001101001010101001100",
11281 => "000001101100001101111010",
11282 => "111111011100011101111011",
11283 => "111011000010010100011001",
11284 => "110110011010001001011111",
11285 => "110010011100001001000000",
11286 => "101110110100001001111010",
11287 => "101100001001110111100110",
11288 => "101011010010100001000010",
11289 => "101100101111011111110000",
11290 => "110000001000011011100110",
11291 => "110011100110001000000100",
11292 => "110110001110000110100010",
11293 => "111000101100011011011100",
11294 => "111010111100101010111001",
11295 => "111100001000111000000110",
11296 => "111011100011100100101010",
11297 => "111001010010000100011101",
11298 => "110101111111100101100110",
11299 => "110010000011000110000010",
11300 => "101110100110110001001100",
11301 => "101100011011010000000100",
11302 => "101011011000110000111110",
11303 => "101100111010000110101010",
11304 => "110001101001101111111000",
11305 => "111000101100010110100000",
11306 => "000000110101100000010011",
11307 => "001000000111011000001010",
11308 => "001110000100011110111100",
11309 => "010010111001101000000010",
11310 => "010110000011110001110000",
11311 => "010111111111010000110010",
11312 => "011000010100001000011101",
11313 => "010110110110000101001110",
11314 => "010101010010111110110010",
11315 => "010100001101011100110110",
11316 => "010011000001011111000010",
11317 => "010001101011001001111010",
11318 => "010000101101010110000000",
11319 => "010000110100000010010100",
11320 => "010001110101110000000010",
11321 => "010010110001111010100010",
11322 => "010001111010111101010100",
11323 => "001111011011110111100010",
11324 => "001101000000111000111000",
11325 => "001001101000100100000100",
11326 => "000100101111001100001001",
11327 => "000000000111000001111011",
11328 => "111100110110000011001101",
11329 => "111011111010111000110000",
11330 => "111100110111111001101000",
11331 => "111101110110001100110000",
11332 => "111101100101100001000000",
11333 => "111011000101010010100100",
11334 => "110111100100010010101111",
11335 => "110100100100101011100000",
11336 => "110001011100111100010010",
11337 => "101110001101110111111100",
11338 => "101011010001010001010000",
11339 => "101001000001011001011110",
11340 => "100111010001000001101001",
11341 => "100100110101011100101110",
11342 => "100010111100101100111111",
11343 => "100010110000011010011101",
11344 => "100011100101010010100011",
11345 => "100110100110110101111100",
11346 => "101100010111000100001110",
11347 => "110010110001010000100010",
11348 => "111000110001000100000110",
11349 => "111110011111000101101100",
11350 => "000011011000101110010111",
11351 => "000111001000100011011000",
11352 => "001010100001110110001000",
11353 => "001101101110000110010000",
11354 => "001111100101100001011000",
11355 => "010000010111100011001110",
11356 => "010001100010111011000000",
11357 => "010010100010010111000000",
11358 => "010001001000110100001110",
11359 => "001101100101110001101010",
11360 => "001011000001011001100110",
11361 => "001010001011111001111000",
11362 => "001001010101100001000100",
11363 => "001001001111011110001110",
11364 => "001010010011110000100100",
11365 => "001011001101100010101010",
11366 => "001100001100100110100010",
11367 => "001101010000101100100000",
11368 => "001110100101100000010000",
11369 => "010000010001101110010110",
11370 => "010010010000011000010000",
11371 => "010101011010001011000010",
11372 => "010111010001001001010000",
11373 => "010110011001010011000010",
11374 => "010011111000011010100010",
11375 => "001110110111001010001010",
11376 => "001001111100100101101000",
11377 => "000110101101010100111111",
11378 => "000010101001101101000010",
11379 => "111010111000100011000000",
11380 => "101101000111101111000010",
11381 => "100010001101011000000001",
11382 => "100001001010111111101111",
11383 => "100001111111000010001000",
11384 => "100010000010111111110000",
11385 => "100011010011101110001101",
11386 => "100011111101111110111110",
11387 => "100100101101101001101011",
11388 => "100101010101010110101111",
11389 => "100111110101100010010101",
11390 => "101111110100110100110110",
11391 => "111010001100101001010100",
11392 => "000010101101110110100100",
11393 => "001001110010011111101110",
11394 => "010001001010110001110010",
11395 => "010110110000001100010110",
11396 => "010111000101111011000000",
11397 => "010010110101111000111110",
11398 => "001101000010110101011000",
11399 => "001001011001111000000001",
11400 => "001001010011100110101110",
11401 => "001001111000011001011010",
11402 => "001000100011101100010101",
11403 => "000101001111010000100010",
11404 => "000001011010001010110010",
11405 => "111111000100111000010110",
11406 => "111110010001110110000110",
11407 => "111100101111011100010000",
11408 => "111001110011001110100010",
11409 => "110111111001111101000111",
11410 => "111001001110000101101100",
11411 => "111100010110100011010100",
11412 => "111101011101011001010001",
11413 => "111100010011011111100001",
11414 => "111011011111100000011001",
11415 => "111100000001101000101011",
11416 => "111110111110000100101100",
11417 => "000011010011001101010010",
11418 => "000110011101111010100011",
11419 => "000111110001010110011000",
11420 => "000110011011000110111101",
11421 => "000011011000010100110100",
11422 => "111111111010101001101011",
11423 => "111011011011110101000001",
11424 => "110110111010011001100001",
11425 => "110100000110000100111000",
11426 => "110011100101000011001110",
11427 => "110011101100010110010110",
11428 => "110010111011101110111110",
11429 => "110001111100111000100010",
11430 => "110000010100111010010100",
11431 => "101111001011011010001110",
11432 => "110000010110010010100010",
11433 => "110010000110011001011100",
11434 => "110010111011011111101110",
11435 => "110010111000000101011010",
11436 => "110001111010111101111000",
11437 => "110000010001000110000110",
11438 => "101111000110010010011000",
11439 => "101111001011010010011010",
11440 => "101111000001011111000000",
11441 => "101111011111100011100010",
11442 => "110011011101111010100010",
11443 => "111010001100101010100001",
11444 => "000001011110111101010000",
11445 => "001000011000010011011000",
11446 => "001110100001100110110000",
11447 => "010100101000011001011100",
11448 => "011010110001000111101001",
11449 => "011110000000111001000011",
11450 => "011101011001001110100001",
11451 => "011100001011100100000001",
11452 => "011011011000001011011000",
11453 => "011010101011110010001011",
11454 => "011010001100000111111101",
11455 => "010111110000000001101110",
11456 => "010011111110110110010010",
11457 => "010001111101101001101000",
11458 => "010001111000000101000000",
11459 => "010010011000111000000100",
11460 => "010010011111110100001100",
11461 => "010001111111011000011110",
11462 => "010000111001001001111000",
11463 => "001111100011000111011000",
11464 => "001101101111101101111000",
11465 => "001001111001000110000011",
11466 => "000100001101010101111111",
11467 => "111101010010010001000111",
11468 => "110101111000010111100001",
11469 => "101111101101000001000000",
11470 => "101000111100100110011000",
11471 => "100010101011011010100101",
11472 => "100001100001100010110011",
11473 => "100010110100101000101111",
11474 => "100011010010010010000111",
11475 => "100011111111011001011101",
11476 => "100101010111110011000011",
11477 => "101000101110001100011110",
11478 => "101100110001110110000100",
11479 => "101111010101010011110110",
11480 => "110010010011110001111110",
11481 => "110100101111101000010101",
11482 => "110100010010110100101001",
11483 => "110010111000000000010010",
11484 => "110010100011100000000010",
11485 => "110010111010100000001010",
11486 => "110010000101000010110010",
11487 => "110000110010101001010010",
11488 => "110001000000110001011010",
11489 => "110001100000000101001000",
11490 => "110001101011010100011010",
11491 => "110010100010101100000010",
11492 => "110100010010101111111100",
11493 => "110110000101100000011001",
11494 => "110111101011010100100101",
11495 => "111010100111111110010001",
11496 => "111110001111011111110001",
11497 => "000001100010101011111001",
11498 => "000101110011110110100111",
11499 => "001010111010010011101110",
11500 => "010000001100110111000000",
11501 => "010101000101100101100010",
11502 => "011001101100001100011101",
11503 => "011101100111100100001010",
11504 => "011110101111001100010011",
11505 => "011110010011010110110011",
11506 => "011101110001100110010111",
11507 => "011100101100101100010011",
11508 => "011100001011100000100000",
11509 => "011100001000000110101011",
11510 => "011010110101110000101100",
11511 => "010110001010010100100000",
11512 => "001111000001010011111010",
11513 => "001000111110000010011010",
11514 => "000100000110100110111110",
11515 => "000000100110110011111110",
11516 => "111110000011000011111101",
11517 => "111001100111001100010010",
11518 => "110100000011110000100010",
11519 => "110000100010011001101010",
11520 => "110001011110001010111110",
11521 => "110101110111100001100110",
11522 => "111010010110101010011110",
11523 => "111110011100100010000101",
11524 => "000010111010000100110011",
11525 => "000111000000110100110010",
11526 => "001000101101111100100001",
11527 => "001000011100001101101010",
11528 => "001001010001101011011110",
11529 => "001011000100110101101001",
11530 => "001100000001001111011000",
11531 => "001011010001000000001100",
11532 => "001000011000001000101010",
11533 => "000011001111111101101011",
11534 => "111100001111010000110111",
11535 => "110101010011110100011001",
11536 => "110000001000101010010100",
11537 => "101110100000110010001100",
11538 => "110000101101101001001010",
11539 => "110010111010011001111110",
11540 => "110100000110110000010100",
11541 => "110110010011100111010001",
11542 => "111001011110000101001010",
11543 => "111100100001100110101010",
11544 => "111111100010111100111101",
11545 => "000011011001000001010111",
11546 => "000110010101101011110001",
11547 => "000111111110111100111010",
11548 => "001010110011000111101010",
11549 => "001101000101101100100010",
11550 => "001011001000101000000000",
11551 => "000101000000100010100000",
11552 => "111111011111011000011100",
11553 => "111110000000011001011000",
11554 => "111110000101111010011101",
11555 => "111110000011111010011011",
11556 => "111110001010010100101000",
11557 => "111101110111011111101101",
11558 => "111100011111100100011010",
11559 => "111001001011010101111100",
11560 => "110100111101001111011001",
11561 => "110001001000100001101110",
11562 => "101110100100111000001100",
11563 => "101110101000010000101000",
11564 => "110000100100111111100000",
11565 => "110011011000001110100100",
11566 => "110110010100010110011011",
11567 => "111000001110000000100000",
11568 => "111001101011101011011100",
11569 => "111100100110011100111000",
11570 => "000000111100010100110111",
11571 => "000100011000011100010101",
11572 => "000110001000111000011011",
11573 => "000110000100011011001010",
11574 => "000011010111110110101011",
11575 => "111111100111111010101001",
11576 => "111100100011100001110000",
11577 => "111011000010111100101100",
11578 => "111011100010101000100001",
11579 => "111101100100011000010100",
11580 => "000010001010101011000010",
11581 => "001001000101010111010010",
11582 => "001111010011110000001010",
11583 => "010011001000011101000000",
11584 => "010101000100011011000010",
11585 => "010110111101110100000000",
11586 => "011001001100001010100011",
11587 => "011001101110100111001001",
11588 => "011000100010010011000001",
11589 => "011000000000000001001001",
11590 => "010111100101111011001010",
11591 => "010100110011011111000110",
11592 => "010000011111101111101010",
11593 => "001100010111101100000010",
11594 => "001001010011101000001011",
11595 => "001000010010010000011011",
11596 => "000111111101000110111111",
11597 => "000110100000110111011100",
11598 => "000011100000110100111111",
11599 => "111111010011010100111001",
11600 => "111010111101110110100111",
11601 => "110110111111110100101011",
11602 => "110011100110000010110110",
11603 => "110000001111000100010110",
11604 => "101100110011111111111010",
11605 => "101010011110010100001110",
11606 => "101001000110000010101000",
11607 => "101000110011011100000110",
11608 => "101001010001001100101000",
11609 => "101001000110010001001100",
11610 => "101001011000110011011010",
11611 => "101011011010110101001110",
11612 => "101111000011000001010100",
11613 => "110011000101011001101110",
11614 => "110101010100100010000110",
11615 => "110110010001000100000010",
11616 => "110111111001100011001011",
11617 => "111001001010100010011000",
11618 => "111000011000000111000011",
11619 => "110110101100101011100100",
11620 => "110101000001111010101011",
11621 => "110010100100001101110100",
11622 => "110000010010101000101010",
11623 => "101110100101101111001010",
11624 => "101100011010011011011010",
11625 => "101011010100101110110010",
11626 => "101100010010111101100000",
11627 => "101110010111000000110110",
11628 => "110001101011110010001100",
11629 => "110110001101011101000011",
11630 => "111011000111100011000111",
11631 => "111111110010010000010001",
11632 => "000011110111100101101100",
11633 => "000111010000101011001011",
11634 => "001001111010011110111001",
11635 => "001100110011101111000110",
11636 => "010000001011001010011110",
11637 => "010010000000010111000000",
11638 => "010010000010110000001010",
11639 => "010001110110101101001000",
11640 => "010001011111001000000010",
11641 => "010000001101111000110110",
11642 => "001101011111110101010000",
11643 => "001010010100100100011110",
11644 => "001000100000000010111110",
11645 => "000111011000010101100000",
11646 => "000110100100111010011101",
11647 => "000110100011111000011010",
11648 => "000101110000100101100000",
11649 => "000011110000010100111101",
11650 => "000001111011011011100101",
11651 => "000001100001001001110000",
11652 => "000011011100101010101101",
11653 => "000110000000100000010000",
11654 => "000101111010100110000010",
11655 => "000010000110110110000001",
11656 => "111101000110110111011001",
11657 => "111010100111001101111010",
11658 => "111010110001100100101101",
11659 => "111011100110110111100010",
11660 => "111100101100011110101010",
11661 => "111110001111010100111010",
11662 => "111111101111001000110010",
11663 => "111111111000101101010011",
11664 => "111110011100110111001110",
11665 => "111101010100010100010101",
11666 => "111101111111101101010001",
11667 => "000000000100010110001100",
11668 => "000010011111111110100001",
11669 => "000101001101101010111010",
11670 => "000111100011000001100010",
11671 => "000111110100101111100110",
11672 => "000110101000100000000111",
11673 => "000110001110011001101001",
11674 => "000111011110001011001010",
11675 => "001001001011110010011001",
11676 => "001010101000000010101111",
11677 => "001100110010111100010000",
11678 => "001101111001010010001110",
11679 => "001011111011110110010110",
11680 => "001001100001001100011011",
11681 => "000111110101111100111111",
11682 => "000101111110010001111101",
11683 => "000011111001110001011111",
11684 => "000001101011100001001010",
11685 => "111111100001001010101000",
11686 => "111011111000001111111110",
11687 => "110101111010100010010111",
11688 => "101110110100000000100110",
11689 => "100111101001110010100000",
11690 => "100100000001001110110011",
11691 => "100100100101001101100101",
11692 => "100110000101111101101100",
11693 => "101001011101000101011010",
11694 => "101111001000000101010110",
11695 => "110100011100100010011010",
11696 => "111000001001001100000010",
11697 => "111011001010001110110110",
11698 => "111111000111000110101010",
11699 => "000011100010010111000100",
11700 => "001000000101001110011011",
11701 => "001100100100111010111010",
11702 => "001110110001011011000110",
11703 => "001101000010101000011110",
11704 => "000111100111110001110100",
11705 => "000001010100100001000000",
11706 => "111100011101101011000010",
11707 => "111001011100101111000000",
11708 => "111001011100001100111101",
11709 => "111011011001100000101100",
11710 => "111110000100000011111001",
11711 => "000001001000011011001010",
11712 => "000010111010110011010110",
11713 => "000011111010010100001000",
11714 => "000100101100110111110111",
11715 => "000110000010101001011000",
11716 => "001001110110011101101100",
11717 => "001110111101001010110110",
11718 => "010100110000100101011010",
11719 => "011010010110000000011101",
11720 => "011100000011000100111010",
11721 => "011010101001011110001101",
11722 => "011001101010000101101011",
11723 => "011000111111101010110101",
11724 => "011000000111000101000011",
11725 => "010111101001101110100100",
11726 => "010110111101100010101100",
11727 => "010110101111000110000000",
11728 => "010101111110010110010110",
11729 => "001111000111001101010110",
11730 => "000100000111100111110011",
11731 => "111100000111000000101011",
11732 => "110111010101011000111111",
11733 => "110100001001111011011000",
11734 => "110001111101101011101010",
11735 => "110000111001100000010110",
11736 => "110001100101111000011100",
11737 => "110010001111000101011010",
11738 => "110010101100111011111110",
11739 => "110100010010110011101110",
11740 => "110110001110011101111110",
11741 => "110111011010101011011110",
11742 => "110110101000110001000010",
11743 => "110011101011101111111100",
11744 => "101111101000100101001010",
11745 => "101010100110100100000010",
11746 => "100101100110000100111001",
11747 => "100011100010111101010101",
11748 => "100100001011100100001111",
11749 => "100100011000001101100010",
11750 => "100100011111011001100011",
11751 => "100101101111110001100111",
11752 => "101000000000110011100100",
11753 => "101011101101100101111010",
11754 => "101111100001000100100010",
11755 => "110010010010101010011010",
11756 => "110100101101100110110000",
11757 => "110110101010100100100111",
11758 => "110111010010110000010000",
11759 => "110110100001110011000110",
11760 => "110110010000000100000011",
11761 => "110111100000010010101101",
11762 => "111010000010001100000100",
11763 => "111101111110101111010101",
11764 => "000010001011111010001000",
11765 => "000110111000001100000001",
11766 => "001101001101001010101100",
11767 => "010011010001010011111010",
11768 => "010111010111000001101000",
11769 => "011010000110000011101111",
11770 => "011100010011110110100111",
11771 => "011101101110111110011111",
11772 => "011101110101111001000011",
11773 => "011100011111001000010100",
11774 => "011001111010100000111001",
11775 => "010110111011100111100010",
11776 => "010011000110100110011010",
11777 => "001111001110001011101000",
11778 => "001110000111010101011100",
11779 => "001110110111110010100000",
11780 => "001111001000101100111010",
11781 => "001111010101100110010110",
11782 => "010000011011100010000000",
11783 => "010010011101010111011100",
11784 => "010011110111001000000100",
11785 => "010011000101000011001100",
11786 => "010000110100101110100100",
11787 => "001101110010011000000000",
11788 => "001010001101101001110000",
11789 => "000111001011110100101001",
11790 => "000011101101100001010100",
11791 => "111110010001101011110111",
11792 => "110111000011000111010100",
11793 => "101101000001001000010010",
11794 => "100011101101100000111101",
11795 => "100001001000101011110111",
11796 => "100001110101100001011011",
11797 => "100001011001110100000011",
11798 => "100001010011111101110111",
11799 => "100001101101011110101011",
11800 => "100010011101010011011100",
11801 => "100011100101000010011011",
11802 => "100011110100101001010001",
11803 => "100100001000011011110011",
11804 => "100111101101110100100001",
11805 => "101110101111000011010010",
11806 => "110101000110001011110110",
11807 => "111001110011110101100000",
11808 => "111110100010011000001011",
11809 => "000010010011101010001010",
11810 => "000100111100101010010110",
11811 => "000111000010000100100110",
11812 => "001000010100101000011110",
11813 => "001001101111101100100100",
11814 => "001011011101010110001011",
11815 => "001100001011111110100000",
11816 => "001010111000110011100100",
11817 => "000111010110100010110001",
11818 => "000011010010001100010111",
11819 => "000001010111000001100011",
11820 => "000010000010000001010101",
11821 => "000011011010000100011000",
11822 => "000100010100010000111110",
11823 => "000101011011110000100110",
11824 => "000111100111100011100011",
11825 => "001001110100100111110000",
11826 => "001010001001110010111111",
11827 => "001000110101011001001011",
11828 => "001000100001010111010111",
11829 => "001011001111111110010010",
11830 => "001111000001010010100100",
11831 => "010001111001111101010010",
11832 => "010100011110010100011100",
11833 => "010101001011111011000010",
11834 => "010011100100000100110110",
11835 => "010000101110000110100110",
11836 => "001100100011100100011110",
11837 => "001001010111010100011100",
11838 => "000111101001101010100101",
11839 => "000100111110011111001110",
11840 => "000001010101010001111000",
11841 => "111100110000111001001000",
11842 => "110111100010011111100010",
11843 => "110011100100110010111000",
11844 => "110010101001000110100100",
11845 => "110100100011110011010101",
11846 => "110110110011110100111101",
11847 => "111000111001001100101001",
11848 => "111011111100001000101101",
11849 => "111111111111000010010000",
11850 => "000100100000101001010011",
11851 => "000111110000000001011000",
11852 => "001010000010110000101000",
11853 => "001101110001001100110010",
11854 => "010010010100011010111000",
11855 => "010101110000110001100110",
11856 => "010110111000111001000010",
11857 => "010101000011000001100000",
11858 => "010000111101100010011110",
11859 => "001011011010010110101000",
11860 => "000100011010111111110001",
11861 => "111101010011111011100000",
11862 => "111000000111000010111100",
11863 => "110100011010000100010011",
11864 => "110000101000011010111110",
11865 => "101100101111110100001010",
11866 => "101010001000010101001100",
11867 => "101001101011000110010110",
11868 => "101010101001100110011100",
11869 => "101101001101111001010100",
11870 => "110010001011000101000110",
11871 => "111000101001110000100010",
11872 => "111110111000110111010011",
11873 => "000011011001100100011100",
11874 => "000110010001101001111011",
11875 => "000110101101110110011110",
11876 => "000011011101111111100101",
11877 => "111111101000011011001110",
11878 => "111101110101110000101110",
11879 => "111100000111110101010100",
11880 => "111000001000000011100110",
11881 => "110010111111111111111100",
11882 => "101111001101001000010100",
11883 => "101010110111010011100110",
11884 => "100101100110100011110100",
11885 => "100011011000000011111011",
11886 => "100011101100011011010111",
11887 => "100100011011011010111011",
11888 => "100101101000111111101111",
11889 => "100111101010011100011111",
11890 => "101011011110111110100000",
11891 => "110000000011111010011010",
11892 => "110101000010001010110100",
11893 => "111011011000110000001010",
11894 => "000000001111011000101110",
11895 => "000001110000101001011111",
11896 => "000001110010110110010101",
11897 => "000001101101000011100110",
11898 => "000001010111011000000011",
11899 => "111111101100100010101010",
11900 => "111101011101100111011111",
11901 => "111100100111101001110000",
11902 => "111101101010000000010011",
11903 => "000000101011101101000011",
11904 => "000100100110001010011010",
11905 => "001000010011111011010111",
11906 => "001100010011101010000100",
11907 => "010000001001110001111100",
11908 => "010011101010100001001010",
11909 => "010111000010110010111000",
11910 => "011001000011101010010011",
11911 => "011001011100101100011111",
11912 => "011001001111100110011001",
11913 => "011000110001000011100010",
11914 => "011000000011101001001001",
11915 => "010111101010011100101010",
11916 => "010111110101101011011000",
11917 => "010111111100010010001010",
11918 => "011000000010110110101111",
11919 => "011000001100010010101101",
11920 => "010111100110010011111000",
11921 => "010111000011000110110100",
11922 => "010110111011110011100100",
11923 => "010101101010110010100010",
11924 => "010010010010000011110010",
11925 => "001100101110011100111010",
11926 => "000101111101101001110101",
11927 => "111110111110101010000101",
11928 => "110111110100101010000000",
11929 => "110000100011000010000110",
11930 => "101000101011000011101100",
11931 => "100010010001010111111101",
11932 => "100000101111110011000011",
11933 => "100001011111100001110001",
11934 => "100001010100110110100100",
11935 => "100001101010010000011111",
11936 => "100010011010010100000111",
11937 => "100010110000100001100111",
11938 => "100011011110000111011110",
11939 => "100100010011011010101111",
11940 => "100100101010101011100000",
11941 => "100101000010100101011011",
11942 => "100111001001010110000100",
11943 => "101011000011101110001010",
11944 => "101110000000111111101110",
11945 => "101111011111000100100100",
11946 => "110000110001010010000010",
11947 => "110001111011011011111110",
11948 => "110010011110111111110000",
11949 => "110001110110010010101110",
11950 => "110010000101011011001110",
11951 => "110101100101000010010000",
11952 => "111001111001100100010100",
11953 => "111100011001100110110011",
11954 => "111101001011101001100001",
11955 => "111101011001101110110010",
11956 => "111111000001101011011011",
11957 => "000010000100111010110110",
11958 => "000100110010011000011100",
11959 => "000111010000100111001011",
11960 => "001010100010000001001001",
11961 => "001110000100110011110000",
11962 => "010001010010111010100000",
11963 => "010100100110110000011110",
11964 => "010110110100000000010100",
11965 => "010110011000010111001010",
11966 => "010100111111011001101010",
11967 => "010100111111011111011000",
11968 => "010110011010100110001110",
11969 => "010111111100011001100010",
11970 => "011000111110111100110010",
11971 => "011010011111111010010011",
11972 => "011100010100001101101111",
11973 => "011100110010001000001110",
11974 => "011100011111101110100111",
11975 => "011100100101011101010010",
11976 => "011100001010011010011000",
11977 => "011011010011001001001111",
11978 => "011010100101001011010101",
11979 => "011001100010001101010001",
11980 => "011000100001011001100000",
11981 => "010111110111111100110010",
11982 => "010111001011000101100010",
11983 => "010110001000001001110010",
11984 => "010100010001010011101000",
11985 => "010001110010000010110000",
11986 => "001111101010101010111010",
11987 => "001101111000010000111100",
11988 => "001010101000110111011000",
11989 => "000101100101001011110010",
11990 => "000000100000101100110011",
11991 => "111010111110011111011110",
11992 => "110011010100001001110110",
11993 => "101010011101010100111000",
11994 => "100011110000110000101001",
11995 => "100001101111011010011111",
11996 => "100001110101011100111110",
11997 => "100001100010110100000011",
11998 => "100001101100001111100010",
11999 => "100001000110111100111101",
12000 => "100001011110000000010011",
12001 => "100110111101010111100000",
12002 => "101110111100000110010000",
12003 => "110101111111100100011000",
12004 => "111100100011111101000001",
12005 => "000010010100110101110100",
12006 => "000111010000111000101000",
12007 => "001010011100101100111111",
12008 => "001010011110000110001001",
12009 => "001001100011010111100100",
12010 => "001000011010010101110101",
12011 => "000100111001100010001001",
12012 => "111111110011010011011101",
12013 => "111010000110100001010011",
12014 => "110011011111101000111100",
12015 => "101101111101001100001100",
12016 => "101010011001101101010110",
12017 => "100110110011110100111001",
12018 => "100011101110010010010100",
12019 => "100011110111010111100110",
12020 => "100101111011110100000011",
12021 => "100111000101101011010011",
12022 => "101000001100101001111110",
12023 => "101010111011110010101000",
12024 => "101111101000101001000100",
12025 => "110101101000100110010100",
12026 => "111011011011001010110111",
12027 => "000000111101111111100100",
12028 => "000110010110100100010100",
12029 => "001001111000101010001100",
12030 => "001010110011011001101001",
12031 => "001010011110010000101110",
12032 => "001001110101100111100000",
12033 => "000111101110111010001111",
12034 => "000100010111011111000100",
12035 => "000001101010011111100011",
12036 => "111111010010100100000100",
12037 => "111100111101010101011000",
12038 => "111011011110001010001010",
12039 => "111011001011001001010011",
12040 => "111101001011101111110011",
12041 => "000001010010111100001000",
12042 => "000110100001011000111000",
12043 => "001100111001001010001100",
12044 => "010010111101011001010110",
12045 => "010111110111010001100010",
12046 => "011011101000100110110011",
12047 => "011100101111011100110111",
12048 => "011011101111100111001001",
12049 => "011010001011100101100011",
12050 => "010111001110011011011000",
12051 => "010010111011001110010000",
12052 => "001110010011001110100100",
12053 => "001010001010000001100001",
12054 => "000111110101111111010010",
12055 => "000110111011101011101000",
12056 => "000110000000110001100111",
12057 => "000101111010111101001111",
12058 => "000111100011010010110000",
12059 => "001001011101011001110011",
12060 => "001010100010001000001000",
12061 => "001011000011100100011110",
12062 => "001010000100000000011001",
12063 => "000110100001101111111111",
12064 => "000000111000111100010000",
12065 => "111010010101111010111000",
12066 => "110101101011101011110010",
12067 => "110001111100010111000000",
12068 => "101010100010111001010010",
12069 => "100011010000010111110011",
12070 => "100001101100110000010001",
12071 => "100010001100101101000111",
12072 => "100010010101011111110001",
12073 => "100011110000110101001111",
12074 => "100100111100001111011100",
12075 => "100101001011101011000111",
12076 => "100110000010011101000001",
12077 => "100111011010001101100101",
12078 => "101000101111011010110000",
12079 => "101010001101010101110000",
12080 => "101100000110001101000100",
12081 => "101110001111101100010010",
12082 => "101111101011011101001010",
12083 => "110000000010111001011110",
12084 => "110000011110000101111110",
12085 => "110001001011111011001000",
12086 => "110001100111011010010110",
12087 => "110011011101100101111100",
12088 => "110111101011111111000011",
12089 => "111100001000101110000011",
12090 => "000000001101000101111101",
12091 => "000100010100011101001001",
12092 => "000111010010110101001110",
12093 => "001000100000000101101111",
12094 => "001000011100101010100100",
12095 => "001000100011110101111001",
12096 => "001001010110111010101110",
12097 => "001001000011101011001011",
12098 => "000111011011101101010011",
12099 => "000110000100101010000001",
12100 => "000101011111010101001011",
12101 => "000100111111101101101010",
12102 => "000011110110010010001010",
12103 => "000011101011001110010000",
12104 => "000101111100110000000010",
12105 => "001001011101110011101000",
12106 => "001110010100111101010100",
12107 => "010100010101111010010010",
12108 => "011000111010011010011101",
12109 => "011011001001011101001101",
12110 => "011100000101000100011101",
12111 => "011100111110001100101101",
12112 => "011101101010101011111001",
12113 => "011100111000001110100011",
12114 => "011011110001011011111011",
12115 => "011011000110001000110001",
12116 => "011001110111111001001001",
12117 => "011001001110111101001101",
12118 => "011000110111111101000101",
12119 => "010110011011100110111100",
12120 => "010010001010000010011000",
12121 => "001100110010111100101010",
12122 => "000110000000010000000001",
12123 => "111101111101111101101001",
12124 => "110101011011111101100010",
12125 => "101110001111101101100000",
12126 => "101001110110000111011110",
12127 => "100111001001011110011001",
12128 => "100101010111101010001101",
12129 => "100110011011000111010110",
12130 => "101010111010100100110100",
12131 => "110000100101100101110100",
12132 => "110110110011110010101111",
12133 => "111101111001010111110110",
12134 => "000100010011000101011000",
12135 => "001000111011110011011011",
12136 => "001100000100010111000000",
12137 => "001110010011011001011000",
12138 => "001111001010110100100110",
12139 => "001101100101101010100010",
12140 => "001011100111110000001100",
12141 => "001010100011000101011011",
12142 => "000111100010101110011110",
12143 => "000010101110100100011010",
12144 => "111110011111101000110110",
12145 => "111001101111110110100110",
12146 => "110010101011110101100110",
12147 => "101010001001111110100000",
12148 => "100011101011001001100001",
12149 => "100001101111110101101101",
12150 => "100010100100100111000001",
12151 => "100011110100010010010111",
12152 => "100101010100000101110101",
12153 => "100111000010001101000010",
12154 => "101000001011110101000010",
12155 => "101001000111010100101000",
12156 => "101100001110100111000100",
12157 => "110001110010000001001110",
12158 => "111000000001111010011110",
12159 => "111111010000100000101001",
12160 => "000110000100100001001110",
12161 => "001001100010100111111011",
12162 => "001010011110110011000111",
12163 => "001001111110010101100101",
12164 => "000111000011001000110011",
12165 => "000010100001001100000010",
12166 => "111110110010001000101011",
12167 => "111100100101001011011101",
12168 => "111010110010101000111000",
12169 => "111001000100001110110110",
12170 => "110111110011010101110001",
12171 => "110111000011001101010111",
12172 => "110111100110011011100101",
12173 => "111001111010101001000101",
12174 => "111101011010110101110101",
12175 => "000001110001100101001110",
12176 => "000111000010100101100000",
12177 => "001101011111000111111110",
12178 => "010011110100101100111010",
12179 => "011000011010010011010000",
12180 => "011100001101000000011101",
12181 => "011110110101111111101101",
12182 => "011110100100100001111111",
12183 => "011101000000100011000110",
12184 => "011100000010010011101100",
12185 => "011011000100111010100101",
12186 => "011001110001110101000001",
12187 => "011000101100000010101111",
12188 => "010111011110010011001010",
12189 => "010100010101111010001100",
12190 => "001111010110110111100100",
12191 => "001010110111011011011110",
12192 => "000111100101011111010100",
12193 => "000101100010001010110100",
12194 => "000101000101111101010101",
12195 => "000101000101111111111011",
12196 => "000100010011010110011100",
12197 => "000011011010111011110111",
12198 => "000011111100010010100010",
12199 => "000101011010011110100000",
12200 => "000101010011100001110010",
12201 => "000001110100010001000011",
12202 => "111011100000100010010000",
12203 => "110101010001011100000110",
12204 => "101111110100000001001010",
12205 => "101000101000010101000000",
12206 => "100010010011100110000110",
12207 => "100001001010100000010101",
12208 => "100010010111110110101001",
12209 => "100010111110100001111000",
12210 => "100011101111101110011110",
12211 => "100100011000101001001111",
12212 => "100100111100001011010000",
12213 => "100101110101001110101001",
12214 => "100110010001110111110110",
12215 => "100110100011010110110000",
12216 => "101000000100100100011000",
12217 => "101011100000000000100000",
12218 => "101111111011100011111010",
12219 => "110011110101001011000110",
12220 => "110110100011011110011111",
12221 => "111000101001100100011001",
12222 => "111011011100110001000010",
12223 => "111111010011010001001111",
12224 => "000011010001111010001110",
12225 => "000110110011011101111110",
12226 => "001001110101100010100101",
12227 => "001101011011010000001000",
12228 => "010010010001001010110010",
12229 => "010110100100101110111000",
12230 => "011000100011011101000101",
12231 => "011000011110000000001010",
12232 => "011000000110110100001011",
12233 => "011000011011100110100110",
12234 => "010111101111000000000110",
12235 => "010101110100111011111110",
12236 => "010100110111100101101100",
12237 => "010100011101110100011000",
12238 => "010011011100000011000110",
12239 => "010010111010100101111110",
12240 => "010011110100110111010100",
12241 => "010101000000010011110100",
12242 => "010101001110110001010100",
12243 => "010101100111000101100000",
12244 => "010111000101000001111010",
12245 => "011000001000111011001111",
12246 => "010111101111011001110110",
12247 => "010110111011101001011110",
12248 => "010110110110111011000010",
12249 => "010101100110011011100010",
12250 => "010000010100000010101010",
12251 => "001000101011000110010110",
12252 => "000001001001000011110101",
12253 => "111000111000010000010101",
12254 => "101111100111100001111000",
12255 => "100111000111011001001100",
12256 => "100010010010110100000101",
12257 => "100001111000010010110001",
12258 => "100010001010001011001011",
12259 => "100001100000110000111001",
12260 => "100001100100010111111111",
12261 => "100001111000011011001010",
12262 => "100001100101000111110111",
12263 => "100001010100010101000101",
12264 => "100010100101101000100011",
12265 => "100110100011110000110001",
12266 => "101011111110100010010100",
12267 => "110001010010011011001100",
12268 => "110110000110101001000111",
12269 => "111001110100100010001101",
12270 => "111101000011100111010001",
12271 => "000001001010100011111100",
12272 => "000101011011010000110001",
12273 => "000111101111000101111111",
12274 => "000111100011111010111010",
12275 => "000110100100110001110111",
12276 => "000101011111101011100101",
12277 => "000011000101111111110101",
12278 => "111111010100011111101101",
12279 => "111100000100110111010000",
12280 => "111010011100101100100100",
12281 => "111001101101010100000011",
12282 => "111001111100000100000111",
12283 => "111011100011000000011100",
12284 => "111101010000111110101110",
12285 => "111111111100110110101010",
12286 => "000101101010011111110100",
12287 => "001100000100010000001110",
12288 => "010000001010001010011010",
12289 => "010010100111110011111110",
12290 => "010100111110011100001000",
12291 => "010110100111001000011000",
12292 => "010101010011111011110110",
12293 => "010001011010010111101110",
12294 => "001101100100111000110000",
12295 => "001010011000000100110100",
12296 => "000111001100100100001010",
12297 => "000011010100101001101101",
12298 => "111101101000011111011100",
12299 => "110110000000100000010011",
12300 => "101101001111010010111100",
12301 => "100101111101110011000011",
12302 => "100011000101101101101001",
12303 => "100011001011011101011100",
12304 => "100100000010110111110000",
12305 => "100111001000110000011111",
12306 => "101101000010111000110010",
12307 => "110011010001010000011010",
12308 => "111000101110011000110010",
12309 => "111110001110111101100101",
12310 => "000010111101011011000000",
12311 => "000110101110010001110000",
12312 => "001011100010011010011101",
12313 => "010000111100111011000100",
12314 => "010100101011111000101000",
12315 => "010101101001011111011010",
12316 => "010011100111011110111100",
12317 => "010000001000011000011010",
12318 => "001100100101101010110110",
12319 => "001001000111011010101010",
12320 => "000110110000011101100100",
12321 => "000101011101100110010110",
12322 => "000100010001001111000010",
12323 => "000011001000010001000111",
12324 => "000001000111111011101000",
12325 => "111110101000100010001000",
12326 => "111101100111001011100000",
12327 => "111101101010101111110000",
12328 => "111110001100011011000011",
12329 => "000000001001001110001000",
12330 => "000011010011110110111001",
12331 => "000110001010000011101100",
12332 => "000111111011101100101010",
12333 => "001001001010000001000000",
12334 => "001001110100100100011100",
12335 => "001001011010111111010000",
12336 => "001000100001110111011010",
12337 => "000111111001001001001011",
12338 => "000111100001101010101000",
12339 => "000101111010001000110101",
12340 => "000000011101000101110000",
12341 => "110111111111010110110101",
12342 => "110000101010100110101010",
12343 => "101011100001100111100010",
12344 => "100110100111001100001101",
12345 => "100011001001101010111101",
12346 => "100011010010110110000101",
12347 => "100100011101110000101011",
12348 => "100100101111000001110110",
12349 => "100101101101011001010001",
12350 => "100110100100010011000011",
12351 => "100111000011000100011011",
12352 => "101010001011000011001100",
12353 => "101111010111001011110000",
12354 => "110011010111010010001000",
12355 => "110101110001111011000111",
12356 => "111000000100110101110110",
12357 => "111010111001000001000101",
12358 => "111100101000110000001101",
12359 => "111100001001000100011101",
12360 => "111011010011111011110100",
12361 => "111100001010011111011111",
12362 => "111111001000000001000110",
12363 => "000011101110110110110100",
12364 => "001001000000101110111100",
12365 => "001111010100100110110100",
12366 => "010111000100010010001000",
12367 => "011100111010001111010101",
12368 => "011101100111101011011101",
12369 => "011100001001111110111111",
12370 => "011011111111111011010101",
12371 => "011011100100011001011101",
12372 => "011010011101111101010001",
12373 => "011010000111111111111110",
12374 => "011001100011101000101001",
12375 => "011000111101011100111011",
12376 => "011001000001010101011101",
12377 => "011000101000100111011011",
12378 => "011000011101101000011001",
12379 => "011000100001100101111011",
12380 => "010110101110110100101100",
12381 => "010010111110110011001110",
12382 => "001110001100100000100000",
12383 => "001001001011001010110110",
12384 => "000100100001000011111010",
12385 => "111111010000111011001001",
12386 => "111000111011010000101001",
12387 => "110001110101110000010110",
12388 => "101010001110111100001100",
12389 => "100100001000100000110101",
12390 => "100001101101010001101011",
12391 => "100001110001000100010111",
12392 => "100010000011110000010001",
12393 => "100011001011010100110001",
12394 => "100110010001110000100000",
12395 => "101001110001100110010010",
12396 => "101100001001111101011100",
12397 => "101101101000000011111000",
12398 => "101110011100011011111110",
12399 => "101110111011111111110110",
12400 => "101110100011010011100110",
12401 => "101100100100110000100000",
12402 => "101010001101011000110010",
12403 => "101000000001101111010100",
12404 => "100101101111010100010101",
12405 => "100100101001111101111001",
12406 => "100101001101011111110101",
12407 => "100101111011011010101001",
12408 => "100110011001101001001001",
12409 => "100111000001101101000101",
12410 => "100111100010110111110011",
12411 => "101000101100100110001010",
12412 => "101011110111111000101100",
12413 => "110000010111100010101100",
12414 => "110101010010011011110010",
12415 => "111011010110111101111110",
12416 => "000010001011110111001011",
12417 => "001000010101011111111001",
12418 => "001101010001101110000010",
12419 => "010001100111101011001010",
12420 => "010110011111001001000010",
12421 => "011011000111001111101100",
12422 => "011101100010110100000100",
12423 => "011101110110011001001111",
12424 => "011101101010011101000011",
12425 => "011110000101110111010101",
12426 => "011101110001000111100111",
12427 => "011010011111010111000011",
12428 => "010101001111011011110110",
12429 => "001111101101101001011010",
12430 => "001010010010111010111101",
12431 => "000110100001011001001000",
12432 => "000101000011101010000100",
12433 => "000100100010000100101011",
12434 => "000100101011111001110000",
12435 => "000110011001100000011111",
12436 => "001001010011110101011110",
12437 => "001011101101111111000000",
12438 => "001101001011001111111000",
12439 => "001110110001101100110100",
12440 => "010000110111010101111110",
12441 => "010011011010011000111110",
12442 => "010101111010011001011010",
12443 => "010111000001101110100110",
12444 => "010110100010101100001110",
12445 => "010100100010110110101010",
12446 => "010000111001100010000010",
12447 => "001100110101011110001110",
12448 => "001001010110010111001100",
12449 => "000110000110000001111111",
12450 => "000010011011001111110100",
12451 => "111101110011110110001110",
12452 => "111000100111101010111011",
12453 => "110011100111000101110110",
12454 => "101110011100001111011100",
12455 => "101000110000100010111000",
12456 => "100100011000100100110101",
12457 => "100011110111001000000111",
12458 => "100110100111101101101101",
12459 => "101010011000111101000100",
12460 => "101110111011011011100100",
12461 => "110100011011001111010000",
12462 => "111001111111111111110100",
12463 => "111111001111010111001111",
12464 => "000100011011100000101011",
12465 => "001001110101101001011001",
12466 => "001111000100101110100100",
12467 => "010011000111111110100100",
12468 => "010101010011001011001000",
12469 => "010101010001000100001100",
12470 => "010010100111100111011100",
12471 => "001101100010011111010000",
12472 => "000111110110101010110100",
12473 => "000011010000000100011111",
12474 => "111111010001010100101100",
12475 => "111011111011011110011000",
12476 => "111010000000000110100001",
12477 => "111000000101100010000110",
12478 => "110101010011011011010100",
12479 => "110011010001110111001100",
12480 => "110010101000011100000000",
12481 => "110010110101111001000110",
12482 => "110011111100110101101000",
12483 => "110100111001010001000001",
12484 => "110100010101100010010110",
12485 => "110011111000111111100100",
12486 => "110101010010111010100100",
12487 => "110111000000101010011110",
12488 => "111000011110010000001000",
12489 => "111011011011011110010011",
12490 => "111111010100100010001111",
12491 => "000001110011101110101110",
12492 => "000001111000101111110011",
12493 => "000000101100010010010110",
12494 => "000000111110011010011111",
12495 => "000011101101010010111101",
12496 => "000110101000001101100111",
12497 => "000111111100000110110110",
12498 => "001001000110010111010001",
12499 => "001100010000011010000100",
12500 => "010000100011010001010100",
12501 => "010100100110110110111100",
12502 => "011000001011100110110001",
12503 => "011001100001100110001010",
12504 => "011000110001011101101101",
12505 => "011000011010110000101111",
12506 => "010111111100000110001000",
12507 => "010111000011010010010010",
12508 => "010110101100011001000010",
12509 => "010101111110001110110000",
12510 => "010110000000000000101010",
12511 => "010101010010000101001000",
12512 => "001100111100011111111000",
12513 => "111110111010001111101100",
12514 => "110011110011010110111100",
12515 => "101011110010100001001000",
12516 => "100100111101101101111011",
12517 => "100001110011001110010011",
12518 => "100001010101001010111011",
12519 => "100010000101001001111100",
12520 => "100110111000010110110101",
12521 => "101111100110010101000010",
12522 => "111000100011000010001101",
12523 => "000000000011100100000100",
12524 => "000101001111111111000010",
12525 => "000111010111101110001011",
12526 => "000110110111000110010000",
12527 => "000100010010111100010011",
12528 => "000001000010101001110001",
12529 => "111110100101101001101101",
12530 => "111100011110101101111100",
12531 => "111001111111000100010101",
12532 => "110111100001000101010110",
12533 => "110101100011000110011100",
12534 => "110011110111011011100100",
12535 => "110001110001001000111010",
12536 => "101111011101001111000010",
12537 => "101101110111101010000110",
12538 => "101100000011000010011100",
12539 => "101000010110100111011110",
12540 => "100100111010110000100111",
12541 => "100100110010000101111000",
12542 => "100110000011110110000111",
12543 => "100110100011111000000001",
12544 => "100111011001100101110011",
12545 => "100111111010011010001001",
12546 => "101000101011101100000100",
12547 => "101110001011100111101010",
12548 => "110111101000111000100001",
12549 => "000000010000000110000000",
12550 => "000111011011011111100000",
12551 => "001101010000101110100000",
12552 => "010000100110010100101010",
12553 => "010010001110100101100100",
12554 => "010010110101111001110000",
12555 => "010010000000110111000100",
12556 => "001111011110011001101100",
12557 => "001011001001110100011101",
12558 => "000110000101011100100010",
12559 => "000001100001010110001101",
12560 => "111101001101111010001011",
12561 => "111001011101000000001001",
12562 => "110111111100001111101000",
12563 => "111000111101110111010010",
12564 => "111010110010100111110000",
12565 => "111100000011101010001001",
12566 => "111100101011101010111010",
12567 => "111101011100100010100010",
12568 => "111111001100100001110010",
12569 => "000001110100101000111101",
12570 => "000100111000011000001101",
12571 => "001000010101011001001111",
12572 => "001011111111010011010101",
12573 => "001111010010110100001010",
12574 => "010001000000110110000100",
12575 => "001111111101000101001000",
12576 => "001101010011100011000000",
12577 => "001011101010110001001000",
12578 => "001011011100101111010100",
12579 => "001010111100001011011101",
12580 => "001001011011001001011101",
12581 => "000111100001001101100011",
12582 => "000101000011101110000001",
12583 => "000001011111111111011000",
12584 => "111101100101011101101100",
12585 => "111010011101000111001011",
12586 => "111000011101010011011100",
12587 => "110111100111111010001000",
12588 => "111000010011110000110000",
12589 => "111010101111100111010000",
12590 => "111110001001101010101101",
12591 => "000001100111101110110000",
12592 => "000101001110000001011110",
12593 => "001000111010101111000000",
12594 => "001100001000100000101010",
12595 => "001110110001100000101000",
12596 => "010001010011000001010110",
12597 => "010011100111101010011010",
12598 => "010100100000101010111010",
12599 => "010011000100010011001100",
12600 => "010000010111000011010000",
12601 => "001101111110111100000000",
12602 => "001100010110000001101100",
12603 => "001011000000010111001011",
12604 => "001000111011001011010101",
12605 => "000101011100010010010011",
12606 => "000001010101001111010100",
12607 => "111100111011101111100011",
12608 => "110111110001101001011111",
12609 => "110011000110001010111110",
12610 => "110000100000111000010110",
12611 => "101111101101110111111010",
12612 => "110000011100111101011100",
12613 => "110011010001100110101110",
12614 => "110111101100010000001010",
12615 => "111100001000111011010000",
12616 => "111111010010101010101110",
12617 => "000000111001001000110111",
12618 => "000001100100000001000010",
12619 => "000010011101000101010000",
12620 => "000100000011010000110111",
12621 => "000100000001011001010111",
12622 => "000000001111010011001010",
12623 => "111010110000101110101111",
12624 => "110110001100101011001110",
12625 => "110011101101110111010100",
12626 => "110100011101011011011011",
12627 => "110111000110100010000000",
12628 => "111001011110000111101000",
12629 => "111011111010001110010100",
12630 => "111110010011001101001010",
12631 => "000000010011100011101001",
12632 => "000011011110111110001001",
12633 => "001000010001010111110110",
12634 => "001101001011010000001000",
12635 => "010000101111001000101010",
12636 => "010011001001101001011100",
12637 => "010110010101100001000110",
12638 => "011001101010000100011101",
12639 => "011010011010011100101101",
12640 => "011001011001000001000011",
12641 => "011000100001001010101000",
12642 => "010111101100000110101000",
12643 => "010110101000001011010010",
12644 => "010011110000100000101010",
12645 => "001101011001100011000110",
12646 => "000101010001101010110110",
12647 => "111101100011110100100101",
12648 => "110111000011101101000010",
12649 => "110010111001011100001110",
12650 => "110000111100001000000110",
12651 => "101111110011011010011100",
12652 => "101111100010110101001010",
12653 => "110001011110000101111110",
12654 => "110101110011100110100010",
12655 => "111010010100000001001000",
12656 => "111101000110000111010011",
12657 => "111111011101101101111000",
12658 => "000010110011110101110100",
12659 => "000110010000111011001001",
12660 => "001000100001100000010011",
12661 => "001000101101000110001010",
12662 => "000110011101010100011100",
12663 => "000010000000111011100110",
12664 => "111011101010111010001011",
12665 => "110011011110110001000110",
12666 => "101010010110110101101010",
12667 => "100011110010101100000101",
12668 => "100010000001011111100011",
12669 => "100010001110100101011011",
12670 => "100010011010011000011111",
12671 => "100011011101011010000111",
12672 => "100100010101110010111000",
12673 => "100101011000001111101011",
12674 => "101001011111001101100000",
12675 => "101111111010110010100100",
12676 => "110101111110111111100001",
12677 => "111010100000001111111011",
12678 => "111100011100001001000100",
12679 => "111100110110111010110000",
12680 => "111101101110110101100110",
12681 => "111110011010010000001110",
12682 => "111110101001110111100000",
12683 => "111111010111010101011010",
12684 => "000000101000101100101000",
12685 => "000011001001011111100100",
12686 => "000110111010011000011010",
12687 => "001010010001100100110001",
12688 => "001100010101000101011010",
12689 => "001101000010011110000110",
12690 => "001100111010101101011010",
12691 => "001100111101011010101100",
12692 => "001101001011010000000110",
12693 => "001100101110101110011000",
12694 => "001011001001101101101000",
12695 => "001001000101100000000011",
12696 => "000111111100100010111111",
12697 => "001000001110000010110100",
12698 => "001001001000011101111010",
12699 => "001001111101111110000000",
12700 => "001011000110011001011110",
12701 => "001101010000110011001000",
12702 => "001111011011011110010010",
12703 => "001111101011110010100100",
12704 => "001101111000001100110000",
12705 => "001010101010101001010001",
12706 => "000110100010010100100001",
12707 => "000010101001001001000011",
12708 => "111111000110001111101101",
12709 => "111010110101001001100011",
12710 => "110110001110111011111101",
12711 => "110010000111001101101000",
12712 => "101110011101100001001000",
12713 => "101011001100011010111010",
12714 => "100111100111110110111101",
12715 => "100100001010100011000101",
12716 => "100010101111100011000011",
12717 => "100011010101010111000100",
12718 => "100100011111011001100001",
12719 => "100101011101000111001110",
12720 => "100110010111100101100001",
12721 => "101000010010100110101000",
12722 => "101011010110000001011100",
12723 => "101110101111101110110000",
12724 => "110010010001001101010110",
12725 => "110101001011100000011110",
12726 => "110111000010101111100011",
12727 => "111000100101100110011001",
12728 => "111010011000100011100100",
12729 => "111101000000111000100010",
12730 => "000000000101100101001010",
12731 => "000001101000111101000110",
12732 => "000001100001110000011000",
12733 => "000001110100110010010101",
12734 => "000011100000101010100000",
12735 => "000101111111010110011011",
12736 => "001000000000011110100011",
12737 => "001001000101010010110010",
12738 => "001010110110001110011111",
12739 => "001101110100100010110100",
12740 => "010000001011101011100010",
12741 => "010001111000101100110010",
12742 => "010100001100111100001000",
12743 => "010111011111111010000100",
12744 => "011011100101001010010100",
12745 => "011110100010010001011011",
12746 => "011110111101001110110111",
12747 => "011110010110000101100011",
12748 => "011101110100001111101101",
12749 => "011101010010010100100010",
12750 => "011100100001000001110111",
12751 => "011010110110111000000011",
12752 => "011000111110111110100011",
12753 => "011000010001001100011110",
12754 => "011000000010000010111101",
12755 => "010110101101011111101110",
12756 => "010100011001011110111100",
12757 => "010001111110000001011010",
12758 => "001110100100100011111100",
12759 => "001000000111111001001101",
12760 => "111110000000000011001001",
12761 => "110010011101110001101010",
12762 => "101001110000111100011000",
12763 => "100110101001110100110101",
12764 => "100111111110011000100101",
12765 => "101010110010110000101000",
12766 => "101101101111111000010000",
12767 => "110001100111101011011110",
12768 => "110111010100101111111000",
12769 => "111101101101101010000011",
12770 => "000010000101000011100100",
12771 => "000011110011010010010100",
12772 => "000100100000110110111101",
12773 => "000011101110100011010100",
12774 => "000000001100110010010010",
12775 => "111011010100000111001110",
12776 => "110110001111100000101110",
12777 => "110001000010101111111110",
12778 => "101100100011011110000000",
12779 => "101010000111101011010000",
12780 => "101011010010100001011110",
12781 => "110000000000111110111010",
12782 => "110101110001000001011000",
12783 => "111010001001001101101000",
12784 => "111100100000110111011001",
12785 => "111110001100011101110000",
12786 => "000000110111010110110100",
12787 => "000100001000000111011000",
12788 => "000110000010101110111101",
12789 => "000101011101011010010000",
12790 => "000100000011111110111001",
12791 => "000100001011110000001111",
12792 => "000100011010101110001000",
12793 => "000010101000101100100001",
12794 => "111111110110101001010010",
12795 => "111100110110010101000111",
12796 => "111001101011011100001101",
12797 => "111000000110111111001101",
12798 => "111000010100001101110100",
12799 => "110111101010011100110101",
12800 => "110101001011011100100111",
12801 => "110010001011111010011110",
12802 => "110000000011011100110110",
12803 => "101110111111011111101100",
12804 => "101110001010000110101110",
12805 => "101111001000100100110000",
12806 => "110100010000001100111110",
12807 => "111010101111011001100000",
12808 => "111111010000110000010101",
12809 => "000010110110100000100010",
12810 => "000110101110001001111111",
12811 => "001010011001101110010100",
12812 => "001100100101110001110110",
12813 => "001100010010001010101010",
12814 => "001010011000001011100010",
12815 => "000111010001010110100001",
12816 => "000001111000010101000101",
12817 => "111010010101101111001101",
12818 => "110010010000100111011000",
12819 => "101011100100001100110000",
12820 => "100111110000010001111011",
12821 => "100111000101110111110111",
12822 => "101000110011100001101010",
12823 => "101100111000000101110110",
12824 => "110100011101100010011110",
12825 => "111110110010111100100111",
12826 => "001001001000110111101001",
12827 => "010010010101100001111010",
12828 => "011001111011100110111001",
12829 => "011110001011110101011011",
12830 => "011110100110101100011000",
12831 => "011101011110110000111111",
12832 => "011100110000001110010111",
12833 => "011011110000011011100000",
12834 => "011001010110100111101101",
12835 => "010101111110100110101010",
12836 => "010010111110101010111010",
12837 => "010000110000100111101000",
12838 => "001110011010010001000110",
12839 => "001011110011011100010100",
12840 => "001001010100000110001111",
12841 => "000110100001000000011101",
12842 => "000011010100011110111000",
12843 => "111111010111101101101101",
12844 => "111010001011100001110000",
12845 => "110100111110001101100100",
12846 => "110000101001101000100110",
12847 => "101100001011111000000000",
12848 => "100111011011110001100101",
12849 => "100100101000100101110001",
12850 => "100100110000000011000010",
12851 => "100101101100001011010000",
12852 => "100110010001111001100101",
12853 => "100110110100100011001000",
12854 => "100111011110111000011011",
12855 => "101001010010111011110000",
12856 => "101100001010110100111010",
12857 => "101110100101011010011000",
12858 => "110000000110111101000110",
12859 => "110000011101111100101100",
12860 => "101111011111111001011010",
12861 => "101101010111011111101100",
12862 => "101010011011011100000100",
12863 => "101000011111011101010110",
12864 => "101000011010011110101000",
12865 => "101000111011100000111100",
12866 => "101001011101001011010100",
12867 => "101001111001010000100000",
12868 => "101010011110011100010100",
12869 => "101100100111010000000000",
12870 => "110000101100011010001110",
12871 => "110101110001101101100000",
12872 => "111100000011010100101101",
12873 => "000011011111101001101101",
12874 => "001010101000100100101011",
12875 => "010001001001010111111110",
12876 => "010111000101110011011100",
12877 => "011011011101100000010011",
12878 => "011101111100101001100111",
12879 => "011110101001100101010001",
12880 => "011110010111111101011101",
12881 => "011110011011100001010101",
12882 => "011110011101110111000011",
12883 => "011110010010100010001101",
12884 => "011110010001000111011110",
12885 => "011110001100001011010111",
12886 => "011110010101100100000101",
12887 => "011110001101011000001011",
12888 => "011101011110101110001101",
12889 => "011101000101100100001101",
12890 => "011100110011101011011100",
12891 => "011100100010011001010011",
12892 => "011100011110111100111010",
12893 => "011100000011100101110101",
12894 => "011011100110100000010100",
12895 => "011011000000001100100101",
12896 => "011001111101001011110111",
12897 => "011001011011011100011111",
12898 => "010111110010000000001110",
12899 => "010001111000001010101010",
12900 => "001001000010000100111011",
12901 => "000001000001001000100100",
12902 => "111010101110010000001111",
12903 => "110100111011111101111011",
12904 => "101111010111010011010100",
12905 => "101010111111011101100000",
12906 => "101000000110111010000100",
12907 => "100100111111100010100011",
12908 => "100001110011101011011001",
12909 => "100001010100011000000011",
12910 => "100010101001011011111010",
12911 => "100011010001100001011000",
12912 => "100011111111101110110111",
12913 => "100101101010101011000011",
12914 => "101000000100001110000100",
12915 => "101011000000100110011010",
12916 => "101110001101100111101110",
12917 => "110001111110001110101010",
12918 => "110110001011111110110011",
12919 => "111010110000111010100010",
12920 => "111111100111001110111110",
12921 => "000011011010101101101011",
12922 => "000101110101011111000101",
12923 => "000110111001110101101101",
12924 => "000101111101100011100101",
12925 => "000100010101001010100010",
12926 => "000011010000000011010111",
12927 => "000000101110101011101101",
12928 => "111011010000111011000010",
12929 => "110101101100111010111000",
12930 => "110011010000011000000000",
12931 => "110010101011101011100110",
12932 => "110001101011111011101010",
12933 => "110000110111001010000100",
12934 => "110010100110100100110100",
12935 => "111000000111011111100000",
12936 => "111111000001101000011100",
12937 => "000100110111000110101000",
12938 => "001010010001100001001100",
12939 => "001111011010000110101010",
12940 => "010010111001100011000010",
12941 => "010100010001010100001000",
12942 => "010100000000001111010000",
12943 => "010011011000110011111100",
12944 => "010100000001000100000110",
12945 => "010100111111101001101000",
12946 => "010011010000011111011110",
12947 => "001111010011110110100100",
12948 => "001011111000101010010000",
12949 => "000111111100001000110110",
12950 => "000010111001100010110011",
12951 => "111111000111110010010001",
12952 => "111100011111101001000011",
12953 => "111001011011110110100010",
12954 => "110110010110001000110010",
12955 => "110100011100000001111100",
12956 => "110011101000001001110110",
12957 => "110011010011001100110010",
12958 => "110100111101101110001000",
12959 => "111010000000101101011100",
12960 => "000001000001101001111101",
12961 => "001000010101110100101000",
12962 => "001111011001101100011110",
12963 => "010101101100110111100000",
12964 => "011001110110100111100010",
12965 => "011010101100100101000001",
12966 => "011000111110110111110001",
12967 => "010101101000110011010110",
12968 => "010000110000100100100100",
12969 => "001010010101110110110001",
12970 => "000010101010101010100011",
12971 => "111011001000001110000100",
12972 => "110101000011000000111001",
12973 => "110000101111001000101110",
12974 => "101110000001011010010000",
12975 => "101100101111110000100000",
12976 => "101110000001000011010110",
12977 => "110001110100100110011010",
12978 => "110101001010010111000110",
12979 => "110110010000100111010100",
12980 => "110110011001111010111110",
12981 => "110110111110010010000110",
12982 => "110111010001000110110010",
12983 => "110110011010000011111000",
12984 => "110101100000011000100111",
12985 => "110101001000001010001110",
12986 => "110100011001011011110100",
12987 => "110011001100000110010000",
12988 => "110010001110111011100110",
12989 => "110010000111111001011100",
12990 => "110010001001101001101100",
12991 => "110001011110001100000010",
12992 => "110000101110000011000010",
12993 => "110000101110101100100000",
12994 => "110001110011011011100010",
12995 => "110010110110000110011010",
12996 => "110010011101111000001110",
12997 => "110001011110111011100100",
12998 => "110000011100010001011100",
12999 => "101110111010100001001110",
13000 => "101101110011010010010100",
13001 => "101110001100100101010110",
13002 => "110000001111100000000110",
13003 => "110011010111010111111110",
13004 => "110111001001010101001101",
13005 => "111011101010110011101000",
13006 => "000000100101000010111100",
13007 => "000101001000011000110010",
13008 => "001000001101110011010011",
13009 => "001001110001100000110000",
13010 => "001011101111101110110010",
13011 => "001111000111001100111000",
13012 => "010010111010100010100100",
13013 => "010101110011111101010000",
13014 => "010111110010100001110000",
13015 => "011010000000100101110011",
13016 => "011011111110000001010101",
13017 => "011100111111100011001101",
13018 => "011101100000111010101101",
13019 => "011101000111101111011100",
13020 => "011100010100001011001011",
13021 => "011011110110110101001100",
13022 => "011011001001111011111011",
13023 => "011010011101010001110000",
13024 => "011001110111110011000011",
13025 => "011001001000100111101111",
13026 => "011000110001110000011100",
13027 => "011000011111000110100101",
13028 => "011000000110101101000101",
13029 => "011000001100110110110011",
13030 => "010111000110000110010010",
13031 => "010010001011010100110010",
13032 => "001010000110011011110110",
13033 => "000001011111110000011101",
13034 => "111010001001100001100111",
13035 => "110100010110011011111011",
13036 => "101101101010111001100110",
13037 => "100101111010000011001011",
13038 => "100001110110010000110000",
13039 => "100001110001110000011111",
13040 => "100001111100100010111111",
13041 => "100010001001001101101011",
13042 => "100011000100101000111011",
13043 => "100110010000001011101111",
13044 => "101100010000110011110000",
13045 => "110001010101111011100010",
13046 => "110101000110110110000111",
13047 => "111010010110000110000000",
13048 => "111111110000101100100111",
13049 => "000011111001000000110110",
13050 => "000110111110100101011001",
13051 => "000111111001110100101001",
13052 => "000111000111001000010010",
13053 => "000110111100101000100000",
13054 => "000110100010001111011010",
13055 => "000100000100011110001110",
13056 => "000001100100101101100001",
13057 => "000000100001100000011101",
13058 => "111111110011010000101010",
13059 => "111111000000011001010010",
13060 => "111101111000100100101100",
13061 => "111100010011110001100001",
13062 => "111010010111110000011111",
13063 => "110111101101101110000001",
13064 => "110101011100001110001010",
13065 => "110100101100101010111100",
13066 => "110100010101110111010111",
13067 => "110011101011010111000000",
13068 => "110100111101101011010011",
13069 => "111000111110000011010000",
13070 => "111011011101011001000010",
13071 => "111011011010011011100000",
13072 => "111101011001010010010010",
13073 => "000010001001100011001000",
13074 => "000111010000000100001111",
13075 => "001011011001000010010110",
13076 => "001101101000011100110100",
13077 => "001110011111001100001000",
13078 => "001101100100011101010100",
13079 => "001001100000010001101101",
13080 => "000100100000110000001110",
13081 => "000001011001000000010001",
13082 => "111111010110010000010001",
13083 => "111101010011010001101110",
13084 => "111100010001001101001110",
13085 => "111100011000011111110011",
13086 => "111100101011001101101000",
13087 => "111101100101010010001101",
13088 => "111111000011011101011101",
13089 => "000000100001101001101110",
13090 => "000010010111001000101000",
13091 => "000011110010111111100010",
13092 => "000100010010111011001001",
13093 => "000100011000111111111000",
13094 => "000011110101011101111111",
13095 => "000010111011011010100011",
13096 => "000010101101001101001110",
13097 => "000011011111010101101101",
13098 => "000100001110010101010110",
13099 => "000100000000110010111100",
13100 => "000100010110010110011110",
13101 => "000110001000101100001111",
13102 => "000111111101000110101011",
13103 => "001000001010001110001010",
13104 => "000101101101101101110101",
13105 => "000001111011100001011100",
13106 => "111110111011110100001101",
13107 => "111100100100101001001110",
13108 => "111010001100111101100011",
13109 => "111000001011111011110001",
13110 => "110111100010101001101000",
13111 => "111000110001010110111011",
13112 => "111011100001001110001010",
13113 => "111111100100111101110110",
13114 => "000011101111101011110111",
13115 => "000110100101110000001100",
13116 => "001000000011111101001000",
13117 => "000111111111110111011100",
13118 => "000101110100001001010100",
13119 => "000000111011100010100101",
13120 => "111001100010011100111010",
13121 => "110000111101000111110000",
13122 => "101001000011010101110110",
13123 => "100100110101100011010011",
13124 => "100101000101001001011101",
13125 => "100110011000110111011100",
13126 => "100110101010111000110001",
13127 => "100111000011000000001010",
13128 => "101000001001111101001100",
13129 => "101000100111111111110100",
13130 => "101001010101111001011000",
13131 => "101110010100100110111000",
13132 => "110110100101100000110101",
13133 => "111101100100011011111110",
13134 => "000011000011001101000101",
13135 => "000111011101001001010110",
13136 => "001001001000001111001100",
13137 => "000111110001000010110001",
13138 => "000100101000111001100111",
13139 => "000001101000011011111100",
13140 => "000000001011011011110110",
13141 => "000000100101100010100111",
13142 => "000011000001000010000101",
13143 => "000111111011110000001111",
13144 => "001110011001111001010010",
13145 => "010100000111100100100110",
13146 => "011000111001100000100011",
13147 => "011100111110111011100111",
13148 => "011110100101100100110011",
13149 => "011101111101010011111011",
13150 => "011100111001010110110011",
13151 => "011011111101010000011001",
13152 => "011011011010001100000011",
13153 => "011010111010101100000010",
13154 => "011010000100100010111100",
13155 => "011000111111000111000010",
13156 => "010111111101011001100110",
13157 => "010111100111010001000000",
13158 => "010111101001011010100010",
13159 => "010111001111100110110100",
13160 => "010110100000111001010100",
13161 => "010110000011001110001010",
13162 => "010100010001010010000000",
13163 => "001101011010111110010100",
13164 => "000011001101000101010111",
13165 => "111011010111000011011010",
13166 => "110101111101100010011101",
13167 => "110001000110010010100000",
13168 => "101101001010111001011000",
13169 => "101001111010011100111010",
13170 => "100111101001001111111111",
13171 => "100110101100110000000011",
13172 => "100110011111010000011101",
13173 => "100111010111110001010111",
13174 => "101000010100100010110100",
13175 => "100110110011001101000111",
13176 => "100011110101111110101001",
13177 => "100010110111101001101101",
13178 => "100011100000110100011100",
13179 => "100011101010011111110101",
13180 => "100011111011011010110111",
13181 => "100101000010000100111001",
13182 => "100111000011111111001111",
13183 => "101001011101001000100100",
13184 => "101010011011100011110100",
13185 => "101010111100001110101000",
13186 => "101100101001110110111010",
13187 => "101110000010100010100010",
13188 => "101110011011111100000000",
13189 => "101111011111100010111100",
13190 => "110010011001110011011110",
13191 => "110110101010001001101001",
13192 => "111010111000111011111110",
13193 => "111110001011100100111100",
13194 => "000000111101111001100000",
13195 => "000110010110110101010101",
13196 => "001110111010101111001100",
13197 => "010101101000010111000100",
13198 => "011001001001010101111010",
13199 => "011100010010001100000011",
13200 => "011110100010101000001000",
13201 => "011110110000000111011100",
13202 => "011110001000111101111011",
13203 => "011101110100100010011000",
13204 => "011100101110101001110100",
13205 => "011001000001011100101111",
13206 => "010011111000011000010000",
13207 => "001111111110110010011100",
13208 => "001100100101111111000010",
13209 => "000111001111001011000101",
13210 => "000001111101011011011101",
13211 => "000001001101110101100110",
13212 => "000011111101011110011100",
13213 => "000110100111110101010001",
13214 => "001000101110000110011011",
13215 => "001010010001101001110100",
13216 => "001010011000011101110110",
13217 => "001000000110000101000110",
13218 => "000100010101100001001010",
13219 => "000001111010010010010111",
13220 => "000001011111010010100011",
13221 => "000010000010001000011000",
13222 => "000010010001000000000010",
13223 => "000000110110001111010011",
13224 => "111110101101100010010101",
13225 => "111101001110100101110001",
13226 => "111100010000011010010111",
13227 => "111011100110111010011111",
13228 => "111011001001000011000010",
13229 => "111010111001110101111101",
13230 => "111010100001001001101001",
13231 => "111001000100000011001011",
13232 => "110110000001111011000110",
13233 => "110001001111101010111010",
13234 => "101011110111000111101110",
13235 => "100111111110001010101011",
13236 => "100110111000110010011011",
13237 => "101000001001100001110100",
13238 => "101010000110000000000010",
13239 => "101101000000111011010000",
13240 => "110001011000100010111100",
13241 => "110101010010100101100101",
13242 => "111000010110110101110000",
13243 => "111011110111011101011010",
13244 => "111111111110010000000001",
13245 => "000011110000110111001010",
13246 => "000110001011000111000011",
13247 => "000111011001101000011010",
13248 => "000111111000101010111001",
13249 => "000111101111001110000010",
13250 => "000110111110010111000011",
13251 => "000100101100000010011100",
13252 => "000001101100110010111100",
13253 => "111111111101101110110010",
13254 => "111110110001010100000111",
13255 => "111100011111001011101101",
13256 => "111000011101100011100010",
13257 => "110011001110111001100010",
13258 => "101110001000111100000100",
13259 => "101010001101100100110110",
13260 => "101000101000101011000010",
13261 => "101001101100111000011000",
13262 => "101100101100001001101010",
13263 => "110001011110010110001100",
13264 => "110111100110110101101111",
13265 => "111110000000100001101001",
13266 => "000011011010111010011011",
13267 => "000110111000011100000010",
13268 => "001000100001101010010110",
13269 => "001001100011001101011101",
13270 => "001011001010110110001010",
13271 => "001100000100001000100100",
13272 => "001010110011011110010110",
13273 => "001001001001101110010110",
13274 => "000111010110010101111100",
13275 => "000100000001000001111011",
13276 => "000000011000101011011001",
13277 => "111110011000100011010011",
13278 => "111110101111101100111101",
13279 => "000001000001000111010000",
13280 => "000100111111011010010101",
13281 => "001011001101010001101101",
13282 => "010010010111010101111010",
13283 => "011000011101101000001011",
13284 => "011100010000010011100010",
13285 => "011100111011101111011000",
13286 => "011011110101000111100100",
13287 => "011010111010110110110011",
13288 => "011010010111000011100101",
13289 => "011001101110101000010101",
13290 => "011001100110000001001011",
13291 => "011001001011101101000101",
13292 => "010100110100110110100000",
13293 => "001100111000000010011000",
13294 => "000110110001111111001001",
13295 => "000100001001110001001011",
13296 => "000010111111111000011110",
13297 => "000010010000111000111010",
13298 => "000001111001000000101101",
13299 => "000010101111001100011100",
13300 => "000100011011011101011011",
13301 => "000101010000000100110001",
13302 => "000101000100110001110110",
13303 => "000100101101100110011000",
13304 => "000011111001110000011111",
13305 => "000001110100101001001000",
13306 => "111110011111001011000011",
13307 => "111001110010010100010001",
13308 => "110011100111000010010110",
13309 => "101101101001101001100100",
13310 => "101001101110001110100100",
13311 => "100111101011000010100100",
13312 => "100101011101000100000010",
13313 => "100010101100110000100111",
13314 => "100010010011010010001111",
13315 => "100011101111100110111101",
13316 => "100100010011000100011001",
13317 => "100100111001001010101000",
13318 => "100101100111101100111001",
13319 => "100101110111010111000001",
13320 => "100110011111011100101001",
13321 => "100110100110011111001001",
13322 => "100110011101011000101101",
13323 => "100111001100000110101111",
13324 => "100111010111001000111100",
13325 => "101000000000100000001010",
13326 => "101100010101101100110110",
13327 => "110011001001100001001010",
13328 => "111001011110001010100111",
13329 => "111111101001010000101100",
13330 => "000101101000101011010010",
13331 => "001001010100001111110110",
13332 => "001010111010110000100011",
13333 => "001100100010001101001010",
13334 => "001111011101001110010000",
13335 => "010011000000101101001000",
13336 => "010100100101111100001110",
13337 => "010011111010001010111000",
13338 => "010010001001111011101000",
13339 => "001111101011001111010000",
13340 => "001111001010100001010100",
13341 => "010001101011001000010000",
13342 => "010011110111010110010100",
13343 => "010100110011001010011110",
13344 => "010110010110010101010110",
13345 => "011000100010001110111001",
13346 => "011001100100111001010001",
13347 => "011000111001110100000001",
13348 => "011000001111010010000001",
13349 => "011001000000001100110111",
13350 => "011010100001101101010001",
13351 => "011011000101101011110001",
13352 => "011010011000011111100001",
13353 => "011001100100110101110111",
13354 => "011001000011111001011111",
13355 => "011000110100110001101111",
13356 => "010111101111010100001110",
13357 => "010100011000001111111000",
13358 => "010000010000010011100010",
13359 => "001100010000000100000000",
13360 => "000111011011110111111110",
13361 => "000010011110011110110110",
13362 => "111101101010111011000110",
13363 => "111000100110110110110001",
13364 => "110011110010011110101000",
13365 => "101111110101100010110110",
13366 => "101100100110010100100010",
13367 => "101000100010011110010000",
13368 => "100011110110101101010101",
13369 => "100001001111100111000010",
13370 => "100000111101001111110111",
13371 => "100001000000101110111110",
13372 => "100000110010011001101111",
13373 => "100000111101111111011100",
13374 => "100001011110100011001011",
13375 => "100001111100010111011001",
13376 => "100100001110101010100001",
13377 => "101010000101111011001010",
13378 => "110001101001100010101110",
13379 => "110111100000001110010111",
13380 => "111010101010110110111001",
13381 => "111101000101010111100111",
13382 => "111111111110001010010100",
13383 => "000010011010001100110111",
13384 => "000010111111010011101101",
13385 => "000000101000001101010001",
13386 => "111100011101001001000011",
13387 => "111001000010110011101010",
13388 => "110111101100001110110100",
13389 => "111000010000100111100011",
13390 => "111001011010100010101110",
13391 => "111011001010010000001111",
13392 => "111110100010111111011011",
13393 => "000010001100011000000000",
13394 => "000100110100111100101011",
13395 => "000110010010110100010110",
13396 => "000110001010111100100010",
13397 => "000101010110101001011010",
13398 => "000100110100001111011111",
13399 => "000101001000100010100110",
13400 => "000111000011011111101110",
13401 => "001001110011000100001110",
13402 => "001100010000001001000100",
13403 => "001110011010010001100100",
13404 => "010000100000010110011100",
13405 => "010010001101111100001010",
13406 => "010011000010000111111100",
13407 => "010011011000110011110010",
13408 => "010011010101000111010000",
13409 => "010010001011000111011100",
13410 => "010000001010111101101000",
13411 => "001101110001001011011010",
13412 => "001011011010011000001100",
13413 => "001001101010001000001001",
13414 => "001000100101010010110110",
13415 => "001000001110101101110000",
13416 => "001000100110010111111100",
13417 => "001001110000110101101000",
13418 => "001011100110101010001011",
13419 => "001101100100011110011000",
13420 => "001110110100100001001000",
13421 => "001101110010010011110110",
13422 => "001001110101101110011101",
13423 => "000011111000110011110011",
13424 => "111101011111100111001111",
13425 => "111000100010101101010111",
13426 => "110100001101010101110000",
13427 => "101110111111010100011000",
13428 => "101011000010110011110010",
13429 => "101010001111010001000000",
13430 => "101100001011100010001110",
13431 => "110000000111000011011000",
13432 => "110101000001100110100000",
13433 => "111010110001010001110101",
13434 => "000001101100111111100010",
13435 => "001001011011011111011101",
13436 => "001111111010100101101100",
13437 => "010010100100011110110110",
13438 => "010010000010101010111100",
13439 => "010000000010100010010000",
13440 => "001100000011011111100110",
13441 => "000110011001011101111101",
13442 => "000000110100111001011000",
13443 => "111100000111111101011001",
13444 => "110111101110011101011000",
13445 => "110011011011010100111010",
13446 => "101111110000001111000110",
13447 => "101011101101001111001110",
13448 => "100110111100100001110001",
13449 => "100100101010111101011100",
13450 => "100101111011101000000111",
13451 => "100110010110101001111111",
13452 => "100100010100101110101101",
13453 => "100011111010001011110011",
13454 => "100101100101101001100100",
13455 => "100110010101011100000100",
13456 => "100110100010010000001100",
13457 => "100110101110101100101100",
13458 => "100111100001000011101111",
13459 => "101010110100111100100110",
13460 => "101110100011001010101110",
13461 => "110000100111010111010000",
13462 => "110011000111111111101100",
13463 => "110111000000000010111010",
13464 => "111011001010100001001100",
13465 => "111101110001001110111001",
13466 => "111101111101100100001111",
13467 => "111110000001111000001000",
13468 => "111110111000101100110111",
13469 => "111110101000110000110101",
13470 => "111101100000100011111000",
13471 => "111101101011100100001101",
13472 => "111111110110101110001010",
13473 => "000011011101110010001101",
13474 => "000111001010001011100111",
13475 => "001001001011000010011000",
13476 => "001010010110011101001010",
13477 => "001100010010010011000010",
13478 => "001101110100010100001010",
13479 => "001110110111100110101100",
13480 => "010000101111010010101110",
13481 => "010010101100001100110110",
13482 => "010011011110011111001110",
13483 => "010010011011011111101100",
13484 => "001111111110000011100100",
13485 => "001101001001010001001000",
13486 => "001010000101011111001100",
13487 => "000111100100011011110111",
13488 => "000110011001111111000011",
13489 => "000101111011111011011001",
13490 => "000101101000011000110011",
13491 => "000101110111000101100111",
13492 => "000111001110000001111110",
13493 => "001000010010011001100010",
13494 => "000110110000100101111011",
13495 => "000011110111011011010101",
13496 => "000010010001101111111100",
13497 => "000001111110110100011101",
13498 => "000001010001100000111111",
13499 => "111111100010001011000000",
13500 => "111101101111001101010000",
13501 => "111100001111101000111100",
13502 => "111011000000111110010100",
13503 => "111010110100101100110101",
13504 => "111011100110000110011111",
13505 => "111100000100011110111001",
13506 => "111011100100111110111101",
13507 => "111010111110111100110000",
13508 => "111010101000101000111000",
13509 => "111001011000111110111100",
13510 => "110111101100000001101010",
13511 => "110110110011010001101011",
13512 => "110110011100001000000011",
13513 => "110110001100001101011110",
13514 => "110110001100010111101010",
13515 => "110111001010011100100111",
13516 => "111001011101100100000011",
13517 => "111100001111001001110100",
13518 => "111110011101111010110000",
13519 => "111110100100111110010101",
13520 => "111100100001100100110001",
13521 => "111011000111101010111001",
13522 => "111011000001001110000011",
13523 => "111010100100100010001111",
13524 => "111010010111011100111100",
13525 => "111100000010111101110011",
13526 => "111111000011100010101001",
13527 => "000001110100001001000110",
13528 => "000011111100100101010001",
13529 => "000101010010010110101111",
13530 => "000110011000000100101011",
13531 => "001001000010101101100101",
13532 => "001100110111001101101000",
13533 => "001111110111001111101010",
13534 => "010001101100100110100000",
13535 => "010010011010001111110110",
13536 => "010001111010101010001110",
13537 => "010000000000001111001000",
13538 => "001100001111000101111110",
13539 => "000111110110010011100100",
13540 => "000101011010010101001110",
13541 => "000101101011000001100001",
13542 => "000110110001011011101110",
13543 => "000111010101110001010101",
13544 => "000111100011000100100100",
13545 => "000111100000100001000010",
13546 => "000111111110100001110000",
13547 => "001001100000111100000000",
13548 => "001011001010101111100110",
13549 => "001100001110011001111100",
13550 => "001011111000101000111001",
13551 => "001001001101111001010110",
13552 => "000100101010110011100010",
13553 => "111111010011101110100101",
13554 => "111010001111000011000101",
13555 => "110101111111001111101001",
13556 => "110010100110111100100010",
13557 => "110000101100000110010110",
13558 => "110000011000111100000000",
13559 => "110001001110010111001100",
13560 => "110010110101100011010000",
13561 => "110100101101101011011110",
13562 => "110110010111101111010100",
13563 => "111000000001000001010111",
13564 => "111010110000000111011011",
13565 => "111110110011011010000111",
13566 => "000010111011101100101101",
13567 => "000110100000101101111101",
13568 => "001001010011111010110111",
13569 => "001011101010100000010000",
13570 => "001110101111000111011100",
13571 => "010001111101001000000100",
13572 => "010100000000000000000110",
13573 => "010101000011100101110110",
13574 => "010101001000110110100100",
13575 => "010011001110111101100100",
13576 => "001110011100001001111110",
13577 => "000110111110110101101111",
13578 => "111110011101010000110100",
13579 => "110110110101111011111011",
13580 => "110000101110011010100100",
13581 => "101011100011010110101010",
13582 => "101000001011011001111010",
13583 => "100111100000001111111011",
13584 => "101000101010101101101100",
13585 => "101011110011010110000110",
13586 => "110001000110000000000100",
13587 => "110110110100111001000010",
13588 => "111100001111000101111101",
13589 => "000001010110000110000110",
13590 => "000100001100100010111101",
13591 => "000010000101110111110101",
13592 => "111011011011000000101111",
13593 => "110011111110001101001110",
13594 => "101110101100011111100010",
13595 => "101011110000101100000100",
13596 => "101001111110010110000000",
13597 => "101000101111010001001000",
13598 => "101000110100000100010100",
13599 => "101010000100001100101100",
13600 => "101011101010010100101110",
13601 => "101110101110100010111110",
13602 => "110100110011010100111100",
13603 => "111100111110000001001111",
13604 => "000100011100011100010111",
13605 => "001010000100011001100001",
13606 => "001111000011001101110010",
13607 => "010011011011010110000010",
13608 => "010101110001111000001000",
13609 => "010101101100110001100110",
13610 => "010100101110101011001100",
13611 => "010100111111011010111010",
13612 => "010101111110100001010010",
13613 => "010101101110000001001010",
13614 => "010011111111001001001100",
13615 => "010001010110010010100000",
13616 => "001110101011001110110110",
13617 => "001100110010101000111010",
13618 => "001011001010011110100110",
13619 => "001001000000110001010000",
13620 => "000110001111011011001010",
13621 => "000011000101100000110001",
13622 => "000000001011001011111110",
13623 => "111101110111010010011100",
13624 => "111011000110101100001110",
13625 => "110111000001001000011010",
13626 => "110011011010110100010000",
13627 => "110010011001111001001110",
13628 => "110011010010101010111110",
13629 => "110100011011011101100110",
13630 => "110101100111001111110000",
13631 => "110111100111101110100100",
13632 => "111001110001011000100110",
13633 => "111010110100101010110100",
13634 => "111011011010010011011110",
13635 => "111011110000100001111101",
13636 => "111011101111110010110111",
13637 => "111100010100000011010100",
13638 => "111100011110000110110010",
13639 => "111010110100101111100110",
13640 => "111000011001111001100001",
13641 => "110110011000110110001110",
13642 => "110101000010011110100010",
13643 => "110100000001000011111001",
13644 => "110010111111001100110110",
13645 => "110001110110011100111010",
13646 => "101111110110000110111000",
13647 => "101101010011011000011010",
13648 => "101011111101011101100110",
13649 => "101100000100100011111100",
13650 => "101101001010011010001100",
13651 => "110000000010111001111010",
13652 => "110101001010100010000011",
13653 => "111011010001111110101001",
13654 => "000001100011010001100001",
13655 => "001000110101000101001010",
13656 => "010001000110100000101000",
13657 => "010111101010011100000110",
13658 => "011010101110111111100111",
13659 => "011100011101100001011011",
13660 => "011110001010111101000000",
13661 => "011110000111110100010111",
13662 => "011100101111011000111101",
13663 => "011100000000101010110111",
13664 => "011011110100100100100010",
13665 => "011011101000001011010101",
13666 => "011011001101011111001001",
13667 => "011010101011000111100110",
13668 => "011001111111011111001011",
13669 => "011000100000000111011111",
13670 => "010111011000110100110110",
13671 => "010111001011011000010110",
13672 => "010100110011101101011100",
13673 => "001111010101101110111000",
13674 => "001001010101101000001011",
13675 => "000100000010001001100111",
13676 => "111111101011111011100110",
13677 => "111101100010001110101011",
13678 => "111101110111011010111100",
13679 => "111110101011100101000101",
13680 => "111110011110010111001001",
13681 => "111101110011010111010010",
13682 => "111100001101011000001000",
13683 => "110111111010010100110010",
13684 => "110001111010011000101110",
13685 => "101101100111101010100110",
13686 => "101011110111111000011110",
13687 => "101010100110000011000010",
13688 => "101000110011110010000010",
13689 => "100111001100000110101110",
13690 => "100101101011111101110110",
13691 => "100011110111000110101111",
13692 => "100011001101111101001100",
13693 => "100101100010111011000101",
13694 => "101001001010111101110110",
13695 => "101100001100100100010010",
13696 => "110000001101100110100010",
13697 => "110101100100111110111111",
13698 => "111001011100101101001110",
13699 => "111010111001101100111000",
13700 => "111100000000100000101111",
13701 => "111101101010000000000000",
13702 => "111110111100110110001110",
13703 => "000000110111111110001101",
13704 => "000100110111101111101100",
13705 => "001000101011111101011101",
13706 => "001010000000011100100011",
13707 => "001010000000111010001000",
13708 => "001001100010100010100010",
13709 => "000111110110100010000010",
13710 => "000110010101010000011111",
13711 => "000111100000001110011011",
13712 => "001001101101010111111110",
13713 => "001001000101000100111101",
13714 => "000110011001000101101100",
13715 => "000100101001010010111101",
13716 => "000011111000001011000110",
13717 => "000011010101011001001110",
13718 => "000010111011000110000000",
13719 => "000011001011011000000110",
13720 => "000101110100010111001001",
13721 => "001010011110100101111000",
13722 => "001110001101101010010000",
13723 => "001111011000101000110010",
13724 => "001110000110110111110100",
13725 => "001100011100100101001010",
13726 => "001100011011110010011000",
13727 => "001011000011001011011011",
13728 => "000101000010101100011011",
13729 => "111100000011100100110100",
13730 => "110001001111100100101110",
13731 => "100110111010000001110111",
13732 => "100010100001110101100101",
13733 => "100011010000011101010001",
13734 => "100100000101001000011100",
13735 => "100100110101000000000011",
13736 => "100101111011000110000011",
13737 => "100111110111000000000110",
13738 => "101101110100000001111010",
13739 => "110111000011101001001111",
13740 => "000000001000011000111000",
13741 => "001000111001101100000110",
13742 => "010000101010001010101110",
13743 => "010101010000111011011010",
13744 => "010111001011100110101010",
13745 => "010111001001000100110100",
13746 => "010100100101100001100010",
13747 => "010000011010111100010000",
13748 => "001100100000100101111100",
13749 => "001001011011000111100010",
13750 => "000110111101100010001100",
13751 => "000101011010001001000100",
13752 => "000100110101010110011111",
13753 => "000100001010000100000011",
13754 => "000011001010010100010100",
13755 => "000011010001001000000010",
13756 => "000100001010010010101011",
13757 => "000100000010110010000001",
13758 => "000010110100010100100101",
13759 => "000000100011001001000010",
13760 => "111100111000111101100011",
13761 => "111001010011011111111100",
13762 => "110110111010101111000100",
13763 => "110100011101011011111000",
13764 => "110001000111111011010110",
13765 => "101110100101010000101100",
13766 => "101110110111110001011000",
13767 => "110001011011110011000010",
13768 => "110100001100110100101101",
13769 => "110110101101010110000011",
13770 => "111001000000000101000001",
13771 => "111001100111001000010101",
13772 => "111000000000110111111011",
13773 => "110110000110110011101010",
13774 => "110100111101010010101000",
13775 => "110011101000011011011010",
13776 => "110001110111010001010000",
13777 => "101111110111111110000110",
13778 => "101100111111101010110110",
13779 => "101001111011100111110000",
13780 => "101000101111010100001100",
13781 => "101001000001100000100010",
13782 => "101001001110100110010110",
13783 => "101010011101101010111000",
13784 => "101101111000110100001010",
13785 => "110001111001100100111110",
13786 => "110101000100110011011001",
13787 => "110111101000100000100101",
13788 => "111001110111111011001101",
13789 => "111011110010000011000011",
13790 => "111101101001111100011011",
13791 => "000000101001101111011010",
13792 => "000101100001111000001010",
13793 => "001011110111110011110000",
13794 => "010011011100000000010110",
13795 => "011010100001101111101011",
13796 => "011101111101111001100011",
13797 => "011110001010101100111111",
13798 => "011110000001000000100101",
13799 => "011101111000001100011111",
13800 => "011101000110000001111011",
13801 => "011100000101111100100110",
13802 => "011011010110000111011101",
13803 => "011011000010000010101101",
13804 => "011011000000011011001101",
13805 => "011010111110100001110000",
13806 => "011010110001000110010011",
13807 => "011010010100001000000001",
13808 => "011010000100110011110010",
13809 => "011010000111100100010011",
13810 => "011010000010001100001111",
13811 => "011010010100111100110101",
13812 => "011001111100101111000001",
13813 => "010101110100100100000000",
13814 => "001110010010111110101000",
13815 => "000110010110001001101010",
13816 => "111110101100001010110010",
13817 => "110111100000111000111010",
13818 => "110001100000000111011010",
13819 => "101100001011000010111100",
13820 => "100111101010011101110101",
13821 => "100101000100100011011001",
13822 => "100100011011000110010101",
13823 => "100100110101111011111111",
13824 => "100101001110001111011100",
13825 => "100101001111010110010111",
13826 => "100101100111010110101011",
13827 => "100101111111011001100001",
13828 => "100101110101010010111101",
13829 => "100110100001100110111111",
13830 => "101000001100111011001100",
13831 => "101000110010010000010010",
13832 => "101000100100000110011100",
13833 => "101001110001111001010110",
13834 => "101100100000111011101010",
13835 => "101111101010011000101100",
13836 => "110010111111010100110010",
13837 => "110110101000000010111001",
13838 => "111010101011000100100101",
13839 => "111110001010110110011001",
13840 => "111111100000110010000011",
13841 => "111111100101000110000110",
13842 => "000000001101110010001110",
13843 => "000000101101101001011100",
13844 => "000000110001010011010110",
13845 => "000001111111101001000000",
13846 => "000100011100111111010001",
13847 => "000111110010110101001010",
13848 => "001100101011010001110100",
13849 => "010001101111011111101100",
13850 => "010101010000011001000110",
13851 => "011000100000001000010111",
13852 => "011100010010111110100101",
13853 => "011110011011100011101001",
13854 => "011101110010011101011011",
13855 => "011100100000111101011011",
13856 => "011100100000110111011001",
13857 => "011101000111100011011001",
13858 => "011100011101011101100100",
13859 => "011001101110011001100101",
13860 => "010110010001100010010110",
13861 => "010011000101100010010000",
13862 => "001111000111000001000100",
13863 => "001011000011011010001100",
13864 => "001000101010101011101100",
13865 => "000110010111011110000000",
13866 => "000010011010010011011001",
13867 => "111100111101110110000111",
13868 => "110101110100000110100111",
13869 => "101110110010000101101100",
13870 => "101010111100111010011110",
13871 => "101010000000010100000010",
13872 => "101010101010010100001010",
13873 => "101100111000011110000010",
13874 => "110000001110111010000100",
13875 => "110100100100101011010001",
13876 => "111001001001100101011101",
13877 => "111100000111100101111011",
13878 => "111110001100110111111001",
13879 => "000001100010100010100110",
13880 => "000100111001001101110000",
13881 => "000101010110111000110111",
13882 => "000010101011000010010101",
13883 => "111110100001110011010101",
13884 => "111010010100010101011101",
13885 => "110111000101010010010001",
13886 => "110100111110110101110001",
13887 => "110011001111101100010010",
13888 => "110010011101000011110000",
13889 => "110100001001001001110000",
13890 => "110111100110110110001010",
13891 => "111010010110011110011111",
13892 => "111011100001000000111011",
13893 => "111100101110001111011000",
13894 => "111110111111100001001001",
13895 => "000000101110010110001010",
13896 => "000000100010100011110110",
13897 => "111111010010110001001100",
13898 => "111101111011110010010111",
13899 => "111100100001001001010101",
13900 => "111011001101000100110110",
13901 => "111010010110101110100001",
13902 => "111001111100110010010011",
13903 => "111001110100000100001110",
13904 => "111010101101100111100100",
13905 => "111101011001101011111111",
13906 => "000000101011100000010000",
13907 => "000010111101110110101011",
13908 => "000100001010001101100101",
13909 => "000100100011001110110011",
13910 => "000011111011001001010100",
13911 => "000001110010100100000101",
13912 => "111110101011100011110100",
13913 => "111100110100000001000001",
13914 => "111100110111100111011100",
13915 => "111100011111000010010110",
13916 => "111010100110010000111010",
13917 => "111001000011111101111100",
13918 => "111000110010100010000111",
13919 => "111000111111000011110101",
13920 => "111001100101111001101100",
13921 => "111010100011001000011100",
13922 => "111010110110111111000110",
13923 => "111010100100110111110101",
13924 => "111010101010010000001111",
13925 => "111011000010011110101010",
13926 => "111011010110011010000110",
13927 => "111100011010001100110100",
13928 => "111111011001101101011010",
13929 => "000011110010101001110010",
13930 => "000111101010101011001000",
13931 => "001010101000100111101011",
13932 => "001101100011000101100000",
13933 => "010000100000100011000000",
13934 => "010011011011110111111010",
13935 => "010101110110111101010100",
13936 => "010111001110110111001000",
13937 => "011000011111110110000111",
13938 => "011001110111110111001011",
13939 => "011010000110000101100111",
13940 => "011001001100011000110001",
13941 => "010111100010101111010000",
13942 => "010101001011101001100100",
13943 => "010011000010110010010100",
13944 => "010000011111010100111100",
13945 => "001011101100111001011100",
13946 => "000110000000001101111010",
13947 => "000001110111010110010100",
13948 => "111110110011100101101101",
13949 => "111011000011100101001000",
13950 => "110110000010010101111111",
13951 => "110000111111010101101000",
13952 => "101110001011010010011010",
13953 => "101101111000001110001010",
13954 => "101110100011100011100010",
13955 => "110000001000101110111110",
13956 => "110011000010110000001110",
13957 => "110110011101011100000111",
13958 => "111001101101001000101101",
13959 => "111100000010101000100010",
13960 => "111100101011111000100110",
13961 => "111100001110001011010101",
13962 => "111011110001100100111111",
13963 => "111011111001001011110110",
13964 => "111100000101101111010000",
13965 => "111011011101111111111101",
13966 => "111010101000001000100010",
13967 => "111010000010000110111011",
13968 => "111000110000001101111100",
13969 => "110111000011010011011111",
13970 => "110101010101100011001000",
13971 => "110010111010001000000100",
13972 => "110001001010011100101100",
13973 => "110010011000100111010000",
13974 => "110101011011101101100001",
13975 => "110111010011111110000010",
13976 => "110111011000011010011111",
13977 => "110111001001101111100000",
13978 => "110111001110000011011011",
13979 => "110111011000010101101000",
13980 => "111000011010110000100000",
13981 => "111011011101101100010011",
13982 => "000000101100101010010110",
13983 => "000110011010101101110000",
13984 => "001010101000110001111000",
13985 => "001101110100111001111000",
13986 => "010000101110010000100000",
13987 => "010011011011010110101010",
13988 => "010111000001101010000010",
13989 => "011010010000110110111110",
13990 => "011010110011010110111111",
13991 => "011010001001110101110010",
13992 => "011001001010000000110000",
13993 => "010101111011100101110110",
13994 => "010001001010001001100000",
13995 => "001100110011101001110100",
13996 => "001001001100100110011100",
13997 => "000110100110100101010110",
13998 => "000101010101110101101100",
13999 => "000101000110111001110100",
14000 => "000101001001001010001110",
14001 => "000100001011001110101010",
14002 => "000001101101011000111101",
14003 => "111111100001100001110110",
14004 => "111111011110101111000000",
14005 => "111111011001001110011100",
14006 => "111011100001100011000010",
14007 => "110100111110111111100011",
14008 => "101111111010010010110000",
14009 => "101110000011010101111110",
14010 => "101110111000110011001100",
14011 => "110000111010100111101000",
14012 => "110010011001000000110100",
14013 => "110010111000101110110100",
14014 => "110011001000001000101010",
14015 => "110011100000111101111010",
14016 => "110011111101011000110100",
14017 => "110100101110100000100100",
14018 => "110101100001010010101011",
14019 => "110101000011010111100000",
14020 => "110011111111010111111100",
14021 => "110011111011010000110110",
14022 => "110011110111110000101000",
14023 => "110011011000011111101010",
14024 => "110100010100100010011010",
14025 => "110111010000001110101011",
14026 => "111011100111010100111100",
14027 => "000001001011001011111100",
14028 => "000111000010111000000001",
14029 => "001011100010110000111100",
14030 => "001101000111101100110100",
14031 => "001100000100010110100000",
14032 => "001010010101111110111100",
14033 => "001000011010001011001111",
14034 => "000100111101110001010011",
14035 => "111111100100110001100100",
14036 => "111001010101000110110101",
14037 => "110011111011011100100000",
14038 => "110000100101010001101110",
14039 => "101110101101000100001110",
14040 => "101100100110011011110110",
14041 => "101011001101111011100110",
14042 => "101101110101101101011110",
14043 => "110100010111010010100110",
14044 => "111011111100111010000101",
14045 => "000011111010010100010110",
14046 => "001011110010111011010010",
14047 => "010001000111111110000100",
14048 => "010010001111100100100000",
14049 => "010000011110011101110100",
14050 => "001110010110101100000110",
14051 => "001011111100101000101101",
14052 => "001000000001100011111100",
14053 => "000100000001101000011000",
14054 => "000001101100101100101001",
14055 => "000000011000010110111111",
14056 => "111111011101100111100011",
14057 => "111111111100101100111100",
14058 => "000011001101101101110001",
14059 => "001000001111100000010111",
14060 => "001011111100010000001110",
14061 => "001101101010010001110010",
14062 => "001110100110101000011100",
14063 => "001110011011001101110010",
14064 => "001101001010010110010000",
14065 => "001100100100111110000000",
14066 => "001101010001001111010010",
14067 => "001101011010011101100110",
14068 => "001100001100110000010110",
14069 => "001011111100001011011010",
14070 => "001101110111100001010010",
14071 => "010000010100101110011000",
14072 => "010010010101110110101100",
14073 => "010011110010110000001000",
14074 => "010100001000001010001110",
14075 => "010010110101111010110100",
14076 => "001111000111001110111100",
14077 => "001000111100001011110111",
14078 => "000001110111101100111110",
14079 => "111011011000011000100101",
14080 => "110110011110010100001001",
14081 => "110010111111001101010110",
14082 => "101111100010100100111100",
14083 => "101100001010111000000110",
14084 => "101010011110101010011000",
14085 => "101010111100010010100110",
14086 => "101100100100011110001100",
14087 => "101110011111111000101010",
14088 => "110000001100101101111000",
14089 => "110001010101101010101000",
14090 => "110010101100000001010100",
14091 => "110100101001111111001101",
14092 => "110101011010001000000110",
14093 => "110011101110101010110100",
14094 => "110001001101110001110000",
14095 => "101111111011011000010000",
14096 => "101111111010111010011010",
14097 => "101111100011001100011010",
14098 => "101110010110101001001110",
14099 => "101101010000110001101010",
14100 => "101100000001100110010010",
14101 => "101010011100110001011100",
14102 => "101001010011000011011100",
14103 => "101000110101111101000110",
14104 => "101001101100100111100100",
14105 => "101011111001110001000010",
14106 => "101110000101101010100010",
14107 => "110000001000000100011010",
14108 => "110010111011011100110110",
14109 => "110111000011111010111100",
14110 => "111100100111101101111101",
14111 => "000010010100010101111001",
14112 => "000111101000111000100001",
14113 => "001110000010011111100010",
14114 => "010100111010100110110100",
14115 => "011001011011110111101010",
14116 => "011010111011110101000111",
14117 => "011011010001101011011111",
14118 => "011011100110111001101011",
14119 => "011011111011101111001001",
14120 => "011100100010001111100111",
14121 => "011100011101000001101111",
14122 => "011010000110110011001111",
14123 => "010110110011001111010110",
14124 => "010100111001000010001000",
14125 => "010101001110001110011000",
14126 => "010111100011001000001010",
14127 => "011001110010110101000001",
14128 => "011010011011000111101001",
14129 => "011010000110010110011111",
14130 => "011000010001011110010011",
14131 => "010100110001010110101010",
14132 => "010001101110111110010000",
14133 => "001110111111111010000100",
14134 => "001011001001101110101010",
14135 => "001000010111010011011000",
14136 => "001000011001011110000010",
14137 => "001000010100111000011000",
14138 => "000101100001100100110000",
14139 => "000001011010011000110010",
14140 => "111101111100110110010110",
14141 => "111011111100000000000011",
14142 => "111011100001110010010010",
14143 => "111010111010111100100000",
14144 => "110111100100111111001101",
14145 => "110000101100001100101100",
14146 => "101000010011110010100000",
14147 => "100010110001011011011110",
14148 => "100001100001111010010101",
14149 => "100001110011111001011001",
14150 => "100001111011010001100011",
14151 => "100001110011010100101011",
14152 => "100001101101111100000111",
14153 => "100010010110001000111011",
14154 => "100011000110010110000001",
14155 => "100100001110010100111111",
14156 => "100110111111001100101100",
14157 => "101010001100100011010000",
14158 => "101101001001011000101100",
14159 => "110001000101101011111110",
14160 => "110101111001000110100101",
14161 => "111010100010000101011011",
14162 => "111101111110101010100000",
14163 => "111111110111110000001000",
14164 => "000001010010011100001110",
14165 => "000010110101101000000110",
14166 => "000100001011101010111000",
14167 => "000100001011000011001001",
14168 => "000010010110011110110010",
14169 => "000000111001110000100010",
14170 => "111111110111000010011111",
14171 => "111100110001010010010010",
14172 => "111001000110001111101110",
14173 => "110111001001101101001101",
14174 => "110110011101100000110010",
14175 => "110111011001010100001100",
14176 => "111010110110110001111110",
14177 => "111111111111011000010110",
14178 => "000100011011011101101101",
14179 => "000111001111011110100111",
14180 => "001011011001000001010100",
14181 => "010001111000110010111000",
14182 => "010110111011010011000110",
14183 => "011001011100111001011001",
14184 => "011011110101110101001101",
14185 => "011101010111100100011011",
14186 => "011011000100011101101011",
14187 => "010101011001001111001000",
14188 => "010000001010000110001010",
14189 => "001100111010000010001100",
14190 => "001010001000110101111010",
14191 => "000111101011100000001100",
14192 => "000110011010010110101111",
14193 => "000101111111101100111101",
14194 => "000101110010011100110110",
14195 => "000110010001101110011111",
14196 => "001001000000111011100111",
14197 => "001110000100000010100100",
14198 => "010011000001010000110000",
14199 => "010110000011101110101010",
14200 => "010111000001111011110110",
14201 => "010110001101100011100000",
14202 => "010011100101100100111100",
14203 => "001110111101110011110100",
14204 => "001001011100000100101010",
14205 => "000100110110010001001101",
14206 => "000001100000111000111011",
14207 => "111110100110101110011000",
14208 => "111011101010110100111110",
14209 => "111001010100001010011110",
14210 => "111000000100011101010001",
14211 => "110110100111011000100101",
14212 => "110011111100110100100010",
14213 => "110001100100110010010100",
14214 => "110000111000110000100000",
14215 => "110001001100100101111010",
14216 => "110001011001110010110010",
14217 => "110001101000101001000110",
14218 => "110010100011110110010110",
14219 => "110011110111110001011010",
14220 => "110100010101001010010001",
14221 => "110011110001101100001110",
14222 => "110011111100001001001010",
14223 => "110100110100100010000001",
14224 => "110100001001110011001001",
14225 => "110010110000110100100100",
14226 => "110010000011110100111000",
14227 => "101111101101001011011100",
14228 => "101011111110011000000010",
14229 => "101001101101110010010110",
14230 => "101000000000010000000010",
14231 => "100110010001010101001101",
14232 => "100110001011111101000110",
14233 => "100111000010010010100001",
14234 => "100111100101010111110001",
14235 => "101000010001101100100110",
14236 => "101001001011111011011000",
14237 => "101001101010111100010100",
14238 => "101001101110001100101000",
14239 => "101001111010001101100000",
14240 => "101001111110111001001010",
14241 => "101010111000111101111010",
14242 => "101111011000010000101100",
14243 => "110110010101110100101110",
14244 => "111100010111010101011110",
14245 => "000001100110000111010111",
14246 => "000110011000100001111101",
14247 => "001001100101110111111111",
14248 => "001011011011110111110000",
14249 => "001100101001100000001010",
14250 => "001110100011010100011100",
14251 => "010010000011001111010000",
14252 => "010101010000011101001100",
14253 => "010110101110100111001100",
14254 => "010111010111000101100100",
14255 => "010111110010100111000110",
14256 => "011000011101011110100010",
14257 => "011010001100001111101100",
14258 => "011100011101100010101101",
14259 => "011101100011000000000100",
14260 => "011101000011101010110101",
14261 => "011100010010010111100001",
14262 => "011011111000111100000100",
14263 => "011011010111011101001010",
14264 => "011010011111010000100100",
14265 => "011001110000111010110101",
14266 => "011001011100101110000001",
14267 => "011001000111110000101011",
14268 => "011000101110111101111101",
14269 => "011000010010111100111001",
14270 => "010111101101110111101110",
14271 => "010111011100010000010100",
14272 => "010110111100101000011010",
14273 => "010110010011011110101110",
14274 => "010110011000101100100000",
14275 => "010011101110010100100100",
14276 => "001100000010010011101110",
14277 => "000100000110100001111110",
14278 => "111110101111101000101101",
14279 => "111010001011101011001011",
14280 => "110011111000001100111100",
14281 => "101010000110011111101000",
14282 => "100001111000111111101000",
14283 => "100000100001000001101111",
14284 => "100001100010100100101001",
14285 => "100001010010110000011001",
14286 => "100001000011000001001010",
14287 => "100000110000000101011001",
14288 => "100001010011010100100111",
14289 => "100010101001001010100100",
14290 => "100011000000010000011001",
14291 => "100011010000001110010001",
14292 => "100011100100110100110001",
14293 => "100101000101001110011011",
14294 => "101011010011011011011010",
14295 => "110011101110110100001100",
14296 => "111001001011010100101100",
14297 => "111011111011011100011100",
14298 => "111101110100110110010001",
14299 => "111110110010000100000110",
14300 => "111101100101110101011111",
14301 => "111010011100011110110111",
14302 => "111000011011111101101101",
14303 => "111001001101110101000100",
14304 => "111011100011011111000011",
14305 => "111101110100101000011011",
14306 => "111110101010000010110010",
14307 => "111111000100000011110001",
14308 => "000001010101110110111100",
14309 => "000101001111000011111000",
14310 => "001001000010001011110110",
14311 => "001011110000011111100110",
14312 => "001110000111101100011000",
14313 => "010001100111100100100110",
14314 => "010101011101101010011010",
14315 => "010111111010100010000110",
14316 => "011000101001011000011001",
14317 => "010111111001000001000010",
14318 => "010111011100000101001110",
14319 => "011001011110111001000111",
14320 => "011100010011111100110010",
14321 => "011100101010010101011010",
14322 => "011011000011011000100000",
14323 => "011010000011010100100011",
14324 => "011001011010101101001101",
14325 => "010110001010100100011100",
14326 => "001111010110111111100110",
14327 => "001000111011011100101110",
14328 => "000110101010111110000110",
14329 => "000110111000001011010110",
14330 => "000110111011010100100010",
14331 => "000111101111011111110011",
14332 => "001001101111010100110111",
14333 => "001011110010111010100100",
14334 => "001101110010111111111000",
14335 => "001111110110110010101110",
14336 => "010001100000001110010010",
14337 => "010000100000000110100010",
14338 => "001010100111011011101110",
14339 => "000001101111010110011111",
14340 => "110111011000010101101111",
14341 => "101011010100110001110110",
14342 => "100010101010101010000101",
14343 => "100001010110111100111111",
14344 => "100010001101000100101001",
14345 => "100001010101010100001100",
14346 => "100001000101101110011101",
14347 => "100001010000001000100001",
14348 => "100000101110011100110110",
14349 => "100011110011000000001111",
14350 => "101100110001001011010000",
14351 => "110111001000111011010110",
14352 => "111111101101011111000011",
14353 => "000110011101001110110101",
14354 => "001001111101011110111100",
14355 => "001001100110100000011000",
14356 => "000111000100000101011010",
14357 => "000011100111110001100010",
14358 => "111111011010111001100010",
14359 => "111010110000100010110000",
14360 => "110111111100001000101010",
14361 => "111000001110100101101000",
14362 => "111000001010111101011100",
14363 => "110101100000001001110110",
14364 => "110010001000000000110100",
14365 => "101110111111001000001000",
14366 => "101100000011001011010010",
14367 => "101001111000110111001110",
14368 => "101000101001100001011110",
14369 => "101000000010011010100100",
14370 => "100111011001101100011001",
14371 => "100111010101100000000001",
14372 => "101000110010011001011010",
14373 => "101010011100110111000000",
14374 => "101011111001011001001100",
14375 => "101110100000011011000110",
14376 => "110010011010011100011110",
14377 => "110110010111101101100100",
14378 => "111000110100010110101011",
14379 => "111010100011101100011111",
14380 => "111101011111010001110110",
14381 => "111111111010001110100001",
14382 => "000000011011001111111001",
14383 => "000000011100010000011000",
14384 => "111111110001111010110001",
14385 => "111101111000100101110010",
14386 => "111011011100100101101101",
14387 => "111001100100000100100100",
14388 => "111001110011111100000000",
14389 => "111011011011001100010001",
14390 => "111100101101111100010110",
14391 => "111110101110010100010001",
14392 => "000001110010011011111110",
14393 => "000100101011100101010001",
14394 => "000111011101010011101000",
14395 => "001010111110000100110110",
14396 => "001111011010111001101000",
14397 => "010011110001110110110110",
14398 => "010111001110101010010000",
14399 => "011001111100101110000111",
14400 => "011011111001000001010001",
14401 => "011101000101001010010110",
14402 => "011101001101100011101101",
14403 => "011100000110010000101001",
14404 => "011011000100110110010000",
14405 => "011010100011001000001001",
14406 => "011001110011111111100101",
14407 => "011000111111000100001001",
14408 => "011000000010011101110111",
14409 => "010111110101100110111110",
14410 => "011000000111010100110000",
14411 => "010101000100011110011100",
14412 => "001111000110101101011110",
14413 => "001010011000111000101001",
14414 => "000110001000101101100001",
14415 => "000001000101110101000011",
14416 => "111100101111000110100100",
14417 => "111001001000001010001000",
14418 => "110110010001111000110010",
14419 => "110011110010001001001110",
14420 => "101111100100010101001000",
14421 => "101001011000110110010100",
14422 => "100100001110010100001011",
14423 => "100010101111000111111110",
14424 => "100011111001011010100101",
14425 => "100110011100000011001111",
14426 => "101010100101100101101000",
14427 => "101101111001100110000110",
14428 => "101110100010010011111110",
14429 => "101110111010110110011110",
14430 => "110000011101010001001000",
14431 => "110010001010001111010010",
14432 => "110100001000100000100000",
14433 => "110110101000100000011101",
14434 => "111000000100011100001010",
14435 => "110110111001100111000110",
14436 => "110011110010111110000010",
14437 => "110000101001001101000110",
14438 => "101110101110000110001000",
14439 => "101110110010010100011110",
14440 => "110001010110110011010000",
14441 => "110110000101110010010010",
14442 => "111011111000001100010111",
14443 => "000001010010101110111111",
14444 => "000101010111100100111011",
14445 => "000111111101001000001001",
14446 => "001001011110001000011010",
14447 => "001011010100010010101010",
14448 => "001110111100111000011110",
14449 => "010100000101110111010000",
14450 => "011000110001010010001011",
14451 => "011011111000001000010001",
14452 => "011101110000000101001101",
14453 => "011101000001110011111011",
14454 => "011001011110101000110111",
14455 => "010110001101111001001110",
14456 => "010100010101100100000100",
14457 => "010100011000010010100110",
14458 => "010111010111101101100110",
14459 => "011010101000101101100000",
14460 => "011011110110100100010001",
14461 => "011011100011010011010011",
14462 => "011001111011001110101101",
14463 => "010111010100101111010010",
14464 => "010100110001110001000000",
14465 => "010011010011001001010100",
14466 => "010011011100101011100000",
14467 => "010011111111111110110110",
14468 => "010010110001110111000110",
14469 => "001110111011111010001100",
14470 => "001000011111101101110000",
14471 => "000000010100011010100100",
14472 => "111000110001001111110101",
14473 => "110011010111001101010000",
14474 => "101111110100010011011110",
14475 => "101100010111010010100100",
14476 => "100111010010111000100111",
14477 => "100010110100010100100001",
14478 => "100001011101010111110111",
14479 => "100001100100100111111110",
14480 => "100001011011010100111011",
14481 => "100001011101100111110101",
14482 => "100011011001000000101101",
14483 => "101000111111010110000010",
14484 => "110001110010100010011010",
14485 => "111011001011010111010110",
14486 => "000001111100010000011010",
14487 => "000101010110111101011000",
14488 => "000111111010101011000100",
14489 => "001001110011000111110000",
14490 => "001001100010000110001010",
14491 => "001000011001101110011001",
14492 => "000101111011001010010000",
14493 => "111111110001010111011110",
14494 => "110111110110111001000010",
14495 => "110000110110101011000000",
14496 => "101010110001111110001100",
14497 => "100110011010110011000010",
14498 => "100101010011011010000111",
14499 => "100111000110010000110101",
14500 => "101010000110111111000000",
14501 => "101110001110111000000100",
14502 => "110011101110011001011000",
14503 => "111000110011010000110001",
14504 => "111100101100001011101100",
14505 => "000000010110101000010101",
14506 => "000100001001110111001011",
14507 => "000110111010011001010100",
14508 => "000110100111010000110100",
14509 => "000100001001010111111000",
14510 => "000001101110101101110001",
14511 => "111110111001100011110010",
14512 => "111100000001101111010100",
14513 => "111011000101001000010111",
14514 => "111011011111010011101001",
14515 => "111011100001110101110111",
14516 => "111011111011001111001001",
14517 => "111101110011111111110010",
14518 => "111111111010100101111001",
14519 => "000001100000110000000001",
14520 => "000011100000000101011100",
14521 => "000101011011111001001001",
14522 => "000110010101101100111010",
14523 => "000110010000101001101110",
14524 => "000101111011011000010101",
14525 => "000110101011010001110000",
14526 => "001000011011100101001111",
14527 => "001001111010000011010100",
14528 => "001011101100010100100110",
14529 => "001110010110001100011100",
14530 => "010000101001100101010010",
14531 => "010010010101010000010000",
14532 => "010011101010011011010100",
14533 => "010011111110010111010100",
14534 => "010011100111111011100010",
14535 => "010100000011010000010010",
14536 => "010100110000101100110010",
14537 => "010011101010011000000110",
14538 => "010000110101010110111110",
14539 => "001110000010110010111010",
14540 => "001011101100010000110110",
14541 => "001001011011011001000100",
14542 => "000111010010000110110010",
14543 => "000101010111101011000110",
14544 => "000011111101101100101001",
14545 => "000011000001010110111001",
14546 => "000001111010010110011001",
14547 => "000000010001110100111000",
14548 => "111110000001000011101010",
14549 => "111011100111101111000001",
14550 => "111010001010100001110100",
14551 => "111000101000011001110001",
14552 => "110101011110110110001001",
14553 => "110001111001100000100110",
14554 => "101111000110110111111110",
14555 => "101101001001110011110000",
14556 => "101100010111001011010010",
14557 => "101101000100001010100010",
14558 => "101101100010110010101010",
14559 => "101010100110011100000010",
14560 => "100110001101000101100011",
14561 => "100101000100000011000101",
14562 => "100110000100110010100011",
14563 => "100110100010110011111011",
14564 => "100110101001100111000111",
14565 => "100111011010110110001010",
14566 => "101001110000001100011010",
14567 => "101100101010010101100000",
14568 => "101110101110111101100010",
14569 => "110001001010011111001110",
14570 => "110101110001000100011000",
14571 => "111100010101001100000001",
14572 => "000010111111001100111001",
14573 => "001000010010001111010100",
14574 => "001100100011001100001000",
14575 => "010000101000011110101100",
14576 => "010100001111011001101010",
14577 => "010110100111010100011110",
14578 => "011000000101101010101111",
14579 => "011010011010010110110110",
14580 => "011101010010100010110111",
14581 => "011101100111011110001101",
14582 => "011100010101110101100111",
14583 => "011100001111001001011011",
14584 => "011011110101100010100111",
14585 => "011010101111001111100011",
14586 => "011001111001111110111101",
14587 => "011001000101011100010010",
14588 => "011000101111111110000110",
14589 => "010111011100000000010100",
14590 => "010011110010001101000100",
14591 => "010000010010110000010000",
14592 => "001110000010101100100010",
14593 => "001011100100101100101010",
14594 => "001001110110011100010001",
14595 => "001010100111100111101011",
14596 => "001101011000001011100000",
14597 => "010000110111100111010100",
14598 => "010011011100000000100110",
14599 => "010100011001101111011100",
14600 => "010011001110101110101110",
14601 => "001110001100010001111000",
14602 => "000110111100110010010011",
14603 => "111111111001011010010010",
14604 => "111001001001101110101111",
14605 => "110010011010010110011110",
14606 => "101001110011000111000010",
14607 => "100010011000011100100011",
14608 => "100000111011111100000101",
14609 => "100001101101000101100001",
14610 => "100001101101100110000101",
14611 => "100001111110001100100001",
14612 => "100001101101011101010011",
14613 => "100001110011000110010111",
14614 => "100011111001001101110011",
14615 => "100110101000100010011111",
14616 => "100111101100010011001110",
14617 => "100111010001000110100100",
14618 => "100111010111000111110010",
14619 => "101000110011010110010010",
14620 => "101011001010000110011110",
14621 => "101110000100101111001000",
14622 => "110001100100111001010010",
14623 => "110100101011010101001100",
14624 => "110110101001011011101000",
14625 => "111000010100000011111000",
14626 => "111001011001010001110011",
14627 => "111001001001111000101010",
14628 => "111000001101101011001111",
14629 => "110111101010011111010110",
14630 => "110110110101101010000111",
14631 => "110100011010011001100110",
14632 => "110010101110110011111100",
14633 => "110100000101000110000001",
14634 => "110111001001001001010110",
14635 => "111011001110110110100100",
14636 => "000001100100001100001100",
14637 => "001010000100110011000100",
14638 => "010010001000100001011010",
14639 => "011000011000100011010011",
14640 => "011100101110010010110001",
14641 => "011110000011101100001001",
14642 => "011100011010110100110001",
14643 => "011000101111000010111111",
14644 => "010100101011000100100010",
14645 => "001111101011110010111010",
14646 => "000111011100111001010111",
14647 => "111110111011001110111111",
14648 => "111000111011111010110111",
14649 => "110100100111000111000011",
14650 => "110010000011111111110100",
14651 => "110001010101110100100000",
14652 => "110010101001010011011100",
14653 => "110101100101000101011110",
14654 => "111001011110110101000010",
14655 => "111111010011011100100100",
14656 => "000110010101010000010001",
14657 => "001100010110100001100110",
14658 => "010000000011001010101110",
14659 => "010001011001111000100010",
14660 => "010001001001000011111100",
14661 => "001111101011010000110010",
14662 => "001101000010110111010010",
14663 => "001001001000101110011011",
14664 => "000101011010111110101100",
14665 => "000011111111001101011010",
14666 => "000101000111001000101011",
14667 => "000110110110000100011111",
14668 => "000110011111100110000101",
14669 => "000100111101000101111001",
14670 => "000100010110000011001010",
14671 => "000100010100001001101101",
14672 => "000100001010110000111001",
14673 => "000011011101100011000001",
14674 => "000010110010110110001101",
14675 => "000010011000010111001000",
14676 => "000001111000100000111101",
14677 => "000001010110001110000000",
14678 => "111111010101110000101101",
14679 => "111100010011111100110000",
14680 => "111010001111010110111100",
14681 => "111010000001101110011110",
14682 => "111100000011101111111011",
14683 => "111101110101010111001001",
14684 => "111101101110110010100110",
14685 => "111101000000100101110101",
14686 => "111100000101100011010010",
14687 => "111011001011001100011101",
14688 => "111001111000001100101101",
14689 => "110111111110011010010010",
14690 => "110110010100110111010001",
14691 => "110100011110100001010010",
14692 => "110000111101110110011100",
14693 => "101100011110101101011000",
14694 => "101001100101000011000000",
14695 => "101000011010110111011100",
14696 => "101000001111000000111000",
14697 => "101000111010111101110010",
14698 => "101001100000011110100000",
14699 => "101010001010111010110110",
14700 => "101010110001001110010100",
14701 => "101011000011110010111100",
14702 => "101011011101100101001100",
14703 => "101011100010001001010000",
14704 => "101101100010101110000010",
14705 => "110010100101100001011010",
14706 => "110111100011111110111001",
14707 => "111011100110001111110110",
14708 => "111111110001111110001000",
14709 => "000101001010101100000000",
14710 => "001011110000111111110010",
14711 => "010001110001011101111110",
14712 => "010111000000010100011110",
14713 => "011011110000101001000010",
14714 => "011110010001100010111001",
14715 => "011110100001000000010001",
14716 => "011110100001010111001000",
14717 => "011110000001111100100100",
14718 => "011100110000001001001001",
14719 => "011011110110011010110101",
14720 => "011011001011000001110101",
14721 => "011010101111101111101001",
14722 => "011010010110110000101101",
14723 => "011001110111100101011011",
14724 => "011001110011101110101111",
14725 => "011001011000101101111011",
14726 => "011001001101001101010100",
14727 => "011001010111010000110101",
14728 => "011000111110010000111111",
14729 => "011000101111101011101011",
14730 => "011000001110100111001011",
14731 => "011000001101110101100111",
14732 => "010110100101000001001000",
14733 => "001110001110100111001100",
14734 => "000100001101100001101001",
14735 => "111111000100001010101100",
14736 => "111011111101101111101100",
14737 => "110111111000000100000100",
14738 => "110100000010000110001000",
14739 => "110010001001001100010100",
14740 => "110000100000110001011000",
14741 => "101100100100010110100010",
14742 => "100111101010011101100100",
14743 => "100100111101000111110011",
14744 => "100101001111011110010101",
14745 => "100101111101001001111010",
14746 => "100101011111101101100101",
14747 => "100101000011101001100110",
14748 => "100101010001000011111011",
14749 => "100110001100101010010011",
14750 => "100111111001000111110001",
14751 => "101001111001001110000010",
14752 => "101100001100111110111000",
14753 => "101110111010011010011000",
14754 => "110000111000101001101010",
14755 => "110001000101001110001000",
14756 => "101111111101111110011110",
14757 => "101101110101100101100010",
14758 => "101011001000110011111010",
14759 => "101001001100001101010110",
14760 => "101000110011110000111100",
14761 => "101010001001011001000110",
14762 => "101101001101001100111010",
14763 => "110010001110110110000100",
14764 => "110111110001101010010100",
14765 => "111011111100010101010101",
14766 => "000000001010110110110011",
14767 => "000101110001110111000010",
14768 => "001100000011011010010000",
14769 => "010001100010001000110010",
14770 => "010100101000001110101000",
14771 => "010110001111110111101000",
14772 => "010111100110000111000010",
14773 => "011000000111111001101000",
14774 => "011000000101111001000100",
14775 => "010111110111101110101100",
14776 => "010110100100001011101000",
14777 => "010011100011011110110000",
14778 => "001111110011001000010010",
14779 => "001100010010000111001100",
14780 => "001001000111011100101110",
14781 => "000110010011000110100100",
14782 => "000011011000001000100001",
14783 => "000000010110100100100100",
14784 => "111101100101011110011000",
14785 => "111011000001001010011011",
14786 => "111001001000010011100101",
14787 => "111000100110000001110010",
14788 => "111001101010001110100101",
14789 => "111011111011000101000110",
14790 => "111111001001100011010101",
14791 => "000011001100010100100001",
14792 => "000110101100111111001000",
14793 => "001000101011001011110010",
14794 => "001000110100001000100101",
14795 => "000111110100111100010110",
14796 => "000111010001100111110101",
14797 => "000110000111101011011001",
14798 => "000010011111001001011101",
14799 => "111100111100000011111101",
14800 => "110111001110000101100111",
14801 => "110010011101011101101100",
14802 => "101110011111101100001000",
14803 => "101100010000011001011000",
14804 => "101100111000001000111110",
14805 => "101111010001100110001010",
14806 => "110011010011111110000010",
14807 => "111000110010011001101000",
14808 => "111110001000010000000001",
14809 => "000011000110001100010010",
14810 => "000110110100101001111100",
14811 => "001001000101110001110100",
14812 => "001011101110111001001010",
14813 => "001101110111011100100010",
14814 => "001101111011010011111100",
14815 => "001100010111010100111010",
14816 => "001001110100001110101000",
14817 => "000111110000011001000000",
14818 => "000110101000000100010000",
14819 => "000101101010111001111001",
14820 => "000101011101110100001011",
14821 => "000110110000111010001110",
14822 => "001001000101100001111001",
14823 => "001001101110011000010000",
14824 => "000111100001001000010100",
14825 => "000101111001001100001111",
14826 => "000101111110100110011010",
14827 => "000100111010000010111010",
14828 => "000001111111100001100010",
14829 => "111111010100101100100110",
14830 => "111101110110011101001110",
14831 => "111100000010010001001100",
14832 => "111000110001000111011110",
14833 => "110101100001011110011000",
14834 => "110100010101110000010010",
14835 => "110100100010010000100110",
14836 => "110011110101111111111010",
14837 => "110001010100001101000000",
14838 => "101100111001010110111000",
14839 => "101000110110001000000100",
14840 => "100111111000100110100101",
14841 => "101000010011001010000010",
14842 => "101000001010011011100000",
14843 => "101000111111111100000000",
14844 => "101100001000011110110110",
14845 => "110000011100010100101000",
14846 => "110100100011011100001001",
14847 => "111000111100111010011010",
14848 => "111101010000001010101011",
14849 => "000000111010011010001011",
14850 => "000101100010100001011011",
14851 => "001010100001100000110001",
14852 => "001110110110001111100000",
14853 => "010100000010101010000110",
14854 => "011000101110111111000000",
14855 => "011011001101000110011011",
14856 => "011100100101000000100110",
14857 => "011100010100000110111110",
14858 => "011011001101011000010000",
14859 => "011010110011011001001101",
14860 => "011001110100001110110011",
14861 => "011001010001100110011110",
14862 => "011000111111101100011001",
14863 => "010110001100010110110110",
14864 => "010001011011101001111100",
14865 => "001011100010000000111010",
14866 => "000101101011011110001000",
14867 => "000000110000101010110101",
14868 => "111100011100100001111110",
14869 => "111010100101011010111010",
14870 => "111010000110111011110110",
14871 => "111001010010111001011000",
14872 => "111001001110111001110000",
14873 => "111001111100111111100010",
14874 => "111101010111100000100000",
14875 => "000011110001101010011000",
14876 => "001010000011111110110010",
14877 => "001110100110011010111110",
14878 => "010000110010100110110010",
14879 => "010001011100000010011000",
14880 => "010000001001110010111100",
14881 => "001100110010111101100010",
14882 => "001001110101100001011011",
14883 => "000111010111011010110001",
14884 => "000100110000011110001011",
14885 => "000001001001110000010011",
14886 => "111011101110010110001111",
14887 => "110101111000101111100100",
14888 => "101111101001000101000000",
14889 => "101010000100010010100110",
14890 => "100111010100001001011011",
14891 => "100101111000100100000001",
14892 => "100100011011010001010010",
14893 => "100011100100110001111011",
14894 => "100011011101001111111111",
14895 => "100011100100100000111111",
14896 => "100011111111011001111001",
14897 => "100101000101000011010111",
14898 => "100101101110101101110110",
14899 => "100101111100010010000101",
14900 => "101001101000000011010110",
14901 => "110010010011011110101000",
14902 => "111011000101110010100100",
14903 => "000000101100001110111101",
14904 => "000100011101010110011011",
14905 => "001000001111011110010000",
14906 => "001100001111110010100110",
14907 => "001110101011010100011000",
14908 => "010000011011100111110000",
14909 => "010010011100111010010110",
14910 => "010010001010011110011110",
14911 => "010000011010100101010000",
14912 => "001110100110111000010010",
14913 => "001011101011101000011000",
14914 => "000111101110100111010011",
14915 => "000100011110011011111010",
14916 => "000101000010110110000000",
14917 => "000111110001011101010000",
14918 => "001000101000011111000010",
14919 => "001000000011100111101001",
14920 => "000111000001010011111111",
14921 => "000110010110000001010011",
14922 => "000110001001101011110010",
14923 => "000110010101010101011101",
14924 => "000111000101110011011111",
14925 => "000110110011111001100101",
14926 => "000110000010101010011110",
14927 => "000110001101100111100001",
14928 => "000110100111100100000000",
14929 => "000101100011010101011100",
14930 => "000010100001101010111011",
14931 => "000000010100010001010010",
14932 => "111110111011001101111010",
14933 => "111100111011001010110000",
14934 => "111011001001011001000101",
14935 => "111000011111110000001110",
14936 => "110100110001111011100110",
14937 => "110001000011101001001100",
14938 => "101110000100100011010110",
14939 => "101011110101111011111010",
14940 => "101001001100101001001000",
14941 => "101000001010010001011010",
14942 => "101001111100110110110010",
14943 => "101101010000001101111110",
14944 => "110010011001000010010100",
14945 => "111000010101100000110111",
14946 => "111101011011001101011101",
14947 => "000001101100011110100000",
14948 => "000110010010000101111111",
14949 => "001010101100011011000000",
14950 => "001011111110011010001000",
14951 => "001010100001010011101111",
14952 => "001000111000100110111100",
14953 => "000110111111000100110000",
14954 => "000011101011011011110101",
14955 => "111111000011011100011000",
14956 => "111010110100110010101101",
14957 => "111000100101010001100000",
14958 => "111000000101100011110110",
14959 => "111000011011101011011110",
14960 => "111011010011100110110100",
14961 => "000001111001011010101110",
14962 => "001001011001010011011000",
14963 => "001111101011110110110100",
14964 => "010100000110100011100110",
14965 => "010110111111111111101010",
14966 => "011000100001100111101001",
14967 => "010111000100011011010000",
14968 => "010011101111101101111100",
14969 => "001111111111110001100010",
14970 => "001011111100110011000100",
14971 => "001000010111001001011000",
14972 => "000101001111011110001011",
14973 => "000100000010010101000100",
14974 => "000100111001010001010110",
14975 => "000110001000100101010100",
14976 => "000111010010001100111110",
14977 => "000110111110011000110101",
14978 => "000101000110100100001101",
14979 => "000010110101101001111110",
14980 => "000000111110000111011111",
14981 => "000000000001011101000000",
14982 => "000000100100110110001101",
14983 => "000011101101011010100000",
14984 => "000110101101111010101011",
14985 => "000111010110101111000100",
14986 => "000111000011100010001110",
14987 => "000110010000011111101011",
14988 => "000110011110110100101111",
14989 => "000111110011110010000111",
14990 => "001000101111110110001001",
14991 => "001001000011000011001111",
14992 => "000111001000010101010100",
14993 => "000011001101001011100101",
14994 => "111110011010010100000001",
14995 => "111001001001100001001001",
14996 => "110011110111111101110000",
14997 => "101110010001001110111110",
14998 => "101010100110011000110100",
14999 => "101001011100110010111100",
15000 => "101000001001001011100010",
15001 => "100110100100010010001101",
15002 => "100101100011110110110111",
15003 => "100110100010100001110001",
15004 => "101010001110000000111010",
15005 => "101110110111011010010000",
15006 => "110011100010100111111010",
15007 => "111000001110111010101100",
15008 => "111100100011111100010011",
15009 => "111111011101100011001101",
15010 => "000000000100001111101010",
15011 => "111110010111011111101001",
15012 => "111011010101011110001000",
15013 => "111001110011010101110001",
15014 => "111010110101101110011111",
15015 => "111011100101111101101111",
15016 => "111010111110111110100010",
15017 => "111010111100111011001110",
15018 => "111010000101111011000011",
15019 => "110110001000011000011110",
15020 => "110010000011000011100000",
15021 => "110000110010010010100000",
15022 => "110000111000100100001100",
15023 => "110000010111110000101000",
15024 => "110001011100111110000110",
15025 => "110101110010000101101110",
15026 => "111001011010101110011110",
15027 => "111100010001110111000101",
15028 => "000000111110011110010100",
15029 => "000101110100111000101000",
15030 => "001010001111101101101100",
15031 => "001101111010001001111000",
15032 => "010001010000101011010100",
15033 => "010011110111011111110000",
15034 => "010010000011100111011010",
15035 => "001110110001001000101010",
15036 => "001101110011010101001100",
15037 => "001100101010110110111110",
15038 => "001010011111111110110110",
15039 => "001000110011110110000000",
15040 => "001000110101100011111111",
15041 => "001001100101000100010100",
15042 => "001011001000010000011000",
15043 => "001110101000000011110010",
15044 => "010000011110110011011000",
15045 => "010000100110111001011000",
15046 => "010010100101000100100010",
15047 => "010100111000010010100110",
15048 => "010100110010111010111000",
15049 => "010001001000000111110100",
15050 => "001011110110000011111110",
15051 => "000111110010011101100100",
15052 => "000011101001110010001111",
15053 => "000000001111111010110011",
15054 => "000000000111011101110101",
15055 => "000000101110011101000010",
15056 => "111111101101011101110101",
15057 => "111111000110111001001001",
15058 => "000000001100011011101000",
15059 => "000000000111010101011111",
15060 => "111100101011100111100011",
15061 => "111001100001010111101010",
15062 => "111001101001111111111000",
15063 => "111001100111010100000111",
15064 => "110110101101011101101010",
15065 => "110010011110111010110010",
15066 => "101110010010001101111100",
15067 => "101010000011011101010110",
15068 => "100101011011110011100010",
15069 => "100010010011000101101101",
15070 => "100010011010101010110101",
15071 => "100011101000110101111001",
15072 => "100100010010011101001001",
15073 => "100100110000110011110010",
15074 => "100101001111011110010001",
15075 => "100101111010101100011101",
15076 => "100110011110111101010010",
15077 => "100111001111000110000011",
15078 => "101001011000001110101110",
15079 => "101100111100111010100100",
15080 => "110000101010101000000110",
15081 => "110011010000100100111000",
15082 => "110101011101101101010001",
15083 => "111001000001101110101000",
15084 => "111101010110011110010101",
15085 => "000000010110000011001101",
15086 => "000010000110000001010000",
15087 => "000100100011101000100000",
15088 => "000111001110110101110000",
15089 => "000111111101111000000111",
15090 => "000111011011001110111011",
15091 => "000111010011101010000010",
15092 => "001000000010001111111110",
15093 => "001001100100001010010000",
15094 => "001011100110111100011010",
15095 => "001110011101111000000110",
15096 => "010001101001010100001110",
15097 => "010100101101001100010000",
15098 => "011001000010011010100101",
15099 => "011101000110110011110101",
15100 => "011110100000110101001110",
15101 => "011110011100101100110011",
15102 => "011101111001010111101000",
15103 => "011101010100111010101101",
15104 => "011100111110000110000011",
15105 => "011100011000100111100000",
15106 => "011011101111011100011111",
15107 => "011011000001101101011100",
15108 => "011010011001010010101011",
15109 => "011000011100001000010001",
15110 => "010011111111000110100000",
15111 => "001111100010010001011010",
15112 => "001100101010110011111110",
15113 => "001011100101111001101011",
15114 => "001100001111110000110000",
15115 => "001101010101101110000000",
15116 => "001110100101010110111110",
15117 => "001110111100101001111100",
15118 => "001011101000101001011100",
15119 => "000100010111110010000100",
15120 => "111100101101010011000010",
15121 => "110110011111100001111001",
15122 => "110000101010000011100100",
15123 => "101011010010011100011110",
15124 => "100101110100100010011111",
15125 => "100001101001011001100001",
15126 => "100001011000000000001011",
15127 => "100001111110100001011001",
15128 => "100001110011000101010111",
15129 => "100010000100010010011011",
15130 => "100010000010001011110011",
15131 => "100010111110011111101101",
15132 => "100110111110111001000000",
15133 => "101101011101111010111100",
15134 => "110011111111011011001110",
15135 => "111001100100001110000100",
15136 => "111110001100010000101011",
15137 => "000000100110001100001101",
15138 => "000010100001001111010100",
15139 => "000101011010100110111000",
15140 => "000110101100100000000011",
15141 => "000101000001011111110001",
15142 => "000001000110000111001100",
15143 => "111101000100110101100001",
15144 => "111010101101000100001111",
15145 => "111001010100110111000011",
15146 => "110111101001000100001111",
15147 => "110100101111001010011111",
15148 => "110001011110000100110100",
15149 => "101110011101110011000110",
15150 => "101011010110011001011100",
15151 => "101001010001100011101000",
15152 => "101000101111001111111110",
15153 => "101000110100001111000010",
15154 => "101001101111010100010100",
15155 => "101100101111001001000100",
15156 => "110001110000011101110010",
15157 => "110111111111110011100111",
15158 => "111110110000101001111101",
15159 => "000100001111111101001000",
15160 => "000111011100100000100011",
15161 => "001001110011001100111001",
15162 => "001101000111111110110100",
15163 => "010000000010000010001010",
15164 => "001111110111111001101100",
15165 => "001101101111111101110010",
15166 => "001011011111101000010110",
15167 => "001001010011101011001100",
15168 => "000110001000100001111101",
15169 => "000001100101011101100000",
15170 => "111110011011001101010010",
15171 => "111100100100100101111010",
15172 => "111010110011101101000111",
15173 => "111010111000000101110000",
15174 => "111100100010100100111101",
15175 => "111110110111011100110001",
15176 => "000001000110000010101100",
15177 => "000011110101001010110110",
15178 => "001000011010101010111111",
15179 => "001100110001010101110000",
15180 => "010000110110111001010110",
15181 => "010101110010110011001100",
15182 => "011010010000110011111111",
15183 => "011101001001100000000110",
15184 => "011101001011010110100111",
15185 => "011011110110100000101011",
15186 => "011011000010111101110011",
15187 => "011010000001111110110101",
15188 => "011001001101100110110110",
15189 => "011000011001010011111101",
15190 => "010111100101110010010000",
15191 => "010111000111001101111000",
15192 => "010100111100111011010100",
15193 => "010001001100100111101110",
15194 => "001101100110011100110000",
15195 => "001001110011010111110001",
15196 => "000110011011101110010101",
15197 => "000100110101011010011110",
15198 => "000011111011110100101000",
15199 => "000010010111110001001100",
15200 => "111111001100011000010010",
15201 => "111010101100011001010000",
15202 => "110110011111111100010100",
15203 => "110001101010001110101100",
15204 => "101011110110101101010100",
15205 => "100110110000111100111111",
15206 => "100011010111110011100001",
15207 => "100010111011000101100011",
15208 => "100011110101011000010111",
15209 => "100100010110100001100101",
15210 => "100101011001000111100101",
15211 => "100110001101100100100001",
15212 => "100110010001001011111111",
15213 => "100110010011101100011111",
15214 => "100111010110000001101111",
15215 => "101001100001011111111010",
15216 => "101011110010011110011110",
15217 => "101110000110100000101100",
15218 => "110000001000111001111110",
15219 => "110010001100110101000110",
15220 => "110011111110011110111010",
15221 => "110011110011101101000110",
15222 => "110010110001010110011000",
15223 => "110010011101010000111010",
15224 => "110011101100110101111100",
15225 => "110110011100110101111001",
15226 => "111010100110110001110001",
15227 => "000000001000010111110010",
15228 => "000100010011100100111000",
15229 => "000110110010010001101000",
15230 => "001001001010010111111010",
15231 => "001100010110110100001010",
15232 => "010000011110101101000110",
15233 => "010011101001011111110110",
15234 => "011000000010101011000111",
15235 => "011100111111100000101101",
15236 => "011110001101001100110111",
15237 => "011110010101001101011011",
15238 => "011110010011100110010001",
15239 => "011101010110011110110010",
15240 => "011100011101000001010101",
15241 => "011010111110100111001001",
15242 => "011010001010110111111011",
15243 => "011010000000101100101111",
15244 => "011001101011111100011011",
15245 => "011001010111001010111001",
15246 => "011000101100011110011001",
15247 => "011000000110010110111111",
15248 => "010111011111111000101010",
15249 => "010111010011000000000110",
15250 => "010110000101101110100110",
15251 => "010011110001100100110110",
15252 => "010010011101001101101010",
15253 => "010000001101011000000010",
15254 => "001100010010101000111000",
15255 => "000101101010010000100110",
15256 => "111110010001111101010100",
15257 => "111000111111010010001101",
15258 => "101110010101111000111000",
15259 => "100010101111000101001010",
15260 => "100000111111011100110011",
15261 => "100001111100011100011001",
15262 => "100001010011001101100111",
15263 => "100001111011001100010000",
15264 => "100001111011000010011010",
15265 => "100001100100011001101111",
15266 => "100010011000100000101011",
15267 => "100010110000111010101100",
15268 => "100100001001110010101101",
15269 => "101011010110110101100100",
15270 => "110100101001010111101100",
15271 => "111010101101110010001000",
15272 => "000000001010010010000101",
15273 => "000011111011101110110110",
15274 => "000011110011011011110010",
15275 => "000001011101101101100010",
15276 => "111110110001100101010001",
15277 => "111100011110001000000010",
15278 => "111000010101011100010111",
15279 => "110100001000011001101010",
15280 => "110010010101110100110100",
15281 => "110000001011010111110000",
15282 => "101110001111101111011110",
15283 => "101110100011010110010010",
15284 => "110000110010000001110110",
15285 => "110100011011000110011100",
15286 => "111000110110001101000101",
15287 => "111110000011100100100100",
15288 => "000011001011001011010100",
15289 => "000111100101000010111001",
15290 => "001011011000110001010000",
15291 => "001110001000111110111010",
15292 => "001110110111011110010110",
15293 => "001101000001001101111010",
15294 => "001010111110011111111010",
15295 => "001001110011110100001110",
15296 => "001000000000000000111111",
15297 => "000110100101111001100011",
15298 => "000110101110110101011101",
15299 => "000110010010010000100101",
15300 => "000010101111000011110000",
15301 => "111101011101010011101101",
15302 => "111001000000100000010011",
15303 => "110101110011101110010001",
15304 => "110100011010111000000101",
15305 => "110100010001001100100110",
15306 => "110100011111001011001101",
15307 => "110101011011001010101011",
15308 => "110110110011110000010100",
15309 => "111000110110110111100100",
15310 => "111010111101111101101100",
15311 => "111011110100011010011011",
15312 => "111100000010101111001001",
15313 => "111101000101001011000000",
15314 => "111111100101001000001110",
15315 => "000010001011101001011111",
15316 => "000010111011001000101100",
15317 => "000010000100110110011001",
15318 => "000001101001100011000000",
15319 => "000010011101111110110100",
15320 => "000011001010001100001001",
15321 => "000010110110100001001110",
15322 => "000010011011100000111110",
15323 => "000011011011100111011111",
15324 => "000101100000100001110011",
15325 => "000110011111010000010101",
15326 => "000110010010001100011100",
15327 => "000110000001100000101011",
15328 => "000110010101100101000000",
15329 => "000111011010101010100011",
15330 => "001000100101011011110111",
15331 => "001001101101101011100110",
15332 => "001010010110000001000111",
15333 => "001010010001000010001010",
15334 => "001010011111011110001011",
15335 => "001010001000101010111110",
15336 => "001000100100110010100100",
15337 => "000111101010001111110001",
15338 => "000111101101101110011100",
15339 => "000111001110101101010110",
15340 => "000101100100100000010011",
15341 => "000010111000000010101001",
15342 => "111111100101001001010001",
15343 => "111100001111111000110110",
15344 => "111001011011000001100000",
15345 => "110111011001010100101111",
15346 => "110101110011110010011100",
15347 => "110101010101100010011010",
15348 => "110110001001000110001111",
15349 => "110110001101010001000110",
15350 => "110101101001110100010010",
15351 => "110101101111100101001000",
15352 => "110110010010101110111110",
15353 => "110111000010011000110110",
15354 => "111000011101001011111110",
15355 => "111011111111001010111011",
15356 => "111111001000111100001111",
15357 => "111110100110110111011011",
15358 => "111100010111001001001110",
15359 => "111000101001110101011111",
15360 => "110010111111111000111010",
15361 => "101110000010111011011110",
15362 => "101011100010010100101100",
15363 => "101100010110100001000100",
15364 => "110000010000000100001100",
15365 => "110110001011110011001111",
15366 => "111100101010101101110101",
15367 => "000010011011011110110111",
15368 => "001000100111100010101111",
15369 => "001111101111000111100110",
15370 => "010110101110010010000010",
15371 => "011100000001011100010100",
15372 => "011110001100010110101111",
15373 => "011110000111000111100101",
15374 => "011101010001000111000111",
15375 => "011100010000010001010011",
15376 => "011011010100011101100011",
15377 => "011010101000111110101101",
15378 => "011010000001111101001101",
15379 => "011001010010111111100011",
15380 => "011000110100110101001101",
15381 => "011000100011110111110001",
15382 => "011000100110100110011011",
15383 => "011000000111111101001110",
15384 => "010111100100101110101010",
15385 => "010111010111010011111010",
15386 => "010001101111001111010010",
15387 => "000111100111010010010101",
15388 => "000000001000100001111000",
15389 => "111001100000110101100100",
15390 => "110011010001001101110110",
15391 => "110000011010100110100110",
15392 => "110000001111101110110110",
15393 => "110001001110000001010100",
15394 => "110000100111011100010000",
15395 => "101111100011111000001000",
15396 => "110010010110101111110110",
15397 => "110111110101111010000100",
15398 => "111010001110011010000011",
15399 => "110110001110011110001110",
15400 => "101110111010111010100000",
15401 => "100111011110000010101110",
15402 => "100010010110001001101010",
15403 => "100001101101101101010011",
15404 => "100010011000011001011011",
15405 => "100010100000011100110010",
15406 => "100011000110111010001011",
15407 => "100100010100101011010000",
15408 => "100110110110100100110111",
15409 => "101001011111011110011000",
15410 => "101011111000011111010010",
15411 => "101110100001110001000010",
15412 => "101111110111010101100000",
15413 => "110000101101011001100000",
15414 => "110010011000101011111010",
15415 => "110100000001010001110000",
15416 => "110101001000100010011101",
15417 => "110101111110100011001001",
15418 => "110111011001011001011001",
15419 => "111010101100001001110000",
15420 => "000000100111110111101001",
15421 => "000111111100100100110111",
15422 => "001110010111001101001110",
15423 => "010011011000000111010110",
15424 => "010111111101010110100100",
15425 => "011011111111000001001110",
15426 => "011101111011001011000101",
15427 => "011110000101001001001111",
15428 => "011101111111101100100011",
15429 => "011100100000001101110011",
15430 => "011000010011111100011110",
15431 => "010011001100011101011100",
15432 => "001110010111000011000110",
15433 => "001000100001011101010110",
15434 => "000010001010110000111100",
15435 => "111110101101110001000110",
15436 => "111111100000011001000101",
15437 => "000010111001000000001100",
15438 => "001000001111111100010011",
15439 => "001110111011001011010000",
15440 => "010100001110110010111110",
15441 => "010111000001010111011110",
15442 => "011000100011110100100011",
15443 => "011001110101000111011111",
15444 => "011001110111111101011101",
15445 => "010110110101011110010100",
15446 => "010001100001010110011010",
15447 => "001011111001001001101011",
15448 => "000110011111010010011100",
15449 => "000000101001011111111110",
15450 => "111001011011100101101110",
15451 => "110010100111111011111100",
15452 => "101101001100110000101100",
15453 => "101000011001010101111100",
15454 => "100101010111110011010111",
15455 => "100011001110011000101001",
15456 => "100001101001011111011100",
15457 => "100001110110101100010011",
15458 => "100010000010101001010111",
15459 => "100010000100011011111001",
15460 => "100010100111101010110111",
15461 => "100011010000111010010101",
15462 => "100100110010100100100101",
15463 => "100111011000101111110000",
15464 => "101011000100110000110110",
15465 => "101110111011110101100010",
15466 => "110001010100100000001000",
15467 => "110010001101110011100100",
15468 => "110011000000010010001100",
15469 => "110101010100110101110010",
15470 => "111000000011000010100110",
15471 => "111001011011001010110010",
15472 => "111001111001011000000001",
15473 => "111010001001000101111011",
15474 => "111010100111111101100000",
15475 => "111010100110110111000010",
15476 => "111001100001001000001000",
15477 => "111000001001011011000000",
15478 => "110111100101100001110010",
15479 => "111000011000000110011000",
15480 => "111000111001111000011101",
15481 => "111000110000011100010000",
15482 => "111001101100000101101001",
15483 => "111100000110001100001111",
15484 => "111111010101000100110111",
15485 => "000010101000001111011101",
15486 => "000110010011100111100000",
15487 => "001010011110010000101011",
15488 => "001110010010111011100000",
15489 => "010001111100010011110000",
15490 => "010101000000011110011010",
15491 => "010110011111010110010010",
15492 => "010110100100110101101000",
15493 => "010110010000111110001100",
15494 => "010101110111010011111100",
15495 => "010101011100111011010010",
15496 => "010101110100110101001110",
15497 => "010110100101000110100010",
15498 => "010111011101111000111100",
15499 => "011000101001010011110110",
15500 => "011001101001100100100110",
15501 => "011011000000100100100011",
15502 => "011011111001011010101001",
15503 => "011011011111110000101101",
15504 => "011010111000101111000111",
15505 => "011010001101011111110001",
15506 => "011001011101101000111011",
15507 => "011000110001101001100100",
15508 => "011000000110100000010011",
15509 => "010111001110100100011010",
15510 => "010110010001101110100100",
15511 => "010101111011000110110100",
15512 => "010101110110101000001000",
15513 => "010101011011100101110110",
15514 => "010010010011100010000100",
15515 => "001011000001110100110000",
15516 => "000001101101111110001000",
15517 => "110111100111101000101011",
15518 => "101110101111001101000000",
15519 => "101001000100101101101100",
15520 => "100101110110110101100001",
15521 => "100100001101110111011011",
15522 => "100100000011000100111001",
15523 => "100110001110110100111001",
15524 => "101001111001100110101010",
15525 => "101110001000000001011000",
15526 => "110011010101010001101100",
15527 => "111000001011001001101111",
15528 => "111100010101111110010101",
15529 => "111111001110000011100110",
15530 => "000001000101001100101100",
15531 => "000010100111110000011011",
15532 => "000000101101100100100101",
15533 => "111100011000011001001100",
15534 => "111000001111000001111001",
15535 => "110011011010110011010010",
15536 => "101110101010011010010010",
15537 => "101011101110111101011000",
15538 => "101010011110101101100110",
15539 => "100110101100011110001111",
15540 => "100010100011000111011001",
15541 => "100011101100100101001001",
15542 => "100101001100010101100000",
15543 => "100101100010111010001101",
15544 => "100110111101110011011111",
15545 => "100111011001101001010111",
15546 => "100111110111111010111111",
15547 => "101000011110100000110110",
15548 => "101010111011010010100110",
15549 => "110001010111111101100100",
15550 => "111001001000110111101000",
15551 => "000001111001100011110010",
15552 => "001011000101100111101001",
15553 => "010011001011001000110000",
15554 => "011001000011110000110111",
15555 => "011011110000001101010001",
15556 => "011100101101100010111110",
15557 => "011010010100101011100101",
15558 => "010100011011100001011010",
15559 => "010000001110001011010000",
15560 => "001111110011101101100100",
15561 => "010000111110011000001110",
15562 => "010000100000100000100010",
15563 => "001110100101010010011110",
15564 => "001100110001011011011000",
15565 => "001010101010101011110100",
15566 => "001001101001111001110011",
15567 => "001010101111011111001100",
15568 => "001100000000000101011100",
15569 => "001011111011011100001101",
15570 => "001100001100001010011010",
15571 => "001110000001000011010110",
15572 => "001110001110010000110000",
15573 => "001011010010111100000000",
15574 => "000111110110010010001010",
15575 => "000110010101010110001001",
15576 => "000111001101100101111111",
15577 => "001001010011100110001001",
15578 => "001100001111011001001010",
15579 => "001111101100100001111110",
15580 => "010010000111111100110110",
15581 => "010010001100011010110100",
15582 => "001111100111000101001100",
15583 => "001011000000000100111100",
15584 => "000100111011001111100000",
15585 => "111110000010100110100111",
15586 => "110111001100000101101010",
15587 => "110001010010110000011110",
15588 => "101011100111110101101010",
15589 => "100101010110000000111001",
15590 => "100001111100111100111010",
15591 => "100001111001110000001101",
15592 => "100001110111101000110100",
15593 => "100011100110110101001001",
15594 => "101000010111110011111100",
15595 => "101101100011000011010000",
15596 => "110001110010111101101000",
15597 => "110101100010101100000100",
15598 => "111000100000111000110010",
15599 => "111001110010100110110110",
15600 => "111010010100011011101000",
15601 => "111010001111010011011011",
15602 => "111001010010001101010111",
15603 => "111000101001000101100010",
15604 => "110111100111010100001000",
15605 => "110101100001010001000101",
15606 => "110010000011011101001110",
15607 => "101110001101100100111000",
15608 => "101100101010101100101010",
15609 => "101100001000101010110000",
15610 => "101011010000111010110100",
15611 => "101010111000001001100110",
15612 => "101010111011110011011110",
15613 => "101011110100111001010100",
15614 => "101101001010010111001010",
15615 => "101111100111001100100110",
15616 => "110011110001001110001010",
15617 => "110111011010111000110100",
15618 => "111010111011001011011100",
15619 => "111111110111110001001000",
15620 => "000100100000100100101111",
15621 => "000110010011010000110000",
15622 => "000101110110110010011010",
15623 => "000110001100100111010111",
15624 => "000111001000000111001110",
15625 => "000110010011111010011110",
15626 => "000101000100011010001111",
15627 => "000101110111011100001001",
15628 => "000111101001011000101100",
15629 => "001000101100010100101010",
15630 => "001001110001001001010110",
15631 => "001011011101010010101101",
15632 => "001100111010111001101010",
15633 => "001101100000010111100100",
15634 => "001110010001010110111000",
15635 => "010000100001010101100000",
15636 => "010011001001111011100110",
15637 => "010110010010110000001010",
15638 => "011010011111111011001111",
15639 => "011100101101010101011100",
15640 => "011100001000111000011111",
15641 => "011011001010000010100001",
15642 => "011010010010110001010101",
15643 => "011001101001100111000101",
15644 => "011001001000100101110011",
15645 => "011000010110111001010011",
15646 => "010111101011011111111110",
15647 => "010111001110010011100010",
15648 => "010110100110110101110110",
15649 => "010100000000101110100010",
15650 => "001110111010110010100110",
15651 => "001001111001000001000100",
15652 => "000101011000100010001101",
15653 => "000001011100100101110111",
15654 => "111111001010000000011000",
15655 => "111101111010100011100110",
15656 => "111111011100111010010100",
15657 => "000011101101011101111011",
15658 => "000110111010110010110011",
15659 => "001001101010000111100100",
15660 => "001101010011011110011000",
15661 => "010001001001101100011010",
15662 => "010100000011100000101000",
15663 => "010100100100101101001010",
15664 => "010011011111001110010100",
15665 => "010000101011010011100000",
15666 => "001011000111010100101101",
15667 => "000010100010101001011100",
15668 => "111000111110001101110011",
15669 => "110010000000111000011100",
15670 => "101010000110001001111100",
15671 => "100010000001001011000011",
15672 => "100000111101110010010110",
15673 => "100001101111111101010011",
15674 => "100000110101000100101001",
15675 => "100001011100101011110011",
15676 => "100001100010010000001111",
15677 => "100001101000100001000001",
15678 => "100010011110101100110111",
15679 => "100011001000001111101001",
15680 => "100100000111000011101001",
15681 => "100100010100101000111001",
15682 => "100100110000101001110001",
15683 => "100101001000010101011011",
15684 => "100101111000000001101011",
15685 => "101011000100111100100100",
15686 => "110001110100111110011010",
15687 => "110101101111000001011100",
15688 => "110111100101010000011111",
15689 => "111000000110000001011100",
15690 => "111000100110111000010111",
15691 => "111010100101101000111000",
15692 => "111101000011101011100011",
15693 => "111110001001110010000011",
15694 => "111110100010011011111001",
15695 => "111111000000001111011000",
15696 => "111110110100010000011011",
15697 => "111111110010101011011001",
15698 => "000010010000011010101010",
15699 => "000100011100101101111100",
15700 => "000111111010010010010111",
15701 => "001110110101001000010000",
15702 => "011000001000001111100100",
15703 => "011110001100000010110010",
15704 => "011110010010011101001001",
15705 => "011100110101111001101001",
15706 => "011011111101111011100011",
15707 => "011010111011101001100010",
15708 => "011010000100100001101101",
15709 => "011001100110011000000111",
15710 => "011001010010110011101011",
15711 => "011000011000010011010011",
15712 => "010111011101000111010000",
15713 => "010100101011001110010000",
15714 => "001100001110001110111000",
15715 => "000001100110100110000101",
15716 => "111010011111000100111111",
15717 => "110111011100011000000110",
15718 => "110111000000011100101101",
15719 => "110111110111011110110001",
15720 => "111010001000101000000000",
15721 => "111100111011001100100001",
15722 => "111101110110111111001101",
15723 => "111100110010001101100010",
15724 => "111010100111001100001010",
15725 => "111000000111110011010010",
15726 => "110101110100111001001111",
15727 => "110011001111000010011010",
15728 => "101111111101110011110000",
15729 => "101100000000100001100100",
15730 => "101000000010001011001100",
15731 => "100100111110101110011001",
15732 => "100010110010101101011110",
15733 => "100001111111010101100111",
15734 => "100011001011111101110111",
15735 => "100101000000110000001111",
15736 => "100110101000100100010001",
15737 => "101000000101111110100110",
15738 => "101000010011111100010000",
15739 => "100111010011001101001010",
15740 => "100110001001000010100010",
15741 => "100101111011001001100110",
15742 => "100111000111100111001111",
15743 => "100111100110111100010010",
15744 => "100111111001110000001101",
15745 => "101011110000101110111010",
15746 => "110010010110101100001000",
15747 => "111000110010111100110000",
15748 => "111110101100100001000011",
15749 => "000100111000111011111110",
15750 => "001011100011011100100010",
15751 => "010001001011101011000110",
15752 => "010101100100111010010000",
15753 => "011001000011011011110111",
15754 => "011010110010111100000101",
15755 => "011011000010001000100101",
15756 => "011001101100101010011011",
15757 => "010111001010010111011100",
15758 => "010100101000111010000000",
15759 => "010010001111110010010100",
15760 => "010000001010110000011010",
15761 => "001110010010100000000100",
15762 => "001100100011001001100010",
15763 => "001010110000010010100010",
15764 => "001000011100000100000110",
15765 => "000110111000101010001000",
15766 => "000110000100100001010010",
15767 => "000101001111011000001000",
15768 => "000101110101010011010001",
15769 => "000111110111101000101101",
15770 => "001010010110110100101010",
15771 => "001100111011001000111010",
15772 => "001110011001101101100100",
15773 => "001110010101000101011000",
15774 => "001101011111101110100000",
15775 => "001100111000110111100000",
15776 => "001100100101001010101110",
15777 => "001010101001000110100001",
15778 => "000110011011011010010100",
15779 => "000001011110011000110101",
15780 => "111011101010001110110110",
15781 => "110101100101000000000110",
15782 => "101111111000101010101010",
15783 => "101000100010000101011010",
15784 => "100010011001001010010011",
15785 => "100001011000000010010011",
15786 => "100010001110101101000010",
15787 => "100010101011110000100011",
15788 => "100011111011100011000111",
15789 => "101000000100110101110000",
15790 => "101111100110111101110100",
15791 => "110111001000111000001100",
15792 => "111110100001010101001100",
15793 => "000110101110000001001010",
15794 => "001101110010111001111000",
15795 => "010011100100010110110010",
15796 => "010111110011100101100100",
15797 => "011010010101100000111011",
15798 => "011010001111010100001100",
15799 => "010111011010011111101000",
15800 => "010110010000101100111100",
15801 => "010101101101001110101100",
15802 => "010010010000001110001110",
15803 => "001110111101110001010010",
15804 => "001101001000100110001010",
15805 => "001011001000111100000100",
15806 => "000111011110000110011100",
15807 => "000010100001111101101101",
15808 => "000000000000101110100010",
15809 => "111111010101000111000000",
15810 => "111110011000011110010110",
15811 => "111111011101011001110010",
15812 => "000010110111010110000100",
15813 => "000110011010000011011001",
15814 => "001001101001010010111100",
15815 => "001101010001110100101100",
15816 => "010000110000010101111110",
15817 => "010010111100010001000100",
15818 => "010100011110010001111010",
15819 => "010100110101000001000000",
15820 => "010001101110110011101010",
15821 => "001010100110000110101001",
15822 => "000001001011011010111011",
15823 => "111000000011010100110101",
15824 => "101110110001100110100100",
15825 => "100110000011111010001111",
15826 => "100010010111110101001011",
15827 => "100010001011111111110111",
15828 => "100010000000010101000011",
15829 => "100010101110110100000001",
15830 => "100011101100110110001111",
15831 => "100100101010000110100100",
15832 => "100101110010010111101001",
15833 => "100111110011101010001111",
15834 => "101110011001000101010100",
15835 => "110111101100010100011000",
15836 => "000000000011110011000110",
15837 => "001000111000000101101101",
15838 => "010001001101011001100010",
15839 => "010110111010000001010000",
15840 => "011010001010101100111001",
15841 => "011011010110111000110100",
15842 => "011010011001010110011011",
15843 => "011000100010010110001010",
15844 => "010111111111100101101000",
15845 => "010101010100100001011110",
15846 => "001101110101111101010110",
15847 => "000110111100111110011110",
15848 => "000010011111000101110011",
15849 => "111110100101100001000001",
15850 => "111011101100111101100110",
15851 => "111001001000111111111110",
15852 => "110111011110000101100000",
15853 => "110111111001010111100110",
15854 => "111000110110110101001001",
15855 => "111000110101110000111110",
15856 => "111000011111100110011100",
15857 => "111010101010001010010110",
15858 => "000000001000001000111001",
15859 => "000101111010100111010111",
15860 => "001010101000001111001011",
15861 => "001110011111100001100010",
15862 => "010000011011100111011110",
15863 => "001111100110001110100000",
15864 => "001100100000101000000000",
15865 => "001001000101100010000000",
15866 => "000110010100101101110001",
15867 => "000001101100101101011110",
15868 => "111010011000000101101000",
15869 => "110011100110000000000100",
15870 => "101110001100100110100110",
15871 => "101000101001011011111000",
15872 => "100011100111000100010000",
15873 => "100001010100001001100111",
15874 => "100001111100111100101101",
15875 => "100011110001001101111101",
15876 => "100111010001000111011101",
15877 => "101100011100001101101010",
15878 => "110000110100000001011100",
15879 => "110100011000001001110001",
15880 => "110111101001001100010100",
15881 => "111010101010101001000001",
15882 => "111110001011101111111001",
15883 => "000000101101000110111111",
15884 => "000001101000110001100001",
15885 => "000001111101100010001001",
15886 => "000001011000000001011111",
15887 => "000000100110001100101100",
15888 => "000000011111001101000111",
15889 => "000001010000000010011000",
15890 => "000100000110001001100011",
15891 => "001000111110111010111001",
15892 => "001101101101001101001010",
15893 => "010001011000001000001000",
15894 => "010101011000011001000100",
15895 => "011001011001101011001011",
15896 => "011011011100100001110001",
15897 => "011011000100010111101111",
15898 => "011000110111011000110001",
15899 => "010110110001010101000000",
15900 => "010110001101001111010010",
15901 => "010101010001010110101000",
15902 => "010011000100100110100000",
15903 => "010001010000000010111100",
15904 => "010000011000110011101000",
15905 => "010000001011010001110000",
15906 => "010000001001110001110010",
15907 => "001111111100001110100000",
15908 => "001111111001010100100110",
15909 => "001111101100101011001110",
15910 => "001110110101010101111110",
15911 => "001100110010011110111010",
15912 => "000111011110110101011110",
15913 => "111111011000100001111000",
15914 => "110111000011111011000010",
15915 => "101101101000001010001100",
15916 => "100100101110000110011110",
15917 => "100001000011110101010011",
15918 => "100001001111110101101101",
15919 => "100001101111010001100110",
15920 => "100001111110111110000100",
15921 => "100001101001010101010001",
15922 => "100001001011111101110111",
15923 => "100001011011110111101101",
15924 => "100001101010000100111101",
15925 => "100010010110000110000110",
15926 => "100101111100110101111111",
15927 => "101010110000011101001010",
15928 => "101101000011001001100100",
15929 => "101111000000110010011000",
15930 => "110001110100101101001000",
15931 => "110010110111110110110110",
15932 => "110011100010110000111010",
15933 => "110100101111010001111011",
15934 => "110100110011000101111000",
15935 => "110100100100100101100111",
15936 => "110101000000010110100001",
15937 => "110101101010110110010011",
15938 => "110110000010101111001010",
15939 => "110110001110111000011100",
15940 => "110111011010100100000111",
15941 => "111001100110110101100011",
15942 => "111011001100111000011111",
15943 => "111100101100000110000011",
15944 => "000001000011011110000100",
15945 => "001000001000100011010000",
15946 => "001110101111111110111000",
15947 => "010011011111010101000010",
15948 => "010110111010011110011100",
15949 => "011010101111000100111101",
15950 => "011110000100100111000011",
15951 => "011110100000000001000010",
15952 => "011101110010101000111111",
15953 => "011101001111001111000011",
15954 => "011100011100100101111110",
15955 => "011100010011000000101100",
15956 => "011010111001011001010111",
15957 => "010101101111100101001100",
15958 => "001111011100101010010100",
15959 => "001100010000111011010110",
15960 => "001001111110111111110100",
15961 => "000100000011111110010001",
15962 => "111100101101010001010111",
15963 => "110110100010000000100100",
15964 => "110010000101001011011010",
15965 => "110001011101110110101000",
15966 => "110100000010001110000100",
15967 => "111000010111001110011000",
15968 => "111101010111111000010100",
15969 => "000001000111100110011011",
15970 => "000100010111011111011000",
15971 => "000111000101000100100101",
15972 => "001000101000111011101111",
15973 => "001011001100000000010101",
15974 => "001110010101000110000010",
15975 => "001111001100110100010110",
15976 => "001101101110010100010000",
15977 => "001100000110000110100000",
15978 => "001010010010010110101101",
15979 => "000110010101111100001111",
15980 => "000000010000011100010001",
15981 => "111000011000111111100100",
15982 => "110000010000110101001000",
15983 => "101010100010100101100000",
15984 => "100101111011010100110000",
15985 => "100010010110101000100011",
15986 => "100010000100100100010111",
15987 => "100010011100001110001011",
15988 => "100010011000000001100111",
15989 => "100100000111011101110011",
15990 => "100110011010000000001010",
15991 => "101001101001111010000010",
15992 => "110000000011010111011100",
15993 => "110111001110001100010000",
15994 => "111100101100011010011110",
15995 => "000000110111111100100011",
15996 => "000100000110000010110010",
15997 => "000110001111110110000010",
15998 => "000110111001011100000100",
15999 => "000101011111001011101000",
16000 => "000010110011100000010011",
16001 => "000000100011010010001000",
16002 => "111110100011000110101011",
16003 => "111011001000001110010000",
16004 => "110110100110110001010110",
16005 => "110010110101000100010000",
16006 => "110000011010010011000110",
16007 => "101111100010100110110000",
16008 => "110000111110101101101110",
16009 => "110011110001100001110100",
16010 => "110110100001111000110110",
16011 => "111010011010011111111110",
16012 => "111111101011000010100111",
16013 => "000100101100101000010111",
16014 => "001001010110100101011011",
16015 => "001101101001011001111010",
16016 => "010000110111100011000110",
16017 => "010010101010010001000010",
16018 => "010010110110110010101110",
16019 => "010001101110111110000010",
16020 => "001111111110111010010100",
16021 => "001110101110111111111110",
16022 => "001110110101111000100010",
16023 => "001111011110000110111000",
16024 => "001111010101110001001000",
16025 => "001110111001111010100010",
16026 => "001111011101011111100110",
16027 => "010000100010010100001100",
16028 => "010000010100011101011000",
16029 => "001110111000011011001100",
16030 => "001110101111010010111000",
16031 => "010000110110111101011110",
16032 => "010011010111111010111010",
16033 => "010101110110110011011100",
16034 => "011000010010111101010001",
16035 => "011000111100100011000100",
16036 => "011000100101000110011111",
16037 => "011000011010011000001011",
16038 => "010111010110001000011010",
16039 => "010110010010100100100010",
16040 => "010101100101111000100000",
16041 => "010010011010111110100110",
16042 => "001011111010011101101101",
16043 => "000011100000000110111101",
16044 => "111010001001010101000111",
16045 => "110000110111011001101000",
16046 => "101001001000001111111110",
16047 => "100011111111011001110100",
16048 => "100001011100011010010000",
16049 => "100000101110101100110111",
16050 => "100000101001101010110010",
16051 => "100000101001110001101000",
16052 => "100001110011110100111100",
16053 => "100100001001111101000011",
16054 => "100110000100000000001011",
16055 => "100111100111010110011101",
16056 => "101001100101101001011110",
16057 => "101011101010011001111010",
16058 => "101110000010011101100000",
16059 => "110000011000011100101100",
16060 => "110001110001001001100110",
16061 => "110011001111101011101000",
16062 => "110101101011110000100100",
16063 => "111000000100101010001111",
16064 => "111010011011101110000000",
16065 => "111100110111111001101010",
16066 => "111101101011000100101111",
16067 => "111100110001001010001010",
16068 => "111011110111011111100010",
16069 => "111010100011111100110000",
16070 => "110111111110000001111011",
16071 => "110101010101011111000011",
16072 => "110011100010001100001000",
16073 => "110001010111010100000000",
16074 => "101110011101001101011010",
16075 => "101101100010100110001110",
16076 => "110000111011110010101010",
16077 => "110111000011101101010100",
16078 => "111101010101110101010000",
16079 => "000011111011100010110001",
16080 => "001100000000110101001110",
16081 => "010011110110101011111010",
16082 => "011000011000100100010100",
16083 => "011001110101010100000111",
16084 => "011010010011001111011001",
16085 => "011010111000110100000000",
16086 => "011011100101010111111011",
16087 => "011010101001110101100001",
16088 => "010110110100100100010110",
16089 => "010001110011111100111110",
16090 => "001101110111100010110100",
16091 => "001011000000100100100100",
16092 => "000111111111010011000001",
16093 => "000100111111001010100000",
16094 => "000011011101010001110101",
16095 => "000011010001001001000010",
16096 => "000010101110011100000010",
16097 => "000001101011010000100110",
16098 => "000001111000010010000100",
16099 => "000011010111011000110100",
16100 => "000100000001001000101101",
16101 => "000011001000100001111011",
16102 => "000000111111110111110010",
16103 => "111100101101011000000000",
16104 => "110110100100110010001100",
16105 => "110010010010100000010100",
16106 => "110010100011101010101010",
16107 => "110101100101011000011110",
16108 => "111001100101001111110100",
16109 => "111110100100101000001110",
16110 => "000010001000110000000000",
16111 => "000001100010011101111010",
16112 => "111111011100101110100101",
16113 => "000000010110110101110010",
16114 => "000011001001100000100001",
16115 => "000011111110100111001100",
16116 => "000011001001101001101100",
16117 => "000011000010000001010100",
16118 => "000011110011001010011011",
16119 => "000100000000111010111010",
16120 => "000010010011110001011100",
16121 => "111111010110111101100101",
16122 => "111101111111100011110001",
16123 => "111111111111011100101101",
16124 => "000011111110001000110001",
16125 => "000110110000000001110000",
16126 => "000110111111110011100110",
16127 => "000110010111100111111100",
16128 => "000110100001011010110001",
16129 => "000111100010101000000100",
16130 => "001000001010010010010111",
16131 => "000111001000011010000110",
16132 => "000101100011110001101101",
16133 => "000101001100111010001100",
16134 => "000101101110100000010001",
16135 => "000100111111001110010100",
16136 => "000000111100110111000001",
16137 => "111010100111101011100101",
16138 => "110011110111011110000100",
16139 => "101100011010111100001100",
16140 => "100110001000101001000100",
16141 => "100100010111001100111001",
16142 => "100101101111100000001001",
16143 => "100111000001110111010111",
16144 => "101000001101100111011000",
16145 => "101010001001010010111010",
16146 => "101101001011000001001000",
16147 => "110010100000010101101110",
16148 => "111010000111110110000010",
16149 => "000001011110011010000100",
16150 => "000110000010101000010000",
16151 => "001000011111101000011001",
16152 => "001011110010010101000100",
16153 => "001111010011000111001110",
16154 => "010000000101011001011100",
16155 => "001111001000111110111010",
16156 => "001110010101001110111010",
16157 => "001101011100110001000010",
16158 => "001100101100100111010100",
16159 => "001011110011110101011111",
16160 => "001010000101001010000100",
16161 => "000111110100000110111011",
16162 => "000110000101010001010010",
16163 => "000110011111001001011010",
16164 => "001000100110001000011100",
16165 => "001010110101100001011110",
16166 => "001110100010011111000100",
16167 => "010011111111101101111100",
16168 => "011000001101011010111001",
16169 => "011001101011100000110001",
16170 => "011000111110111010011111",
16171 => "010111110111110100010110",
16172 => "010111011011010010001110",
16173 => "010110010011011101111000",
16174 => "010101001011001001000010",
16175 => "010100110111000010000010",
16176 => "010010001110101011010000",
16177 => "001100110000100100011100",
16178 => "000110010010111101100011",
16179 => "111110011010111011011000",
16180 => "110110111001110011100001",
16181 => "110000110100011101010010",
16182 => "101001100000100111111010",
16183 => "100011010100101111011110",
16184 => "100010000001100001100101",
16185 => "100010011100001010100011",
16186 => "100010010001111011001111",
16187 => "100011000101111111101111",
16188 => "100101110000111100001001",
16189 => "101011011110011110011110",
16190 => "110011001001000000010010",
16191 => "111000111110000110011101",
16192 => "111011111111100111110001",
16193 => "111100110111000110101111",
16194 => "111011011011000101001110",
16195 => "111000010000010111110100",
16196 => "110100011000110110100000",
16197 => "110000101010101001001000",
16198 => "101101000000000111000000",
16199 => "101000101000001111110110",
16200 => "100101000100100110110011",
16201 => "100100010001100111001001",
16202 => "100100011101001001011101",
16203 => "100100001100000110111011",
16204 => "100100110111110101000111",
16205 => "100110011011111001111011",
16206 => "101000110010000011001110",
16207 => "101101010100110110100000",
16208 => "110011101000100000100110",
16209 => "111010101000100011110110",
16210 => "000001101001110011001100",
16211 => "000111010001100111110110",
16212 => "001011011000010100110100",
16213 => "001111001110000010101000",
16214 => "010011000100000100101110",
16215 => "010101100110100011111000",
16216 => "010110110010100100010000",
16217 => "011001011110111111010011",
16218 => "011101100100100100000011",
16219 => "011111011100001010000111",
16220 => "011111011010100111100111",
16221 => "011111011111011001000101",
16222 => "011110111101110110111111",
16223 => "011101110100110011001011",
16224 => "011100011000000100100110",
16225 => "011010001011011101010111",
16226 => "011000010010000101100001",
16227 => "010110101011100101011010",
16228 => "010011011110111100010110",
16229 => "001111000000000101100110",
16230 => "001011000111101011011110",
16231 => "001000110000001000110000",
16232 => "000111001100110000001101",
16233 => "000100111100011010111101",
16234 => "000010111110100100101110",
16235 => "000011010001001110111100",
16236 => "000100010011000110111110",
16237 => "000011101110110000101111",
16238 => "000001110000110001110110",
16239 => "111110110111101010000000",
16240 => "111010111010010010111011",
16241 => "110110010000011111010010",
16242 => "101111100100111101111000",
16243 => "100110111000110101101000",
16244 => "100010001000111111100100",
16245 => "100010101110001111110010",
16246 => "100010100111000001101100",
16247 => "100001011011100010010110",
16248 => "100001110100000100011010",
16249 => "100010011010011110110100",
16250 => "100011001110011111011001",
16251 => "100100100111111110000111",
16252 => "100100110111100010011011",
16253 => "100101010000010101101111",
16254 => "101000101101111110100110",
16255 => "101101101001001011100110",
16256 => "110000111110010111100100",
16257 => "110010111111110000000100",
16258 => "110101011100101000110110",
16259 => "111001010001011000100010",
16260 => "111101001011010110100101",
16261 => "111111011110110000110010",
16262 => "000001011111110111010010",
16263 => "000101010110000110101100",
16264 => "001011000100001001111111",
16265 => "010000001001101010111100",
16266 => "010010000100001100101010",
16267 => "010001000101110000111100",
16268 => "001110101100010111100100",
16269 => "001100111011111001101110",
16270 => "001100111110101101011100",
16271 => "001100110001001110111100",
16272 => "001011001011100111010100",
16273 => "001010101100011111111100",
16274 => "001101000001000110101010",
16275 => "001111111101010100001010",
16276 => "010001001100011010101110",
16277 => "010001101000010111101100",
16278 => "010010111101101101101100",
16279 => "010101101000011110100110",
16280 => "011000110101000110001011",
16281 => "011011101011110101011011",
16282 => "011101100110100000100011",
16283 => "011110000000101100010011",
16284 => "011101110010000110110101",
16285 => "011100101100110000111011",
16286 => "011001101011111001010111",
16287 => "010111010100110100100100",
16288 => "010111001000001000101000",
16289 => "010110011100010100001100",
16290 => "010100011110010100101000",
16291 => "010011000001010000011000",
16292 => "010010011100010000010110",
16293 => "010001000010111101101100",
16294 => "001101100000000000001010",
16295 => "001000010101001011111111",
16296 => "000010010001010111111111",
16297 => "111011100100101000111111",
16298 => "110101100000100000010000",
16299 => "110000110011110001011010",
16300 => "101100111101101011010110",
16301 => "101011000000011101100010",
16302 => "101011110011010110000110",
16303 => "101110010010000101111010",
16304 => "110010000110010100001000",
16305 => "110111010111111010101101",
16306 => "111101011101101110011010",
16307 => "000011000010110001011101",
16308 => "000110100010010000101000",
16309 => "000111100000101111011110",
16310 => "000110001011010001010110",
16311 => "000010110001000110001110",
16312 => "111110001100110010000010",
16313 => "111000111110010000101100",
16314 => "110010001010111110111110",
16315 => "101001110101001000001110",
16316 => "100011010110011111101101",
16317 => "100001100000000011000000",
16318 => "100010101001101100101010",
16319 => "100101000101110100101001",
16320 => "101001001110010100001010",
16321 => "101110100011101011111000",
16322 => "110011101111110110101100",
16323 => "110111011100011011010000",
16324 => "111000011011011000100010",
16325 => "110111100000110110110110",
16326 => "110110111001101101001100",
16327 => "110111101010100011111100",
16328 => "111001010010110010111000",
16329 => "111010101110101000000001",
16330 => "111100000011110101011010",
16331 => "111101100101000101111100",
16332 => "111101111001010011101101",
16333 => "111011111000101011111010",
16334 => "111000100101010111011110",
16335 => "110101100011001111110000",
16336 => "110011010000011001111000",
16337 => "110001101000100010000010",
16338 => "101111001100011101100010",
16339 => "101010011111001010101000",
16340 => "100110001100001110010101",
16341 => "100100111101110100110001",
16342 => "100110000000111111100011",
16343 => "101000100010010010111010",
16344 => "101100000000110010010110",
16345 => "110000110100000011000100",
16346 => "110111110000000011111111",
16347 => "111111110100110001110000",
16348 => "001000010000100011010010",
16349 => "010000110101010110010000",
16350 => "011000000001010010010011",
16351 => "011100000110010001110001",
16352 => "011101011111100000110011",
16353 => "011101000100100001010011",
16354 => "011001110100101011100110",
16355 => "010100001000110010011110",
16356 => "001110000000000101101000",
16357 => "001000111010011010101100",
16358 => "000110101010000010011101",
16359 => "000110100011101100110010",
16360 => "000110010001000110000010",
16361 => "000110111011101110011010",
16362 => "001010010001000101111010",
16363 => "001111010000010110010110",
16364 => "010100111111010011101100",
16365 => "011001011101110011100011",
16366 => "011010010101110110111101",
16367 => "011001100011000011001111",
16368 => "011000110110001001011111",
16369 => "010111111011101010111000",
16370 => "010111011110111111111100",
16371 => "010110010110110011011100",
16372 => "010011000101001101010100",
16373 => "001110011001110100101110",
16374 => "001001101101111100100110",
16375 => "000110010010100111010000",
16376 => "000011110111011100011101",
16377 => "000000111111000001001011",
16378 => "111100100100111101011000",
16379 => "111000001010110100000001",
16380 => "110101100111001011110000",
16381 => "110011111001010100110010",
16382 => "110000110000111100101100",
16383 => "101001011100010110110110",
16384 => "100010001010010101110111",
16385 => "100001010011001110100001",
16386 => "100001111111110011100001",
16387 => "100001011110110000010011",
16388 => "100010010110011011111001",
16389 => "100011001010010000001011",
16390 => "100011111001100000010011",
16391 => "100100010101101001011111",
16392 => "100100001011100100011111",
16393 => "100100101010001100001001",
16394 => "100101010010010100100001",
16395 => "100110010010001011100001",
16396 => "100111000000011101111000",
16397 => "100111001101101100110100",
16398 => "100111011101000110000011",
16399 => "100111111010101011001010",
16400 => "101010101101011001101000",
16401 => "101110001110010100001100",
16402 => "110000001011111001110010",
16403 => "110010011010110011111010",
16404 => "110110010011101101111111",
16405 => "111100001110110000000110",
16406 => "000001010100000111101111",
16407 => "000011100101101011110010",
16408 => "000101010010010010000100",
16409 => "001000000000000000011000",
16410 => "001100100111101010010110",
16411 => "010000101101101000010000",
16412 => "010001111101100011111110",
16413 => "010010100111000110000110",
16414 => "010011111000001111101000",
16415 => "010101100110010011110000",
16416 => "010110011111110000110100",
16417 => "010110000010010111101010",
16418 => "010110001000001000110000",
16419 => "010110111101111011111100",
16420 => "011001001011000011100101",
16421 => "011100100101000011010001",
16422 => "011101110111001100111000",
16423 => "011101001000011101111011",
16424 => "011100110001110000000000",
16425 => "011100100101011001100111",
16426 => "011100001101100011100101",
16427 => "011011101111000010111011",
16428 => "011010110001000110100101",
16429 => "011001111110010000110101",
16430 => "011001101101011010001100",
16431 => "011001010000011101011101",
16432 => "011000011001001001101001",
16433 => "010111000111101011101000",
16434 => "010110001101100010000010",
16435 => "010101010010001000000000",
16436 => "010010011010000000100000",
16437 => "001110110110011100111100",
16438 => "001011111100101100101110",
16439 => "000111111000011110011110",
16440 => "000010000110111001001101",
16441 => "111011100100010001101010",
16442 => "110100111111000101111100",
16443 => "101111001111110000111110",
16444 => "101010010010011101000000",
16445 => "100101010111011111111101",
16446 => "100010001000110100111100",
16447 => "100010010001101101101111",
16448 => "100010110101011101010101",
16449 => "100010001010110011111111",
16450 => "100011010011011010011111",
16451 => "100110111110001100001111",
16452 => "101010101001001101100110",
16453 => "101100111101001100100010",
16454 => "101101110100011010100110",
16455 => "101100010000110000011110",
16456 => "101000110010100011001110",
16457 => "100110100001100011100001",
16458 => "100101010011010110000001",
16459 => "100011100110011100101111",
16460 => "100011111000010011011110",
16461 => "100110110000111111101101",
16462 => "101001111110110111001100",
16463 => "101101110011000111011110",
16464 => "110010010000100101000110",
16465 => "110101001100000100011110",
16466 => "110110001101100111000100",
16467 => "110110111011101100101000",
16468 => "110111111001011110011010",
16469 => "111000101111111111100100",
16470 => "111001110010001011110110",
16471 => "111011000111111001000110",
16472 => "111011111100100011011001",
16473 => "111011000001101111111101",
16474 => "111001000110110000011110",
16475 => "111010110101001111010000",
16476 => "000000100101001100000100",
16477 => "000011110000110001000010",
16478 => "000100111010010101110110",
16479 => "001001011000010000110101",
16480 => "001101111110101000001110",
16481 => "001110100000100001011010",
16482 => "001101000101001001010000",
16483 => "001100000010100101001100",
16484 => "001011100011110011011110",
16485 => "001011011110001010100000",
16486 => "001011001101111001001000",
16487 => "001001111111000111110100",
16488 => "001000101111010011000111",
16489 => "001000111000101000111000",
16490 => "001001011100111011011010",
16491 => "001001101010111101100110",
16492 => "001011000110100101011010",
16493 => "001110110110000011001110",
16494 => "010011001111110000100010",
16495 => "010101100111001000000000",
16496 => "010101110011010001000110",
16497 => "010110001110110101111110",
16498 => "010111000000110111101000",
16499 => "010110001100100111111100",
16500 => "010100110101110001110100",
16501 => "010100001101011010100110",
16502 => "010100001001001000111010",
16503 => "010101101101100011001110",
16504 => "010111100110100011011110",
16505 => "010111101010100101010100",
16506 => "010111000111110110110010",
16507 => "010110110000001000011010",
16508 => "010101111110000101100100",
16509 => "010100111110100100101010",
16510 => "010010110010101111111110",
16511 => "001101001100111000000100",
16512 => "000110110011111001000001",
16513 => "000011100001100011110011",
16514 => "111111100000011101010001",
16515 => "111000100100111011100011",
16516 => "110011100010111100101010",
16517 => "110001100100000001000100",
16518 => "101111100000111000111010",
16519 => "101100011100111110001110",
16520 => "101011000101101110011010",
16521 => "101101001001000110110100",
16522 => "110000010001100100111100",
16523 => "110001001100110111000010",
16524 => "101101010001011101000110",
16525 => "100110100011101111110001",
16526 => "100010111011001001010111",
16527 => "100011000110111101111101",
16528 => "100011111101101010100101",
16529 => "100100011001001011110010",
16530 => "100101001001110010101111",
16531 => "100110000101100010110101",
16532 => "100110100011100010011110",
16533 => "100111001001110110100010",
16534 => "100111100110110110101011",
16535 => "100111110100100010010011",
16536 => "101010000010110010100000",
16537 => "101111010000001110110010",
16538 => "110100100101111101111010",
16539 => "110111111001100011000110",
16540 => "111010111100110011001010",
16541 => "111110000101110000101010",
16542 => "000000110001110001000001",
16543 => "000100000111100011001001",
16544 => "000110111111011110110110",
16545 => "001001111001101100111100",
16546 => "001110001000000110000110",
16547 => "010001000001000110110000",
16548 => "010001011100001001101110",
16549 => "010000001011010010010010",
16550 => "001110101010100000110100",
16551 => "001110010110010100111100",
16552 => "001101011110111010010010",
16553 => "001011010101100011101000",
16554 => "001001111101000111101100",
16555 => "001010101110001110111000",
16556 => "001100010011101100110000",
16557 => "001011101010000111001011",
16558 => "001001100000100111001001",
16559 => "001000010111011100010110",
16560 => "001000011011010111110011",
16561 => "001010010000010111101001",
16562 => "001101001111100100100110",
16563 => "010000101001110010101100",
16564 => "010101111011010110101010",
16565 => "011010101111000011011000",
16566 => "011011011100000000101011",
16567 => "011010000111101000000111",
16568 => "011001001000100001110011",
16569 => "011000000010110010100011",
16570 => "010111000111000110011000",
16571 => "010110010101111010010110",
16572 => "010100100000001111100100",
16573 => "001111111011000010010010",
16574 => "001001000101111100000000",
16575 => "000010000100000011100011",
16576 => "111001100101111011011110",
16577 => "101111111011101101010110",
16578 => "101000101001100111101000",
16579 => "100100000001110110000000",
16580 => "100001110111100000101011",
16581 => "100001101011110110110011",
16582 => "100001010101011011111001",
16583 => "100001010100110011100010",
16584 => "100001100010011111011100",
16585 => "100010101101110111101110",
16586 => "101000101111111010010000",
16587 => "110001111010111001101010",
16588 => "111001101101100101100101",
16589 => "000000100100110011100000",
16590 => "000111001101010101010111",
16591 => "001011000001110000011111",
16592 => "001010110000011110101100",
16593 => "001001001101100101001110",
16594 => "001000010010010010110010",
16595 => "000110110000001100000100",
16596 => "000100001001100110010000",
16597 => "000001001100011100011010",
16598 => "111110010010001011011011",
16599 => "111011000110011001100001",
16600 => "111000001010000011000110",
16601 => "110110001101111010001100",
16602 => "110011110011101111100110",
16603 => "110001101000010001011110",
16604 => "110010101100010111110000",
16605 => "110101011100110100000001",
16606 => "110110010101101111101100",
16607 => "110110010101100001010100",
16608 => "111000100111011110000010",
16609 => "111100100111101110101011",
16610 => "000000000011001101101100",
16611 => "000010100100101110110111",
16612 => "000011011111110110100110",
16613 => "000010000111000111110000",
16614 => "111111001010101000110101",
16615 => "111100000101100001001100",
16616 => "111001100011001101011101",
16617 => "110110100001011100110111",
16618 => "110100000010011010110001",
16619 => "110100000011101000000011",
16620 => "110100100110100001100000",
16621 => "110100000101100010111011",
16622 => "110100011100101100110000",
16623 => "110111000001100001101110",
16624 => "111010011010111001111111",
16625 => "111101110101100001001101",
16626 => "000010011000101110000000",
16627 => "000111001010101000111100",
16628 => "001010100111001111101110",
16629 => "001101100100011010111000",
16630 => "010000001110100101010100",
16631 => "010001100010100001101100",
16632 => "010001010110110011101100",
16633 => "010001000111101010011110",
16634 => "010010100000010111111010",
16635 => "010011111010000001001110",
16636 => "010011010000001100001010",
16637 => "010010110001011110011000",
16638 => "010011100111010010001000",
16639 => "010011001111100111010000",
16640 => "010001000101000101101010",
16641 => "001111010000110100101010",
16642 => "001110101101111100101000",
16643 => "001101010011011100011100",
16644 => "001010101101010110100110",
16645 => "001001110000111111001110",
16646 => "001010010110011110011101",
16647 => "001011011101111001010100",
16648 => "001100001000001111010100",
16649 => "001010011110000111010000",
16650 => "001000010110011111111011",
16651 => "000111000000110000111111",
16652 => "000101011110010011110110",
16653 => "000011001000100011000000",
16654 => "111110011110001101110101",
16655 => "111000111101000101101100",
16656 => "110100001011011000010000",
16657 => "101111010111000101011000",
16658 => "101011100000010111010110",
16659 => "101001000001010010101010",
16660 => "100111100010000000110111",
16661 => "100110111011111000100101",
16662 => "101000000101011000001100",
16663 => "101010101000111000101100",
16664 => "101001110001100000100000",
16665 => "100110010101101011010110",
16666 => "100101111011110101011101",
16667 => "100111000011010010011101",
16668 => "100111010100011011110111",
16669 => "100111101010111100001000",
16670 => "100111111010111110011111",
16671 => "101000001010100000101110",
16672 => "101000110100011011010110",
16673 => "101001000010111011010110",
16674 => "101001010110011101011100",
16675 => "101100100110001110100110",
16676 => "110011000100110010001100",
16677 => "111001111110101000101011",
16678 => "000000011101111110111011",
16679 => "000111110001001001010100",
16680 => "001111110010001101100110",
16681 => "010110001011100110001100",
16682 => "011001100000001010000111",
16683 => "011010101000100010101011",
16684 => "011010101101001011110101",
16685 => "011010111100101001110001",
16686 => "011011101100100001000001",
16687 => "011011101000001110110101",
16688 => "011010000011111001110000",
16689 => "010111011100101111010000",
16690 => "010101011010010111111000",
16691 => "010101110011111101111110",
16692 => "010111010100100011010010",
16693 => "010111101110011001010000",
16694 => "011000010000111101010011",
16695 => "011010000000101010111001",
16696 => "011011000100110101111101",
16697 => "011010010110011001110001",
16698 => "011001100010001101011011",
16699 => "011001010111100010000011",
16700 => "011000100111101111000011",
16701 => "011000001010010100110001",
16702 => "010111100010111001100010",
16703 => "010100110100001000001000",
16704 => "010001101011000000101100",
16705 => "001101110011000101110000",
16706 => "000110110111011011011001",
16707 => "111101111110001010111000",
16708 => "110110011011011011000100",
16709 => "110001001000110000011010",
16710 => "101001100110010100010100",
16711 => "100010001000101011010011",
16712 => "100001000101001100001000",
16713 => "100001110100111001001101",
16714 => "100001100010101110111011",
16715 => "100001111110110110100101",
16716 => "100001110100011000001001",
16717 => "100001100100001001111101",
16718 => "100001100101101110101011",
16719 => "100010001111100010101101",
16720 => "100010111011000011000111",
16721 => "100010110111110111000100",
16722 => "100101000001111000110001",
16723 => "101001010010011001101110",
16724 => "101110001010000111111010",
16725 => "110010010111101011110110",
16726 => "110100010100001001010100",
16727 => "110110110111010100111011",
16728 => "111010111001010100011110",
16729 => "111110000110101101111001",
16730 => "111111101010011011011001",
16731 => "111111110100110011111011",
16732 => "111111111000011100010101",
16733 => "111111011111110000101010",
16734 => "111110010100101111010000",
16735 => "111100101010100100011110",
16736 => "111011010110011000110101",
16737 => "111100011001001111001010",
16738 => "111110100101010000111111",
16739 => "000000011001001101011001",
16740 => "000010011111110011101000",
16741 => "000110111110100001011100",
16742 => "001111000111111111000000",
16743 => "010110011011001110000010",
16744 => "011010110001011101110001",
16745 => "011101111010011110001111",
16746 => "011110101111000010110101",
16747 => "011110100101111011100001",
16748 => "011110111010010101111101",
16749 => "011110010110110101100000",
16750 => "011101011000101101011111",
16751 => "011011101100101011001110",
16752 => "011000000100011100001011",
16753 => "010011001011000100010000",
16754 => "001101110100110011000100",
16755 => "000111001001101001100101",
16756 => "111111000111001100001000",
16757 => "111000011101111101011001",
16758 => "110100110101000110000111",
16759 => "110011101011110111100110",
16760 => "110100101100110111100101",
16761 => "110110100100011010001100",
16762 => "111000000001110001100100",
16763 => "111010011001111111001110",
16764 => "111110101111001111000011",
16765 => "000010111000100110011101",
16766 => "000100111010110100000010",
16767 => "000110001010110111111100",
16768 => "001000101110101011001010",
16769 => "001011110001110010001110",
16770 => "001100100001110000000100",
16771 => "001001111001001001010110",
16772 => "000100000000100101111100",
16773 => "111011100101001011110110",
16774 => "110011011010010100111000",
16775 => "101100110011010000010100",
16776 => "100110101101010111100101",
16777 => "100010100110000001011111",
16778 => "100001011000001111011001",
16779 => "100010001011111111001101",
16780 => "100110001111010001010001",
16781 => "101100000010110011011000",
16782 => "110001011001000000111100",
16783 => "111000011011110000101110",
16784 => "000000011110100110110100",
16785 => "000111000011100100000011",
16786 => "001100011001110011000010",
16787 => "010000101011011101000010",
16788 => "010011101001100011001000",
16789 => "010011110000110111101110",
16790 => "010000100011101111000110",
16791 => "001100000010011000010100",
16792 => "000111001001010010100100",
16793 => "000010001101100011011000",
16794 => "111101100110000101101000",
16795 => "111001111111000110001000",
16796 => "110110110110111100010000",
16797 => "110010111100000001010010",
16798 => "101111110000101001110100",
16799 => "101110001111001000000000",
16800 => "101101001111011011010110",
16801 => "101011111011111011000110",
16802 => "101011100100101111100010",
16803 => "101101010111110100100000",
16804 => "101101000011110000110110",
16805 => "101001100100111101001100",
16806 => "101000010010110001100110",
16807 => "101001011010011100011110",
16808 => "101010100111101001100000",
16809 => "101101110000110100111100",
16810 => "110100111010010010000010",
16811 => "111101111010001100000100",
16812 => "000100111101100100001000",
16813 => "001000101110111110000111",
16814 => "001001011110001000001100",
16815 => "001001011000110101001100",
16816 => "001010000001110110111111",
16817 => "001001110000000010011010",
16818 => "001000010110011111111110",
16819 => "000111110010010101001010",
16820 => "001001011111011111001010",
16821 => "001100011110000110101010",
16822 => "001110100001111101101100",
16823 => "010000110010010001001100",
16824 => "010101100010111111011010",
16825 => "011010001001000101110101",
16826 => "011010101011010110011011",
16827 => "011001110001101011001010",
16828 => "011001110110000100101111",
16829 => "011001010100001101010111",
16830 => "011000111111110110010011",
16831 => "011000110001100111100111",
16832 => "011000001011011101111100",
16833 => "010111110101110111100110",
16834 => "010101110110001000011000",
16835 => "010011010001010010001100",
16836 => "010011001111011000000110",
16837 => "010100001100010011000110",
16838 => "010010100000010010110110",
16839 => "001110110101000000110110",
16840 => "001100011110000100001110",
16841 => "001010111100111110110111",
16842 => "001000011000011100001000",
16843 => "000010111100011100100010",
16844 => "111011101111101000011111",
16845 => "110101001010001011001110",
16846 => "101011001110000111101110",
16847 => "100001110011000111111011",
16848 => "100000101101111100001001",
16849 => "100001111011001011000001",
16850 => "100001110010111011000001",
16851 => "100010011011111010011001",
16852 => "100010100101111100001101",
16853 => "100010101000000111111111",
16854 => "100011101101010110100101",
16855 => "100111110100100000000011",
16856 => "101110100000111110000110",
16857 => "110100000010111011101100",
16858 => "110110100100110100101111",
16859 => "110101101101011000100110",
16860 => "110100001011110010000100",
16861 => "110010111110000000100100",
16862 => "101111010110011001000110",
16863 => "101010011000111110101110",
16864 => "100110011110100010001000",
16865 => "100100100000101110001111",
16866 => "100100000111110000111101",
16867 => "100100010110110001000001",
16868 => "100101000101110010001111",
16869 => "100101111101110011001001",
16870 => "100111100111110001101111",
16871 => "101010000100011011111100",
16872 => "101100100110010100010110",
16873 => "101111011000000101000110",
16874 => "110001101001011100001000",
16875 => "110100101101001101111111",
16876 => "111010001101000001110111",
16877 => "000000100010111011000101",
16878 => "000110110010011110000100",
16879 => "001101100000111011011110",
16880 => "010100110111111100001100",
16881 => "011011000010100111011011",
16882 => "011101111011100111111001",
16883 => "011110000000010100011101",
16884 => "011101010111110111111011",
16885 => "011110001011011110001001",
16886 => "011101110111000100000111",
16887 => "011000100001101010101101",
16888 => "010001101001010001111010",
16889 => "001100111010111111111100",
16890 => "001000110101111000001001",
16891 => "000100100111111000101110",
16892 => "000001001110011101000100",
16893 => "111111101001000000011001",
16894 => "111111101100000111110101",
16895 => "111111110011110110101000",
16896 => "111111101010010000001011",
16897 => "000000101110000100100101",
16898 => "000011100011101001010100",
16899 => "000110010110100001010100",
16900 => "001000010100001010111011",
16901 => "001010101101110000001010",
16902 => "001101101100111001110000",
16903 => "010000111011110010101010",
16904 => "010011110100000110010100",
16905 => "010100110011001111001000",
16906 => "010011001010011011110000",
16907 => "001111110011001000101100",
16908 => "001100101101110100110010",
16909 => "001001110100000000100111",
16910 => "000101100100111111000001",
16911 => "000001011000111010100011",
16912 => "111110011100111100111100",
16913 => "111100000101001000111001",
16914 => "111010001110011110001010",
16915 => "111000110110110000101100",
16916 => "110111101101010010101111",
16917 => "110111010110010010011110",
16918 => "111001000001100010101100",
16919 => "111011110111000110101101",
16920 => "111101111010011100001011",
16921 => "111111111011000101010110",
16922 => "000010011011100011001000",
16923 => "000101000010000000101110",
16924 => "000111110001111111011110",
16925 => "001010001110111101011110",
16926 => "001100101000011000001100",
16927 => "001110100100010010100100",
16928 => "001111100000111001101100",
16929 => "001111100010100000111100",
16930 => "001100001100001111110100",
16931 => "000100100000011010111101",
16932 => "111011101101110111110110",
16933 => "110100011111100000000100",
16934 => "101110011100011111000110",
16935 => "101000011011011010111000",
16936 => "100100110101001110111100",
16937 => "100101111110011011000101",
16938 => "101000100001101110001000",
16939 => "101001111110111100100000",
16940 => "101101000101101110010010",
16941 => "110011000101110100111000",
16942 => "111001101011001011010100",
16943 => "111111001111001001111001",
16944 => "000010011010111111011010",
16945 => "000010011001100100001001",
16946 => "000000111111100000111110",
16947 => "111111100111010111100000",
16948 => "111110000111000000111010",
16949 => "111100100010101000010001",
16950 => "111011101101011111001011",
16951 => "111100110000100010010110",
16952 => "111110100000000000000011",
16953 => "111111001000000100100011",
16954 => "111111110110111001100111",
16955 => "000010001111100000111000",
16956 => "000110010101011010111110",
16957 => "001011001111111000110010",
16958 => "001111001110010100100010",
16959 => "010001101000010001001110",
16960 => "010011010101110110111010",
16961 => "010101010100011111111000",
16962 => "010111101111110100010100",
16963 => "011001001100011110100111",
16964 => "011000111000101111110101",
16965 => "011000010100111111011011",
16966 => "011000001101111010101110",
16967 => "010111110010010011011010",
16968 => "010110111001001001011000",
16969 => "010110000101000100101000",
16970 => "010101100000100111100110",
16971 => "010100111000111110011010",
16972 => "010100111011100100111010",
16973 => "010100100101001101111000",
16974 => "001111101110000011110110",
16975 => "000111000011001010111001",
16976 => "111110110101010010110101",
16977 => "110110010110100110011100",
16978 => "101101010001010010011110",
16979 => "100111010010001010110011",
16980 => "100100110011001000000001",
16981 => "100011101000001101011101",
16982 => "100100000000110000001100",
16983 => "100111000110111000111111",
16984 => "101101000011010100111010",
16985 => "110011111001000000011010",
16986 => "111000010111111100110010",
16987 => "111001100110000001011000",
16988 => "111001000010011100100011",
16989 => "111000000010101010101100",
16990 => "110110101111110011110101",
16991 => "110100010100100010100001",
16992 => "101111110101111000101100",
16993 => "101001110010111111101000",
16994 => "100101000100010111110011",
16995 => "100011001100010010010010",
16996 => "100010100101101111111111",
16997 => "100010111111001101010111",
16998 => "100100111000010000010111",
16999 => "100111101101101000100111",
17000 => "101010111100011010100100",
17001 => "101100010110110101010000",
17002 => "101010011010111110111010",
17003 => "101000000001110101110100",
17004 => "100111110100000101101001",
17005 => "101000101001000011100110",
17006 => "101001001101100101110000",
17007 => "101001101000000100101010",
17008 => "101011000111010100011000",
17009 => "101111101101100011001110",
17010 => "110110111010110000010101",
17011 => "111110110111100011110010",
17012 => "000110111011010010111011",
17013 => "001110010110000110100100",
17014 => "010101100000111101000010",
17015 => "011011110100101100000001",
17016 => "011110101111011011100011",
17017 => "011111000010111100110100",
17018 => "011111000000100111001111",
17019 => "011111011010001101111001",
17020 => "011111000010010010100110",
17021 => "011010111101111000110000",
17022 => "010100011001110111100010",
17023 => "001111011001010111110100",
17024 => "001100010100010000101010",
17025 => "001001110101000110001000",
17026 => "000111010100010100100010",
17027 => "000100001001100110100001",
17028 => "000001000100101011110111",
17029 => "111111101010000110101000",
17030 => "111111001011010101010010",
17031 => "111110011100110001001111",
17032 => "111110001001011001100011",
17033 => "111110100011011010110110",
17034 => "111111100111101011000101",
17035 => "000000110001000100111001",
17036 => "000000111011101001111001",
17037 => "000001000111011010010100",
17038 => "000001001111111000010111",
17039 => "111111010010000000000000",
17040 => "111100001001000110100000",
17041 => "111010000011000111101010",
17042 => "111000100001000010111010",
17043 => "110101111110011001011000",
17044 => "110010110101001010111000",
17045 => "110000101111111100000000",
17046 => "101111011110010110101000",
17047 => "101101110111010111010100",
17048 => "101100100101101111100010",
17049 => "101100100000111100101000",
17050 => "101100111111011011110110",
17051 => "101101101011011010101000",
17052 => "101111100011011101001010",
17053 => "110010000101001100000100",
17054 => "110011010011101010111010",
17055 => "110011101111101111100000",
17056 => "110101010000111000001110",
17057 => "111000100000011010001110",
17058 => "111101001011101011100000",
17059 => "000010001010000010000000",
17060 => "000110000100000100110010",
17061 => "001000000101000011000001",
17062 => "001001011101100100111010",
17063 => "001100001010111110010000",
17064 => "001110110110111101110110",
17065 => "010000001010000101000100",
17066 => "010001101001011001010010",
17067 => "010100001001110100000100",
17068 => "010110010101001000011010",
17069 => "010110111100110010100000",
17070 => "010110101010010101001100",
17071 => "010101101100100100001000",
17072 => "010011011110100010101010",
17073 => "010001011100010010101010",
17074 => "010001010000111001101110",
17075 => "010010100011000001010110",
17076 => "010011100100111011010110",
17077 => "010100101100010111110110",
17078 => "010111100100100101110110",
17079 => "011001110110011111100001",
17080 => "011000110101100101101001",
17081 => "010101110110111100101010",
17082 => "010011101010010000101010",
17083 => "010010111101101001001010",
17084 => "010000011100011011011100",
17085 => "001001111101010101110110",
17086 => "000001011110110010111011",
17087 => "111010001111110111110011",
17088 => "110110011110111100110000",
17089 => "110101001000000010100000",
17090 => "110101000101011001011100",
17091 => "110101011000010010110000",
17092 => "110100000010100010110110",
17093 => "110001101100011001100110",
17094 => "101110110110100100001100",
17095 => "101100110000000000001100",
17096 => "101110010100101000111110",
17097 => "110011001100111010110000",
17098 => "111001000000010000111000",
17099 => "111101111011000010100101",
17100 => "000011000100010111110001",
17101 => "001001011101011010110100",
17102 => "001101110110110111101100",
17103 => "010000001110111101000100",
17104 => "010011110010101001000110",
17105 => "010111011010101111001100",
17106 => "011000010000100110010001",
17107 => "010111011111110010110100",
17108 => "010110111001011100100100",
17109 => "010001110001000010100000",
17110 => "000101011001111000110010",
17111 => "111000101100010111000110",
17112 => "110000001110111000000100",
17113 => "101001101000100010000110",
17114 => "100100001100100100111111",
17115 => "100001111001101000011101",
17116 => "100010001010100100010101",
17117 => "100010111100001001001001",
17118 => "100100010000101011111011",
17119 => "100111011011000001010101",
17120 => "101101000101111111001000",
17121 => "110100000000010101001000",
17122 => "111011010001000010010000",
17123 => "000100000101110011011001",
17124 => "001101101110011100111010",
17125 => "010101001000001000101110",
17126 => "010111111001100000010000",
17127 => "010101100011110100001010",
17128 => "010000010110111110111000",
17129 => "001011111001011000110011",
17130 => "001001110011101101001011",
17131 => "000111100101100110110000",
17132 => "000010110011111111101010",
17133 => "111100111100010011111010",
17134 => "110110111000110110000000",
17135 => "101111011000101100100000",
17136 => "100111011100111000110101",
17137 => "100010111000111001010111",
17138 => "100010110001010101010010",
17139 => "100100001110000111101001",
17140 => "100110001001010101100001",
17141 => "101010010111101011010000",
17142 => "110001000100110011100100",
17143 => "110111000111111101100010",
17144 => "111011010001000000000001",
17145 => "000000101011111111010001",
17146 => "000111111101000010000000",
17147 => "001101111101110111010100",
17148 => "010001110100011001101100",
17149 => "010100011000110100000010",
17150 => "010101101110111010101110",
17151 => "010100110001111000100010",
17152 => "010001000111100011010000",
17153 => "001100001101000000010110",
17154 => "000111101010000001001111",
17155 => "000100001111010100010001",
17156 => "000001110000110001001001",
17157 => "000000010001101111000001",
17158 => "000001000010100111000111",
17159 => "000100000010100000110101",
17160 => "000111000011011010101111",
17161 => "001000011010101110010000",
17162 => "001000100101001110011011",
17163 => "001001000000100000010111",
17164 => "001010001000001100001001",
17165 => "001010101110110010101010",
17166 => "001001110000111101010011",
17167 => "000111001111111010010101",
17168 => "000100001001010110000001",
17169 => "000010100111011001111101",
17170 => "000011101011101110011101",
17171 => "000101110001111100111010",
17172 => "000111010010111000011110",
17173 => "000111111100110111001111",
17174 => "001000010001111100100110",
17175 => "001000100010100010000011",
17176 => "000111100111100101101100",
17177 => "000100101000000101100001",
17178 => "000000111100001110101010",
17179 => "111110000110000001001111",
17180 => "111011001100110110111110",
17181 => "110110110110000011011011",
17182 => "110001010000011010101110",
17183 => "101100000111011111001100",
17184 => "101000010110101111110100",
17185 => "100100101010101111001001",
17186 => "100001011011110111001001",
17187 => "100001001101011001100110",
17188 => "100010111111011101001111",
17189 => "100100000001011000000011",
17190 => "100100100011010100100001",
17191 => "100101001011000010100000",
17192 => "100101110100001100100111",
17193 => "101000000101101010000110",
17194 => "101100000101110000010010",
17195 => "101111100111111110001110",
17196 => "110010110001110110001010",
17197 => "110110011010110001100110",
17198 => "111010010011001111001110",
17199 => "111110101110100011110011",
17200 => "000010101111010000001011",
17201 => "000100100010100011011100",
17202 => "000100100111001100000001",
17203 => "000100110011000010110110",
17204 => "000101011011010100001101",
17205 => "000101010111000101100001",
17206 => "000101001000100100100110",
17207 => "000110100101111110011000",
17208 => "001001011001100100110010",
17209 => "001011101100000110100100",
17210 => "001100111111001101001010",
17211 => "001101111000100001111010",
17212 => "001110100001000110000010",
17213 => "001111001100010100011110",
17214 => "010000010011010110101000",
17215 => "010001101000001010000100",
17216 => "010010110101010010101010",
17217 => "010011101111110001000110",
17218 => "010100101110010000000100",
17219 => "010101101100110100100100",
17220 => "010110000101000011110000",
17221 => "010110000100110101101000",
17222 => "010101110010111100011100",
17223 => "010101110111000001011100",
17224 => "010110100110101010100000",
17225 => "010100111101101010110110",
17226 => "001110101111111011000000",
17227 => "000110111110100010101010",
17228 => "000001100111001001001110",
17229 => "111111011101001101111001",
17230 => "111111101001001110111100",
17231 => "000010011000010001111001",
17232 => "000111100110111010010111",
17233 => "001100000110110011011110",
17234 => "001100101101010000100110",
17235 => "001011010011000000010010",
17236 => "001011011100001001000001",
17237 => "001101001000111111001010",
17238 => "001110000110100100111110",
17239 => "001101001011100001000010",
17240 => "001100010101101011010110",
17241 => "001101000010001100000110",
17242 => "001100010100010010100010",
17243 => "001000010000000000100010",
17244 => "000010110011100100010011",
17245 => "111110001100000110111010",
17246 => "111011011101100010001001",
17247 => "111000100111011011010001",
17248 => "110011000000011101110000",
17249 => "101100111011111100111010",
17250 => "101000101100111000000110",
17251 => "100100111101001011100111",
17252 => "100010001101010101110101",
17253 => "100001100011100010011111",
17254 => "100001100000010110010011",
17255 => "100001010101001000011111",
17256 => "100001011000111100101000",
17257 => "100010011101000110110100",
17258 => "100101011010010111100111",
17259 => "101000010111000000100010",
17260 => "101010001001010111101010",
17261 => "101101011010001100011100",
17262 => "110010110111011010101010",
17263 => "111000101111011001011100",
17264 => "111110000101000010011000",
17265 => "000010010001010111010011",
17266 => "000101001000001000000101",
17267 => "000101001110001000101011",
17268 => "000000011101101010010100",
17269 => "111001011010000100110000",
17270 => "110100111100100111010001",
17271 => "110011100000001000000100",
17272 => "110001101111110111010100",
17273 => "101110101001010001100010",
17274 => "101101010101110011000010",
17275 => "101111011101101110010100",
17276 => "110010100111111110001100",
17277 => "110101001101101100011001",
17278 => "111000011101100000000000",
17279 => "111101110101111110111110",
17280 => "000011101101111111011010",
17281 => "000110110001110100001100",
17282 => "000111111010110011100111",
17283 => "001010010010100101100001",
17284 => "001101001101111100101110",
17285 => "001110111000001110111100",
17286 => "010000000100010110100100",
17287 => "010001011000101000010000",
17288 => "010010010101100101110110",
17289 => "010011011001001101101000",
17290 => "010101000000110001010000",
17291 => "010110111101011010101010",
17292 => "011000011011101101111001",
17293 => "011000000111100011110001",
17294 => "010110000001101100010110",
17295 => "010010110000110100111110",
17296 => "001110101010101100100000",
17297 => "001010110111010001110001",
17298 => "001000000010101111100100",
17299 => "000110110110101000110111",
17300 => "001000000011110011111011",
17301 => "001010100001100110101011",
17302 => "001100100111110010111110",
17303 => "001110100000000011010010",
17304 => "010001011001011010100100",
17305 => "010100001001111010110000",
17306 => "010011001110001110000010",
17307 => "001110001001111110001110",
17308 => "000111011100101000011010",
17309 => "000000000110001000110011",
17310 => "110111111100011000010100",
17311 => "110000000110001001000010",
17312 => "101010001100111011001010",
17313 => "100101110111100010110111",
17314 => "100010101010010111010111",
17315 => "100001011100110011110011",
17316 => "100001001100111110100111",
17317 => "100001000000111111010001",
17318 => "100010001001110000101011",
17319 => "100100101001010100111011",
17320 => "100110111100001000011111",
17321 => "101000000011101111011000",
17322 => "101000010101001101111000",
17323 => "101000001111101000010100",
17324 => "100111011001101110010110",
17325 => "100110010000001011100001",
17326 => "100110001111010011001101",
17327 => "100111010110000110101001",
17328 => "101000010111110011111110",
17329 => "101001000110010011001110",
17330 => "101001101010001001000110",
17331 => "101010001001101000001100",
17332 => "101100111011110101101110",
17333 => "110011100110101010110110",
17334 => "111011010010111011000011",
17335 => "000001111111001111111101",
17336 => "001000011110111111011110",
17337 => "001110010010100010110100",
17338 => "010010100001111101101000",
17339 => "010101110011000010100110",
17340 => "011001001001001001011001",
17341 => "011100010100010101010100",
17342 => "011101100100000111100000",
17343 => "011101001101011010010101",
17344 => "011101000101100000101110",
17345 => "011100101110101010100111",
17346 => "011011011011111100100011",
17347 => "011001111100101101001101",
17348 => "011001011000101010110101",
17349 => "011010000111111101101110",
17350 => "011001111101001100001010",
17351 => "010111010111000000100100",
17352 => "010100011111111001110010",
17353 => "010010110011011010110010",
17354 => "010001000110000001110100",
17355 => "001110101011111111100010",
17356 => "001100101101011000111010",
17357 => "001100011000100111100100",
17358 => "001101011000101011000000",
17359 => "001110100110110111000100",
17360 => "001110111010011110000110",
17361 => "001101100001110011111010",
17362 => "001011000001000001100010",
17363 => "001000111111001111100101",
17364 => "001000011100110100110001",
17365 => "001000000001011110110111",
17366 => "000100100000010001100101",
17367 => "111100110011101001101001",
17368 => "110100100111110100101100",
17369 => "101111110011111110000000",
17370 => "101101010110000100111000",
17371 => "101100000001001110010110",
17372 => "101101000010010011100110",
17373 => "101111001100111110111100",
17374 => "110000001011001100110110",
17375 => "101111001101110001000110",
17376 => "101100000010100100000010",
17377 => "101000001110001011111100",
17378 => "100111000001010001100110",
17379 => "101000010101111111010000",
17380 => "101000110001100000110000",
17381 => "101000101111111110101000",
17382 => "101011011110110101101000",
17383 => "101111111000111101100110",
17384 => "110011111001110011001110",
17385 => "111000101001110111010001",
17386 => "111111100111101111001110",
17387 => "001000010001111111000110",
17388 => "010000010000100100100110",
17389 => "010110011101000110110000",
17390 => "011010111011101101100000",
17391 => "011011111100010011011011",
17392 => "011001100100010100101011",
17393 => "010111001110101111001100",
17394 => "010101100101000001011000",
17395 => "010001111011111011101010",
17396 => "001101000000111011010100",
17397 => "001010011100110001001101",
17398 => "001001011011100101000011",
17399 => "000110001100001100100010",
17400 => "000000101100011110111000",
17401 => "111011001011001100000010",
17402 => "110110101110001001001111",
17403 => "110100111000110001110110",
17404 => "110111001110100110101101",
17405 => "111011110001111000100110",
17406 => "111111001011001011000110",
17407 => "000001011011110000101110",
17408 => "000100000100010000110000",
17409 => "000110000111010110100110",
17410 => "000110010101100000011110",
17411 => "000110010100000111101100",
17412 => "000111000100000110110011",
17413 => "000110001101111110110110",
17414 => "000001101100001110100010",
17415 => "111011000100010101000100",
17416 => "110101001111100001011000",
17417 => "101111111000111010111010",
17418 => "101010011010100001000110",
17419 => "100110111100110010100010",
17420 => "100101000100110111010111",
17421 => "100011011000101101110011",
17422 => "100010110011000101001111",
17423 => "100011000010101000101111",
17424 => "100100010011110010111011",
17425 => "100111110000111001110110",
17426 => "101101011010011010000110",
17427 => "110101010111101001011100",
17428 => "111110000010011001010110",
17429 => "000100100101100100101011",
17430 => "001001011011111000010011",
17431 => "001110101010001011111100",
17432 => "010010010001001100010010",
17433 => "010001101101110000110000",
17434 => "010000011011110110111110",
17435 => "010000100100010000011100",
17436 => "001111110101000011111110",
17437 => "001110010110011011000000",
17438 => "001100111011111100101000",
17439 => "001011101010010110010111",
17440 => "001010100011011000101101",
17441 => "001001010010101110100010",
17442 => "001000100010111111011011",
17443 => "000111000010101011010110",
17444 => "000100110110000111010100",
17445 => "000101110100001111010000",
17446 => "001000101101001101100011",
17447 => "001000110010100100100010",
17448 => "000101111100100000110010",
17449 => "000010111011000011001000",
17450 => "000001010001101101101101",
17451 => "000000100011100001101100",
17452 => "111111110110110111000111",
17453 => "111110110111000101001110",
17454 => "111101100111001101100110",
17455 => "111100000000110110100100",
17456 => "111001100110110000010110",
17457 => "110110000101001111000110",
17458 => "110001101011000111111100",
17459 => "101101111110000101000010",
17460 => "101011111011110101111100",
17461 => "101010100111101010111000",
17462 => "101001101101100000110110",
17463 => "101001000111010100110100",
17464 => "101001001010111011011000",
17465 => "101010100010111000011000",
17466 => "101100000101101100110100",
17467 => "101101001000101101001000",
17468 => "101101011011011111011010",
17469 => "101100101011001101111010",
17470 => "101100001101101101000110",
17471 => "101011111001001010010000",
17472 => "101011001001110000100110",
17473 => "101011110001001000101110",
17474 => "101110101100000111101110",
17475 => "110011010011101111110100",
17476 => "111000010110000110000000",
17477 => "111101010110101110011101",
17478 => "000011011011100011110100",
17479 => "001001110101100001101110",
17480 => "001111010010101001010110",
17481 => "010100001001000011100100",
17482 => "010111101100000111011010",
17483 => "011001100011111010111111",
17484 => "011010011110000000011101",
17485 => "011010000010000011110011",
17486 => "011000111011111110111111",
17487 => "011000010001000011000111",
17488 => "010111010001111110010000",
17489 => "010110100001100110101100",
17490 => "010111011011010001101100",
17491 => "011001000001101001101001",
17492 => "011001111111111010100011",
17493 => "011010101111111100001110",
17494 => "011011001101101101011110",
17495 => "011010110000000101000001",
17496 => "011010001101111000100010",
17497 => "011001111101111001100010",
17498 => "011001010110100101001111",
17499 => "011000110100101100001110",
17500 => "011000101010111010100110",
17501 => "011000010110110101110001",
17502 => "010111100110101011000010",
17503 => "010111010100100010101000",
17504 => "010110011110111011101110",
17505 => "010001011000011100011110",
17506 => "001000111110000100110101",
17507 => "111101110010010100001100",
17508 => "101110000100100111011110",
17509 => "100010100100111100111110",
17510 => "100001010110011011001101",
17511 => "100010001000011101001001",
17512 => "100001010100000010010000",
17513 => "100001100001111001000111",
17514 => "100001100111100001100101",
17515 => "100001011000111101111001",
17516 => "100010000110001001011111",
17517 => "100010110010101111000001",
17518 => "100010111011101100111111",
17519 => "100011001011001101010011",
17520 => "100011000101101110011010",
17521 => "100011101110110101000101",
17522 => "101000000010101000001100",
17523 => "101111101001011001100110",
17524 => "110111100011100110100111",
17525 => "111100110100001111110101",
17526 => "111110101000011110011010",
17527 => "111111110101111100101001",
17528 => "000001111100101111011010",
17529 => "000011100100100101101001",
17530 => "000011001100011111011011",
17531 => "111111101001100010010010",
17532 => "111001100100100011101011",
17533 => "110011011010010010101010",
17534 => "101111011101000000100010",
17535 => "101110001111000010111010",
17536 => "101110110011001111110010",
17537 => "110000100110101001100010",
17538 => "110100010001010011000101",
17539 => "111010001000000111111011",
17540 => "000000001110001101110101",
17541 => "000101011100001110000010",
17542 => "001010110011010101101001",
17543 => "010000110100110101000110",
17544 => "011000000010010001011011",
17545 => "011101100101100100110010",
17546 => "011110011001101011100011",
17547 => "011110000110110001010010",
17548 => "011110101010101111110001",
17549 => "011110101010110111110111",
17550 => "011110101100111011100111",
17551 => "011101110100001001111101",
17552 => "011011111111010001100111",
17553 => "011011001101010001110001",
17554 => "011001000100110100010110",
17555 => "010010101011100010010000",
17556 => "001011011110110000001010",
17557 => "000111010011010010011111",
17558 => "000100100011100111101100",
17559 => "000001110100000000101010",
17560 => "111111101111010011000000",
17561 => "111110101001011101010001",
17562 => "111110101101011111001011",
17563 => "111111000110101100011110",
17564 => "111111000111110011001001",
17565 => "111110101001110000000111",
17566 => "111110101001010010101101",
17567 => "000001000101000000011100",
17568 => "000100010111011100100011",
17569 => "000110011101010110011111",
17570 => "001000011000011010110100",
17571 => "001010010000111000101010",
17572 => "001010111100000110000001",
17573 => "001000001100111111100000",
17574 => "000001011010011111010100",
17575 => "111000101110010110000001",
17576 => "101110110110110001100100",
17577 => "100101110010001101111010",
17578 => "100001100111111011000101",
17579 => "100001110000100011010101",
17580 => "100010000100001000010111",
17581 => "100001110101100110000101",
17582 => "100001110110110110010111",
17583 => "100010010100111110110101",
17584 => "100110011011110001000010",
17585 => "101101111000110010101100",
17586 => "110100010101010111000110",
17587 => "111010101001111001110101",
17588 => "000000101010001110001001",
17589 => "000011101100011100111110",
17590 => "000100011001011100100000",
17591 => "000010101010101001010011",
17592 => "111111101000011010001101",
17593 => "111100010100101000101010",
17594 => "111000001001111100110010",
17595 => "110110110101000111101000",
17596 => "111000111010111101101110",
17597 => "111001110101110001011111",
17598 => "111001001110101011101100",
17599 => "111000111010010010100111",
17600 => "111000111010011100100011",
17601 => "111000001001110000010101",
17602 => "110110100111100011111001",
17603 => "110110010110011100011110",
17604 => "110111110101100100100010",
17605 => "111010011000110100000010",
17606 => "111110010000011011011000",
17607 => "000010111110011010000011",
17608 => "000111100000011011101001",
17609 => "001011101100110111101010",
17610 => "001111110011101000100110",
17611 => "010011010000000100100010",
17612 => "010110000101110111000100",
17613 => "011001011100010010000111",
17614 => "011011011011100110101101",
17615 => "011001100100011111100001",
17616 => "010101110101101001011010",
17617 => "010010011010010010100010",
17618 => "001110110001111011000110",
17619 => "001010100010001101011101",
17620 => "000110111010100011110001",
17621 => "000101111101011011100001",
17622 => "000111001000110001010110",
17623 => "001001001010001010110101",
17624 => "001100101111110101010000",
17625 => "010001010100100100101100",
17626 => "010101100111111011011110",
17627 => "011000010111110100000101",
17628 => "011000010110111000011110",
17629 => "010111011001100001011110",
17630 => "010110110011100001110100",
17631 => "010101111010011011101100",
17632 => "010100111000000110110000",
17633 => "010100001010110110011110",
17634 => "010011101001010101111010",
17635 => "010000101010101100011000",
17636 => "001010001001000011100010",
17637 => "000100000001000101110011",
17638 => "000001001101110101111001",
17639 => "000000111100010101101000",
17640 => "000000100101100011000110",
17641 => "111111010010001011010000",
17642 => "111101101100000000001011",
17643 => "111001111100011101011000",
17644 => "110011010100001000101000",
17645 => "101011100111001010000010",
17646 => "100101000101010100111110",
17647 => "100010000100001001011001",
17648 => "100001110100011000001001",
17649 => "100001110100010101111101",
17650 => "100001011000010001111111",
17651 => "100001011101010101010001",
17652 => "100001101111011000101111",
17653 => "100001011011100101010110",
17654 => "100010001000010101000101",
17655 => "100010110010110010000000",
17656 => "100100100010100000111011",
17657 => "101100110101000111010110",
17658 => "110111011110101010101110",
17659 => "111111000011001000111111",
17660 => "000101010111011101100101",
17661 => "001000101101000101000110",
17662 => "000111111100001001000100",
17663 => "000110000100010100101101",
17664 => "000100000001011100010001",
17665 => "000000010010110011010001",
17666 => "111010001011101101100101",
17667 => "110100001001111011101011",
17668 => "101111110010000100000110",
17669 => "101101100100101111001010",
17670 => "101110010010110010001110",
17671 => "101111111000011101110110",
17672 => "110000100100110001100100",
17673 => "110000000110110110000110",
17674 => "101111111011111100000110",
17675 => "110010011110111111011010",
17676 => "110110100000011001101010",
17677 => "111010111010001100110011",
17678 => "000000010010000110011101",
17679 => "000110100110101111110000",
17680 => "001101011000111010010110",
17681 => "010001100000111010101000",
17682 => "010001111110011001111100",
17683 => "010001001110110100101110",
17684 => "001111100001001000001110",
17685 => "001101100011110101111010",
17686 => "001100110110010010100110",
17687 => "001100100011001000011110",
17688 => "001011101101111001010110",
17689 => "001001101000111001011010",
17690 => "000101111010101101000001",
17691 => "000010000101100100001000",
17692 => "111111011001100010111110",
17693 => "111101010100001110111010",
17694 => "111011101100010011111011",
17695 => "111011000000100010011000",
17696 => "111011101010110001101000",
17697 => "111101001110011110111101",
17698 => "111110010100110100111100",
17699 => "111111011000011000000000",
17700 => "000001101001110100110010",
17701 => "000101010111111101000000",
17702 => "001001100011010010110000",
17703 => "001100000101001010100100",
17704 => "001101101000110101101010",
17705 => "001111001111110100101000",
17706 => "001110101011111101011000",
17707 => "001011110100100010010111",
17708 => "001000101001010001101100",
17709 => "000101110010101111101000",
17710 => "000010111000010010100000",
17711 => "000000011001000101001010",
17712 => "111111111010100000011010",
17713 => "000000111011100001001100",
17714 => "000010001010000010010100",
17715 => "000010100100110101101011",
17716 => "000001010110101100101010",
17717 => "111111111011100001111100",
17718 => "111110010100101111000011",
17719 => "111100010011111100001111",
17720 => "111011001111111111110011",
17721 => "111010000000011101100101",
17722 => "111001000100001100000010",
17723 => "111010001011111011000000",
17724 => "111011101100011011001111",
17725 => "111100111011111010011001",
17726 => "111111010010101111011001",
17727 => "000010011010101111001001",
17728 => "000100110100010100001000",
17729 => "000110011000110001110001",
17730 => "000110100100001101110011",
17731 => "000011101001000100101101",
17732 => "111110110001111111001011",
17733 => "111010010101011110110001",
17734 => "110110010110000011100010",
17735 => "110000100110000011100010",
17736 => "101000110000011111001010",
17737 => "100100000010011000110111",
17738 => "100100001111010100000011",
17739 => "100101001001001000010101",
17740 => "100101011000011010110000",
17741 => "100101110011100110111101",
17742 => "100110110110100100010101",
17743 => "100111110101010010111111",
17744 => "101000101110110001111000",
17745 => "101101011011011000010110",
17746 => "110110010101100101111000",
17747 => "111110110110100110101000",
17748 => "000101010111100101101011",
17749 => "001010011111011001011111",
17750 => "001110011001101110111000",
17751 => "010001011000011010010000",
17752 => "010011010101111101010110",
17753 => "010011111110111101000010",
17754 => "010011100001110110100110",
17755 => "010010111101011111010010",
17756 => "010010011111111101111010",
17757 => "010010000000010010100110",
17758 => "010010010110101011010110",
17759 => "010011100000110100100000",
17760 => "010100101000000000010110",
17761 => "010101010010001011000100",
17762 => "010101101010110110111100",
17763 => "010111001001000111101100",
17764 => "011000111010010100110101",
17765 => "011000101001011010001001",
17766 => "010111110100010111000000",
17767 => "011000000100001000001101",
17768 => "011000010100001010001111",
17769 => "010111101100100000111100",
17770 => "010110100001101011010110",
17771 => "010110001000101011101110",
17772 => "010110000100000111000000",
17773 => "010101111010100110101000",
17774 => "010110000011110000110110",
17775 => "010100111101111110101110",
17776 => "010100100111000110000010",
17777 => "010011011011101101101010",
17778 => "001010001010010101011111",
17779 => "111011111100000111100001",
17780 => "101110110000100110000100",
17781 => "100100100010101010011001",
17782 => "100000111101001011010011",
17783 => "100001010100001000111100",
17784 => "100001001010011111000011",
17785 => "100001001011110101010011",
17786 => "100001001100111110011101",
17787 => "100001000110000111100011",
17788 => "100001110110010001001100",
17789 => "100100001000011011100111",
17790 => "100101101001110111011101",
17791 => "100100101101010101001000",
17792 => "100100011110101001011101",
17793 => "100100111000111011011111",
17794 => "100100100001001101010111",
17795 => "100100101011100110000001",
17796 => "100101001111110001000100",
17797 => "100110000100110100101011",
17798 => "100110011000010011011111",
17799 => "100110011000000111101101",
17800 => "100110111001000101111111",
17801 => "100111111110000100001001",
17802 => "101011011001000111001010",
17803 => "101110010100001101001100",
17804 => "101111011110001010110000",
17805 => "110011111010101100010110",
17806 => "111001101010001100001110",
17807 => "111100100110000111000000",
17808 => "111110001011010111111110",
17809 => "000000111111101010110011",
17810 => "000110001101111000001100",
17811 => "001011110011110100110100",
17812 => "010000100110111100011010",
17813 => "010100100001000010110110",
17814 => "010111110011010110011010",
17815 => "011011110001000001000011",
17816 => "011110001110010001101111",
17817 => "011110011011000110001111",
17818 => "011110001110001001010111",
17819 => "011101110011101101010001",
17820 => "011101111110010100000111",
17821 => "011101111010111111101011",
17822 => "011100111101000001101101",
17823 => "011100011001100001011111",
17824 => "011100001101011111101000",
17825 => "011010011000011100011101",
17826 => "010100011010001010000000",
17827 => "001101000100101011101100",
17828 => "000111100101111111011110",
17829 => "000010001100010011010110",
17830 => "111110010110001000111111",
17831 => "111100100010100010101011",
17832 => "111001110100001100111001",
17833 => "110111001010100010011100",
17834 => "110110000010100011010101",
17835 => "110110101110000010000100",
17836 => "111000100110100011010111",
17837 => "111010011011110010000000",
17838 => "111100100010001000100010",
17839 => "111100111011001001001010",
17840 => "111010010001100000001101",
17841 => "110111100010001010010110",
17842 => "110101100000000000011111",
17843 => "110010100011011110010110",
17844 => "101110001100100001101110",
17845 => "101001001101011110101000",
17846 => "100100111011011111110011",
17847 => "100010001010001000110111",
17848 => "100001111010101011011001",
17849 => "100011011001101110101100",
17850 => "100100010001101010011101",
17851 => "100101000010001101000001",
17852 => "100110001010010101010011",
17853 => "100111100000101001011111",
17854 => "101010010111011110010110",
17855 => "101110010100000111111000",
17856 => "110010110111110101000100",
17857 => "110111001110100000101100",
17858 => "111001011111101101000010",
17859 => "111011100110110001010011",
17860 => "111111000000001011000110",
17861 => "000010001100100011011100",
17862 => "000100111100001111011101",
17863 => "000111011100101000001110",
17864 => "001010011011111000001110",
17865 => "001101010111001000010010",
17866 => "001111100001011000001010",
17867 => "010010010011000111111110",
17868 => "010100011011011100000110",
17869 => "010101000001010111100100",
17870 => "010101100010111000001000",
17871 => "010101011001110000000010",
17872 => "010011110100101101001100",
17873 => "010000111000100101000100",
17874 => "001101111000111000100100",
17875 => "001100011111011100111010",
17876 => "001100100101101010000010",
17877 => "001101011111110100101110",
17878 => "001101101111010010000000",
17879 => "001101101101111001100110",
17880 => "001110101101011101100100",
17881 => "001110101110100101010110",
17882 => "001101001000001111000010",
17883 => "001011110001010000111110",
17884 => "001011100000100011110000",
17885 => "001011100001010010000010",
17886 => "001011011101010000010111",
17887 => "001100110111110010101010",
17888 => "001110100110001000011010",
17889 => "001111000001101001001110",
17890 => "010000000101001111100000",
17891 => "010001101101101100000000",
17892 => "010010001000000011011010",
17893 => "010001001000100001011000",
17894 => "001111011011001001100000",
17895 => "001101011100100001000100",
17896 => "001010110001000111111100",
17897 => "000110111010101101101111",
17898 => "000001100010110111100101",
17899 => "111011100011110110011111",
17900 => "110110010101101000110011",
17901 => "110010000011111011101100",
17902 => "101111101001111111010010",
17903 => "101111011101101101111100",
17904 => "110001110001010100101010",
17905 => "110111010011011011000111",
17906 => "111101110101010000011011",
17907 => "000011110100011111001100",
17908 => "001001010100101010111010",
17909 => "001100111000101001100000",
17910 => "001110010011100100110100",
17911 => "001110010101000010010100",
17912 => "001101000101111111110000",
17913 => "001011000001001011001010",
17914 => "001000000111101100001110",
17915 => "000011101111110100101110",
17916 => "111101000100000011110101",
17917 => "110101001110011011101101",
17918 => "101111011000010011000110",
17919 => "101100010011010110110110",
17920 => "101011011101010001100100",
17921 => "101101011011001111010110",
17922 => "110000100000111001001000",
17923 => "110011010100101100011010",
17924 => "110111010100000100001010",
17925 => "111010111110000101000000",
17926 => "111011110110111011000000",
17927 => "111010111000000001011111",
17928 => "111001111010101010110101",
17929 => "111010100011100100100011",
17930 => "111011001111001100110011",
17931 => "111001010110101011111000",
17932 => "110100110111100001101100",
17933 => "101111001010010001010110",
17934 => "101011000000100100000110",
17935 => "101000010101100100111100",
17936 => "100111000000100000001111",
17937 => "101010000101101001111010",
17938 => "101110111010000111110010",
17939 => "110001001111001011100010",
17940 => "110001000100100011010100",
17941 => "101111001101001110101010",
17942 => "101110001010011100101010",
17943 => "101110110111000101011000",
17944 => "110001000000100000010010",
17945 => "110100111100001010001001",
17946 => "111001110001110000111001",
17947 => "111111111011011000010000",
17948 => "000110011010110001000000",
17949 => "001011111101001100101001",
17950 => "010001100111000011111100",
17951 => "010111010011101000001100",
17952 => "011100011000101100010010",
17953 => "011110100101011011110101",
17954 => "011110001101000001110100",
17955 => "011101011111110011110001",
17956 => "011000101000010011111001",
17957 => "010000000001011010110000",
17958 => "001001110101011100100100",
17959 => "000110110010110110110100",
17960 => "000101000010101100011100",
17961 => "000011010000111010101110",
17962 => "000010110100110111100101",
17963 => "000101100011010000111110",
17964 => "001001000101011011011011",
17965 => "001011111110100111100001",
17966 => "001101111111011000000100",
17967 => "001110011011001111100010",
17968 => "001110000110101100110110",
17969 => "001110000111111110100110",
17970 => "001110011100110000100110",
17971 => "001101010010011010011000",
17972 => "001010001011100111010111",
17973 => "000101110110110111100001",
17974 => "000000000010101010010011",
17975 => "111010111011011111100001",
17976 => "111000011010011101000100",
17977 => "110111100100101001111101",
17978 => "110111101001010001100000",
17979 => "110111111001100010011011",
17980 => "111000100110000010011101",
17981 => "111001100011101000111110",
17982 => "111001101111011001011101",
17983 => "111001101111110001101110",
17984 => "111000110111101111001011",
17985 => "110110010001001010110101",
17986 => "110011101010100010011000",
17987 => "110001000111111010111110",
17988 => "101100101100000001011110",
17989 => "100110111111110101010000",
17990 => "100011101000101111010110",
17991 => "100011011111111011000010",
17992 => "100100001101010001010101",
17993 => "100101010000011001101101",
17994 => "100110001111001000100001",
17995 => "100110101101001100001011",
17996 => "101000111110110110011000",
17997 => "101101001000100001111000",
17998 => "110000100111000001100010",
17999 => "110010101000111110000100",
18000 => "110011011000100110100000",
18001 => "110011100111111010011010",
18002 => "110100010000111111000010",
18003 => "110101101100011111101100",
18004 => "110111111001100001111010",
18005 => "111001111101110000111101",
18006 => "111100010001101010010011",
18007 => "111111011100010001000001",
18008 => "000010110011101101000111",
18009 => "000110111110010010001001",
18010 => "001100000111001011110100",
18011 => "010001011000011101101010",
18012 => "010101101101000001111000",
18013 => "010111011101110110100100",
18014 => "010110110100100110001000",
18015 => "010011111011100110011110",
18016 => "001111001100010010010000",
18017 => "001011001001111000010101",
18018 => "001001001000011100011101",
18019 => "001000111101011110010010",
18020 => "001001001111100100111101",
18021 => "001001100101101110100000",
18022 => "001011110000111010111101",
18023 => "001110100110000011101000",
18024 => "010001000000011001110100",
18025 => "010011110001010100111100",
18026 => "010110111000011001011000",
18027 => "011010110100111000011101",
18028 => "011101011000010100001111",
18029 => "011100111111101001010001",
18030 => "011011111100111011000011",
18031 => "011010101110100101010101",
18032 => "011001101101010011010101",
18033 => "011001000111010000011011",
18034 => "010111111111100010011100",
18035 => "010110111011111010001000",
18036 => "010110010011111010110010",
18037 => "010110000100011101101100",
18038 => "010101101000110100100010",
18039 => "010101001011101000100010",
18040 => "010100101111111011100000",
18041 => "010000101011110111000110",
18042 => "001000100111101101100111",
18043 => "000000111000010110010101",
18044 => "111010111111000010101100",
18045 => "110101100000000110110101",
18046 => "110000000010111101110000",
18047 => "101101110111011010011110",
18048 => "101111010011101010001000",
18049 => "101111100011011010010000",
18050 => "101110100110100101011110",
18051 => "110000101111011010011100",
18052 => "110110001010001100101100",
18053 => "111010110001010100010110",
18054 => "111101101111010010010011",
18055 => "000010000111101101011011",
18056 => "000111001110101011101010",
18057 => "001001100011011111101000",
18058 => "000110011100011011100111",
18059 => "111110110000100110001110",
18060 => "110101010101100011100000",
18061 => "101010001010001110101110",
18062 => "100001110110001010010111",
18063 => "100000111111011000101000",
18064 => "100001101110110010010010",
18065 => "100001000111011000111100",
18066 => "100001100100101011110110",
18067 => "100010011001001010011111",
18068 => "100011110010111011011001",
18069 => "100111000001110011111111",
18070 => "101010110110101010100100",
18071 => "101101110011000101000110",
18072 => "110001101110011011011010",
18073 => "110110010101000100110000",
18074 => "110101100100000010100111",
18075 => "101111011110010010111100",
18076 => "101011000101001101010010",
18077 => "101010111011101100110110",
18078 => "101100100001100010010000",
18079 => "101110100010101001101100",
18080 => "110011100100011010100110",
18081 => "111100000110101101000011",
18082 => "000011100011000100001110",
18083 => "000110100111010010010001",
18084 => "000111000010111001101001",
18085 => "001001000111000100111000",
18086 => "001100110000000011000100",
18087 => "001101110001101110011010",
18088 => "001011100110011111010111",
18089 => "001001101010010011011001",
18090 => "001010111101000000011101",
18091 => "001110011011010111111110",
18092 => "010001001001000010110000",
18093 => "010011110110101001011010",
18094 => "011000010111000111110101",
18095 => "011100100100100100111100",
18096 => "011101010110110111111000",
18097 => "011011110101100101010101",
18098 => "011010110101100000001111",
18099 => "011010011001110001110101",
18100 => "011010000011000000001011",
18101 => "011001101001111101010000",
18102 => "011000001111001000100011",
18103 => "010100101000101111100010",
18104 => "001111110111001100000010",
18105 => "001100100110011000110000",
18106 => "001010010111011001111100",
18107 => "000111011101011010110100",
18108 => "000011010100000010110001",
18109 => "111101101011101110010111",
18110 => "111001100100110100101100",
18111 => "111000001000010111110001",
18112 => "110110111100000110000011",
18113 => "110110111100011101001010",
18114 => "111000001100110001101110",
18115 => "110111011110111011111011",
18116 => "110100000000011010001100",
18117 => "101111100011011101101010",
18118 => "101011111010100101001100",
18119 => "101001111100100010010110",
18120 => "101001111000101101101000",
18121 => "101010101110101111111010",
18122 => "101010001110111111001000",
18123 => "101000001011000000001010",
18124 => "100110111101101011100001",
18125 => "100111100000000111000001",
18126 => "101000100100010110000100",
18127 => "101010010110011001001010",
18128 => "101100011110010111110110",
18129 => "101101100000100101110000",
18130 => "101101100111000000101000",
18131 => "101011110101110010000010",
18132 => "101000011111100010101100",
18133 => "100110100111000001100101",
18134 => "100110110010010100110110",
18135 => "100111111010000100001011",
18136 => "101000110000111010011100",
18137 => "101010000001100011111010",
18138 => "101110100101001000100000",
18139 => "110101101000000011110100",
18140 => "111100001010100001100111",
18141 => "000001111010101011000011",
18142 => "000111111111111010100110",
18143 => "001110010010101110000100",
18144 => "010011101000100001101010",
18145 => "010111110100001111000000",
18146 => "011010100011011000101011",
18147 => "011011111111101000010111",
18148 => "011100111001001010100000",
18149 => "011100000001111010100010",
18150 => "011001001000001001010111",
18151 => "010101111100110010100000",
18152 => "010100000100100111110100",
18153 => "010011110011100111000110",
18154 => "010011000111111101000110",
18155 => "010000110101101101100000",
18156 => "001101010100011000111110",
18157 => "001000111010011101000001",
18158 => "000101001111110111010010",
18159 => "000011001011001010100000",
18160 => "000010010010111000110010",
18161 => "000010010000000001110111",
18162 => "000001101000000110101001",
18163 => "111111111101101101100101",
18164 => "111111000110011010001001",
18165 => "000000001001111100010110",
18166 => "000010001101011000001000",
18167 => "000100010000111101111000",
18168 => "000110000010001010000001",
18169 => "000111010110101110000101",
18170 => "000111101101011010010100",
18171 => "000110011111000010101110",
18172 => "000100110000011000110100",
18173 => "000011110000001101101001",
18174 => "000010110101101100011011",
18175 => "000001011100110111110000",
18176 => "111111011010011111011100",
18177 => "111100001110110011011111",
18178 => "110111010000110101100010",
18179 => "110001001011101100011010",
18180 => "101100010011111010001110",
18181 => "101001010111000010011100",
18182 => "100111101001110001000101",
18183 => "100110011001001101101111",
18184 => "100100111110010011100111",
18185 => "100100111111100101000010",
18186 => "101000001101111111010010",
18187 => "101101111000001111111010",
18188 => "110100010110011001101100",
18189 => "111100011000000001011000",
18190 => "000110101110011000101110",
18191 => "001111110001000000110000",
18192 => "010101100000100110010110",
18193 => "011001111100001111101001",
18194 => "011100101110011101111010",
18195 => "011100101110110100111101",
18196 => "011011010011110110100101",
18197 => "011010100001011011101001",
18198 => "011010010110000001110101",
18199 => "011001100111010100101101",
18200 => "010111110110111001111100",
18201 => "010011111111001010011100",
18202 => "001110110000000100111110",
18203 => "001001011110000100111100",
18204 => "000011010101011011010000",
18205 => "111101111110111000110111",
18206 => "111011110100100000101001",
18207 => "111100100101010000000100",
18208 => "111110001111010101010110",
18209 => "111110110000000111010001",
18210 => "111111011111111111011100",
18211 => "000010001011100010001010",
18212 => "000101011110110010001101",
18213 => "000111111011000101110110",
18214 => "001001111110011000001000",
18215 => "001011111100010000001111",
18216 => "001001110000110111110111",
18217 => "000001100101101000101001",
18218 => "111001000110111101110000",
18219 => "110011101100011101100100",
18220 => "101110100110110110000100",
18221 => "101000010001010010000100",
18222 => "100011101010110110001001",
18223 => "100010100000011101000101",
18224 => "100010101111111011000101",
18225 => "100011101011110010101011",
18226 => "100100010100000101111101",
18227 => "100101000001011011000001",
18228 => "101001100100010111010000",
18229 => "110000111011111111101100",
18230 => "111000001001010010101111",
18231 => "111111100111111111001101",
18232 => "000111011100001111000101",
18233 => "001111001010011101101100",
18234 => "010101110101111111101110",
18235 => "011010010111111000101100",
18236 => "011100011100011011110101",
18237 => "011100000001010100011101",
18238 => "011010101001101011111101",
18239 => "011001100101011101111011",
18240 => "011000101000010000010111",
18241 => "010110110110010111111100",
18242 => "010010111000101011100110",
18243 => "001110101011000011111010",
18244 => "001011110010001001011010",
18245 => "000111001110010101000100",
18246 => "000001011010100011101010",
18247 => "111110111101101000001101",
18248 => "000000010010010110110010",
18249 => "000000011100111111011110",
18250 => "111100100000010000101110",
18251 => "111001101011000010110000",
18252 => "111011110010001000010010",
18253 => "111101100000111001100001",
18254 => "111100100101010101100110",
18255 => "111100111100110111110111",
18256 => "111111010100000010000111",
18257 => "000000101101100011011100",
18258 => "111111010011010011000011",
18259 => "111101001010110011011100",
18260 => "111100100010111010101100",
18261 => "111100010000100110010100",
18262 => "111011011101000001100101",
18263 => "111010010011101010000010",
18264 => "111000110001101111011000",
18265 => "110101111000100001010000",
18266 => "110000111100000100111100",
18267 => "101101000001100010001010",
18268 => "101100010000111111100110",
18269 => "101100000010100110001100",
18270 => "101010001011111010010110",
18271 => "101000011100001010111110",
18272 => "101001010110001100100010",
18273 => "101011000110001110011010",
18274 => "101010101010111101010100",
18275 => "101001010010100110100000",
18276 => "101001111011000011001010",
18277 => "101101011011000010110110",
18278 => "110001100111111000010110",
18279 => "110101000101111111001010",
18280 => "111001001010101000101110",
18281 => "111110011110001110001001",
18282 => "000011110011000010001110",
18283 => "000111010011111110001110",
18284 => "001000111100001011111001",
18285 => "001010011000000110111100",
18286 => "001100100101101111010110",
18287 => "001111010110100001010110",
18288 => "010001110001101010111010",
18289 => "010100000100101111110000",
18290 => "010101110001000000011000",
18291 => "010101001111110000000000",
18292 => "010011101001100100100110",
18293 => "010010011100100111100010",
18294 => "010001111000100110010000",
18295 => "010001001100011111101110",
18296 => "001111000001111001011110",
18297 => "001100100001000110010000",
18298 => "001010001111010111001010",
18299 => "001000001101011100010110",
18300 => "000111110011101111010001",
18301 => "001000100111101001010111",
18302 => "001010011011001111000000",
18303 => "001101110101110000011110",
18304 => "010001110111100111000000",
18305 => "010100001001010100100000",
18306 => "010011010110010111011010",
18307 => "010000111101111001110100",
18308 => "001101110101100000110100",
18309 => "001001110101111110010010",
18310 => "000100011110101101101100",
18311 => "111101000010011001101100",
18312 => "110100011110111010010110",
18313 => "101010101000111001111000",
18314 => "100010110000110000000111",
18315 => "100001010101100011010000",
18316 => "100001111011111000010111",
18317 => "100001011111101101010111",
18318 => "100001101000000100011101",
18319 => "100001101100101110110110",
18320 => "100010001011100111000101",
18321 => "100010110111000101111001",
18322 => "100011011011010110101100",
18323 => "100100011011100110110001",
18324 => "100100110000110110110011",
18325 => "100110100010000110011010",
18326 => "101100000010111000100110",
18327 => "110010100110010010100000",
18328 => "110110110111111011000111",
18329 => "111000010100010010100100",
18330 => "111001100110001100000000",
18331 => "111100010110010000011101",
18332 => "111110110100001111101111",
18333 => "000000101010011110011100",
18334 => "000010111011010111001101",
18335 => "000100100000111001000110",
18336 => "000100010101110101000100",
18337 => "000011100010101110000110",
18338 => "000011000011010101010110",
18339 => "000010101000101001100000",
18340 => "000010101111110001010100",
18341 => "000100010000001001110010",
18342 => "000110010011011110101010",
18343 => "000111010111001010000000",
18344 => "000111101001011111111110",
18345 => "001001001010100001010000",
18346 => "001101101010010110110000",
18347 => "010010001101000111100010",
18348 => "010100011010010100001010",
18349 => "011000101110100000111011",
18350 => "011101111010100011101001",
18351 => "011110101101101001101001",
18352 => "011110001111100001000010",
18353 => "011110010011001101111001",
18354 => "011101001111110101011001",
18355 => "011011001111100001100001",
18356 => "010111001011111010010100",
18357 => "010001001100001101001010",
18358 => "001001011111110000100001",
18359 => "111111110010101101100110",
18360 => "110110000011100100110101",
18361 => "101111010011110011000010",
18362 => "101110001001011011111010",
18363 => "110000110110000111100000",
18364 => "110100010110000110111011",
18365 => "111000001000101110011000",
18366 => "111011001100001001000111",
18367 => "111101100100101110101010",
18368 => "111111010100100100101110",
18369 => "000000011100000111010001",
18370 => "000010110001100101010010",
18371 => "000101101011101000011000",
18372 => "000111111011001100111100",
18373 => "001010101010000110011101",
18374 => "001110110101111101000010",
18375 => "010010001101011000110000",
18376 => "010001100100110100011110",
18377 => "001111011100010100010000",
18378 => "001110111010110000101000",
18379 => "001110001011011011101010",
18380 => "001010100101010011001000",
18381 => "000011000010001100001010",
18382 => "111000110001111101000111",
18383 => "101101011101011101110100",
18384 => "100100011001101110101100",
18385 => "100001011100101110100101",
18386 => "100001101001010110010001",
18387 => "100001011111010100000111",
18388 => "100001100101110001101011",
18389 => "100010111100110010101011",
18390 => "100111110100101101000101",
18391 => "101110110010111100110010",
18392 => "110011101000001110011110",
18393 => "110110101101101011110000",
18394 => "111001110001001111000100",
18395 => "111101111101001111100000",
18396 => "000011100101011000010000",
18397 => "000111101100001101011100",
18398 => "001001000111100101010010",
18399 => "001001010110000111101010",
18400 => "000110110111010011100100",
18401 => "000000111010010001100000",
18402 => "111011100011111101101110",
18403 => "111001110110111101010001",
18404 => "111001110011110100100101",
18405 => "111000011011000100100100",
18406 => "110110101110001111000111",
18407 => "110110101101010011010110",
18408 => "110110101110110011110010",
18409 => "110101101010111001110010",
18410 => "110100110000111011000100",
18411 => "110101001111011001110000",
18412 => "111000000100000011010111",
18413 => "111100010111001111001100",
18414 => "000000101100011110101010",
18415 => "000100111101111110111000",
18416 => "001001001001101110010000",
18417 => "001100010101000110101110",
18418 => "001101011100001110110110",
18419 => "001110101000111010000100",
18420 => "010010011010011011010110",
18421 => "010110100010101011000100",
18422 => "011000111100110000010101",
18423 => "011010010110100101100111",
18424 => "011010101001100010011001",
18425 => "011000010110110110010100",
18426 => "010011110100101101111010",
18427 => "010000000111101000111000",
18428 => "001110100111100101111110",
18429 => "001110001011100011110000",
18430 => "001101111111011011000010",
18431 => "001110001100101101000110",
18432 => "001111110000111110111110",
18433 => "010010110101000110011110",
18434 => "010110000011100101101000",
18435 => "010111111001111000000100",
18436 => "011000000111001101010110",
18437 => "010111110000101101001110",
18438 => "010111011101011110000000",
18439 => "010110111011110110010010",
18440 => "010011101101011000011010",
18441 => "001011111010010010110111",
18442 => "000011000010111011101100",
18443 => "111011110111010001100110",
18444 => "110101101100001010100010",
18445 => "110001011010100111110100",
18446 => "101111001000110110110010",
18447 => "101100011010100111100100",
18448 => "101000110101011000100000",
18449 => "100110011010111011011100",
18450 => "100100101101001011001101",
18451 => "100010100001101101011101",
18452 => "100001101010111110110001",
18453 => "100001101111111010000111",
18454 => "100001010010001110001101",
18455 => "100001010100000011001101",
18456 => "100001101011111110111001",
18457 => "100010011110000001110111",
18458 => "100011011100010111000101",
18459 => "100011111011111011001110",
18460 => "100111100111110110010000",
18461 => "101111011011011001110100",
18462 => "110110011010100100101001",
18463 => "111011000110000100010101",
18464 => "111111011001100001010101",
18465 => "000100000000000100011110",
18466 => "000111001010110111000001",
18467 => "000110100110001010011000",
18468 => "000011001100000101111000",
18469 => "111111001100110011001001",
18470 => "111100000110110000001000",
18471 => "111010010000101001001100",
18472 => "110111110101011010011111",
18473 => "110100110101101001111000",
18474 => "110011110011001111110100",
18475 => "110101101111100111011110",
18476 => "111001110110001000010100",
18477 => "111101110001101110001110",
18478 => "000000101001011100100000",
18479 => "000100011011101000001111",
18480 => "001001101011110001010000",
18481 => "001110100000100001011000",
18482 => "010001001010011110000100",
18483 => "010010101111100010110000",
18484 => "010100111010001101000100",
18485 => "010101110010101001111010",
18486 => "010100010000110110001100",
18487 => "010010100001110011101010",
18488 => "010001100111000000000010",
18489 => "001111100101000000110010",
18490 => "001011001011000110101010",
18491 => "000111000111101100000010",
18492 => "000101100001110111111000",
18493 => "000100110011101110011011",
18494 => "000011110001001010001101",
18495 => "000010001011011010010110",
18496 => "000000001101010110110100",
18497 => "111110100111111000101100",
18498 => "111101010001101010100001",
18499 => "111011010010011000110100",
18500 => "110111100101001110111100",
18501 => "110001110111110010110100",
18502 => "101011101001011000001100",
18503 => "100110101111010010001111",
18504 => "100100001000110001001101",
18505 => "100101001010100010110100",
18506 => "101010100011010111110110",
18507 => "110001111001010111101000",
18508 => "111001000110010010100111",
18509 => "111111101111011001111010",
18510 => "000011111100100110000100",
18511 => "000101100101111001101111",
18512 => "000111001000000011010010",
18513 => "001000111011110100100110",
18514 => "001000110000010101010110",
18515 => "000101101111001000000010",
18516 => "000011110011111010111010",
18517 => "000101100000100011011100",
18518 => "000111100100010110110110",
18519 => "001000000010100101100000",
18520 => "001000101001101110110100",
18521 => "001010110100111100000101",
18522 => "001101110010000111010000",
18523 => "001111001111100101101100",
18524 => "001101111010010101000000",
18525 => "001010001111100111001010",
18526 => "000110001101001011001000",
18527 => "000011100001010000011000",
18528 => "000001110111100000100101",
18529 => "000001000011001000101111",
18530 => "000001000110010011010001",
18531 => "000001000000110011111110",
18532 => "000001011011011011110001",
18533 => "000011010111010010101011",
18534 => "000100101100001101011110",
18535 => "000100001011101110011011",
18536 => "000010111101000111111001",
18537 => "000001001101010101001110",
18538 => "111111110110111000101001",
18539 => "111111011100011010001110",
18540 => "111110110111111011000011",
18541 => "111101100010100101000101",
18542 => "111001110010101101101000",
18543 => "110010101011110111000000",
18544 => "101010100100001000010010",
18545 => "100101001010010100100101",
18546 => "100100001111000010001001",
18547 => "100101111010000100101111",
18548 => "101001011011111111011010",
18549 => "101110001101111000000000",
18550 => "110010001001011110101010",
18551 => "110110111010000110001110",
18552 => "111011111011011101011110",
18553 => "111110001011111000010010",
18554 => "000000100100101001001110",
18555 => "000101000110100011100101",
18556 => "001001001000000111111011",
18557 => "001011000110001000110001",
18558 => "001011100001011100001100",
18559 => "001010100000100100100100",
18560 => "000111011011011100100100",
18561 => "000100000100101010100000",
18562 => "000011000000110111010011",
18563 => "000011111111011010101011",
18564 => "000101100101010010010010",
18565 => "001000000101011001111100",
18566 => "001100100111010000101010",
18567 => "010000111101101001001000",
18568 => "010011000001111011011010",
18569 => "010100101100010010110000",
18570 => "010110110011101001000100",
18571 => "011000000010000011011111",
18572 => "010111111010011111001100",
18573 => "011000000000011110011011",
18574 => "011000110000110010101001",
18575 => "011000101100011111010001",
18576 => "011000010111011111010001",
18577 => "011000000000010111110010",
18578 => "010111100001100011001000",
18579 => "010111011010100111100010",
18580 => "010101111101111111111100",
18581 => "010010110000110001001110",
18582 => "001100011011010110101100",
18583 => "000001010101010100001110",
18584 => "110100111100110111110010",
18585 => "101001100100110001100110",
18586 => "100010000000110011010100",
18587 => "100001000001110000011101",
18588 => "100001101010111001011011",
18589 => "100001100101101110001001",
18590 => "100010110111110101110101",
18591 => "100011101101010100011101",
18592 => "100101001010101010011111",
18593 => "101010011100101000110110",
18594 => "110001001000100000100100",
18595 => "110110011101101110110110",
18596 => "111001111111101011100110",
18597 => "111010101100110111011110",
18598 => "111001011110010110011011",
18599 => "110111101001011111001001",
18600 => "110100100100101000000100",
18601 => "110001000000111011000100",
18602 => "101110001100011010100000",
18603 => "101100000000011000101100",
18604 => "101010001101110001001010",
18605 => "101000110011110001010010",
18606 => "101000100100010011110000",
18607 => "101001100110101111110000",
18608 => "101011101010011100111010",
18609 => "101110111000111100001000",
18610 => "110010011110011111010100",
18611 => "110110001000111110001001",
18612 => "111001100111110011100101",
18613 => "111100010001001011111100",
18614 => "111110111011110010110100",
18615 => "000010011100001101100000",
18616 => "000110011011101010100001",
18617 => "001010010010010001110011",
18618 => "001110010101001100001100",
18619 => "010010110101111010011010",
18620 => "010111001010000000110100",
18621 => "011011010011011101011011",
18622 => "011110000111001111001010",
18623 => "011110100011010110110001",
18624 => "011110010101010110110100",
18625 => "011101110001001110001000",
18626 => "011100100111101000000001",
18627 => "011011111101110011000100",
18628 => "011011100010111011000101",
18629 => "011010111101000100110111",
18630 => "011001101110101000100111",
18631 => "010110001001011111000110",
18632 => "010000011010000001000010",
18633 => "001010110001001111110101",
18634 => "000101101111000001000100",
18635 => "000001010111011100001110",
18636 => "111110110110011011011100",
18637 => "111101111100010011000100",
18638 => "111101011101101000010111",
18639 => "111100100100011100101010",
18640 => "111100000000110001101110",
18641 => "111100011011101111000001",
18642 => "111011010000111111101000",
18643 => "110111110011011100111110",
18644 => "110001101001101010100100",
18645 => "101000000101010000000010",
18646 => "100001100110110100011001",
18647 => "100000111110000101001011",
18648 => "100001001100100111000111",
18649 => "100001110001110100000011",
18650 => "100010110010011110111110",
18651 => "100011110001101110111001",
18652 => "100101110110110100111010",
18653 => "100111000010011011100000",
18654 => "100111011110101010001111",
18655 => "101010000100111101011000",
18656 => "101110010001010111101100",
18657 => "110010000000001100110000",
18658 => "110100101101000100111010",
18659 => "110111001100101001000000",
18660 => "111010001000001011011000",
18661 => "111101011100001011100001",
18662 => "000000001110100101111110",
18663 => "000001101111111111010000",
18664 => "000011110001111100000011",
18665 => "000111001010000001001000",
18666 => "001010010111000011001100",
18667 => "001100100100011010111010",
18668 => "001101010101110010101100",
18669 => "001101100111011011001110",
18670 => "001110110111101111011110",
18671 => "010000101011101001011100",
18672 => "010010001010001101001000",
18673 => "010010001101011110010000",
18674 => "010001011111101100100000",
18675 => "010010010101001010000110",
18676 => "010011100000000101100100",
18677 => "010010100100000110001000",
18678 => "010000010000001010111110",
18679 => "001110010000000111010110",
18680 => "001100110011101000010110",
18681 => "001011101000111111100110",
18682 => "001100001110100110110010",
18683 => "001111001111000101010110",
18684 => "010010101010011100111000",
18685 => "010101011110110010000010",
18686 => "010110101010011011000100",
18687 => "010101010111100111001110",
18688 => "010011011101010011111000",
18689 => "010010011110001010000010",
18690 => "010010111000001100111100",
18691 => "010011101101000111011010",
18692 => "010011010101110111001000",
18693 => "010010010001100111001010",
18694 => "001111101111111100000000",
18695 => "001011110100101001111001",
18696 => "001001001111101100111110",
18697 => "000111010000000101011011",
18698 => "000100010001010100010001",
18699 => "000001001100001101000110",
18700 => "111110010101110010011100",
18701 => "111010111110110001001011",
18702 => "110101100110000011111111",
18703 => "101110101111100010100010",
18704 => "101000111110011001010100",
18705 => "100101101100111000011001",
18706 => "100101100100110101111100",
18707 => "100111110101000110101101",
18708 => "101100000111011100001000",
18709 => "110010110000001101001100",
18710 => "111001001000101110011001",
18711 => "111101011001100111100100",
18712 => "000000011110001010111001",
18713 => "000010111001010000010010",
18714 => "000100001010001000111100",
18715 => "000011000011000000111011",
18716 => "000000010001110000111011",
18717 => "111101101111001001011011",
18718 => "111010111000010000111000",
18719 => "110110111110110011100110",
18720 => "110010000001000010101100",
18721 => "101100001110111111100110",
18722 => "100111100100101111100011",
18723 => "100101011011101001001101",
18724 => "100101101101001011100111",
18725 => "100111101001101100111111",
18726 => "101001101010000101000100",
18727 => "101011001001010001011100",
18728 => "101101001000110011001100",
18729 => "110000100001000111011100",
18730 => "110100110010111111010010",
18731 => "111000100111110010101011",
18732 => "111011001011100110100101",
18733 => "111011111111111011011000",
18734 => "111100010100000010110111",
18735 => "111110001000111001111100",
18736 => "000000100111110010110001",
18737 => "000010011111100100111110",
18738 => "000010111101001011000111",
18739 => "000001010100111011111001",
18740 => "111111010111101111000010",
18741 => "111110000001101010110101",
18742 => "111100110110111000101011",
18743 => "111100000111011000111100",
18744 => "111011001111100010111011",
18745 => "111010010001110011011111",
18746 => "111001010010001001100010",
18747 => "110111110111011010011010",
18748 => "110110110100110100001100",
18749 => "110110110101010110100000",
18750 => "111000111011010100100000",
18751 => "111101011000011110100001",
18752 => "000010111101110101010100",
18753 => "001000111110001100000000",
18754 => "001110011010111011001010",
18755 => "010011011100010110100100",
18756 => "011000001011011000011011",
18757 => "011010110101100101000110",
18758 => "011011101101110110100001",
18759 => "011011101111100111101000",
18760 => "011010000000111011011101",
18761 => "010110001010011100111000",
18762 => "010001000110011110000110",
18763 => "001100101010110100111110",
18764 => "001001010100101011101010",
18765 => "000110001011101011100001",
18766 => "000011110001111011111011",
18767 => "000011001011111010001001",
18768 => "000101001001011011100100",
18769 => "001001010110111001010110",
18770 => "001101100100101010001100",
18771 => "001111111100101011011110",
18772 => "010000100100001100100000",
18773 => "010000000100111000110100",
18774 => "001110110101001010011010",
18775 => "001100011110111110001010",
18776 => "001000001101000011001111",
18777 => "000010111111001110011000",
18778 => "111110110110111111001101",
18779 => "111011110101110001100000",
18780 => "111000101111101001101010",
18781 => "110100101011110011111100",
18782 => "110000111000110000001000",
18783 => "101110111011010011110100",
18784 => "101101011110000110101100",
18785 => "101100011011010000010100",
18786 => "101011100110111101100010",
18787 => "101000001001010001000000",
18788 => "100100000011101010100110",
18789 => "100011010000101111000001",
18790 => "100011111000010110100001",
18791 => "100100001010100010100111",
18792 => "100101001111111110011101",
18793 => "100110100000010100000101",
18794 => "100110110011010110001101",
18795 => "100111001001101110000111",
18796 => "100111110011111011011011",
18797 => "100111111100001001000011",
18798 => "101001000011001000111100",
18799 => "101100100110000000100110",
18800 => "110000101110000110110110",
18801 => "110100010101001011111010",
18802 => "111000101001101100101100",
18803 => "111100110011010010110111",
18804 => "111111001000011001000101",
18805 => "000000100111011110001001",
18806 => "000010000000100111110001",
18807 => "000011001100110010110000",
18808 => "000100011011101000000000",
18809 => "000101001000001110010101",
18810 => "000100011010111000101101",
18811 => "000010011001110011000110",
18812 => "000001001110100110111001",
18813 => "000010101101111001101100",
18814 => "000101010001111101100100",
18815 => "000111011001011111011010",
18816 => "001001111000110111011110",
18817 => "001101111111111011111000",
18818 => "010011010011010011111000",
18819 => "010111101011100111000010",
18820 => "011001111010110001011011",
18821 => "011001010011101001100111",
18822 => "010110101111110110100110",
18823 => "010101010101111110101100",
18824 => "010101000111110010011100",
18825 => "010100100100111001001110",
18826 => "010100101101010001100000",
18827 => "010110001011101011011100",
18828 => "010111101100000000100110",
18829 => "010111100010011111110110",
18830 => "010110011010010100010110",
18831 => "010110011110010111101000",
18832 => "010111100111011110110100",
18833 => "011000010111011010101001",
18834 => "011000001011000011111101",
18835 => "010110111000100010101100",
18836 => "010011111010100101101100",
18837 => "001111101100101111010000",
18838 => "001100011001001001101000",
18839 => "001010111001000011111100",
18840 => "001010001000100100101011",
18841 => "001001010110010001111101",
18842 => "001000011001101000001111",
18843 => "000110111100010100001100",
18844 => "000100100000100010010110",
18845 => "000001011001101011111011",
18846 => "111110011101110111001100",
18847 => "111100110000011000011101",
18848 => "111100000010110101000100",
18849 => "111010100001100010011101",
18850 => "111000111000110110011100",
18851 => "111000111001001010000110",
18852 => "111001011001000111100100",
18853 => "111000100101010001000000",
18854 => "110101100010011000000010",
18855 => "110001010100010100101100",
18856 => "101110100000001001011100",
18857 => "101101110111100001001110",
18858 => "101111000110100101110010",
18859 => "110001011001001110001010",
18860 => "110011111110011111010110",
18861 => "110111100100010100011110",
18862 => "111010101100110000000110",
18863 => "111010011111010011111011",
18864 => "111000000111100011111010",
18865 => "110101100111001110100110",
18866 => "110010010000101110101110",
18867 => "101110010011100001011100",
18868 => "101011001111011001010000",
18869 => "101000111110011100010100",
18870 => "100111000000010111010001",
18871 => "100110001010001010101111",
18872 => "100111110110100010000011",
18873 => "101100001101010100100110",
18874 => "110001100111011001010000",
18875 => "110110010111111011011010",
18876 => "111001101110011001000111",
18877 => "111100010000100111110111",
18878 => "111110110011110110101110",
18879 => "000000100110011011000000",
18880 => "000000100001110111111101",
18881 => "111110111001000110001101",
18882 => "111101011000111100101110",
18883 => "111101011000000110100000",
18884 => "111101111101000100010010",
18885 => "111110100100110000100001",
18886 => "000000110101010000001111",
18887 => "000101000111111011010100",
18888 => "001001010111101000011101",
18889 => "001011110011101000000100",
18890 => "001101000111100001111110",
18891 => "001110110011111011011100",
18892 => "010000000001110000101100",
18893 => "001110101111110000111100",
18894 => "001011111001010010000100",
18895 => "001010010000101001011100",
18896 => "001010100000101010100100",
18897 => "001011100001010111111010",
18898 => "001100001010010111001000",
18899 => "001100011001000111000010",
18900 => "001101011110010111101010",
18901 => "001111111010101010011010",
18902 => "010011100000111110110100",
18903 => "010111100001111111000100",
18904 => "011001101000010001110111",
18905 => "011001011000110101110001",
18906 => "011000110111100101001001",
18907 => "011000000100110100000011",
18908 => "010110000011000101110110",
18909 => "010011001111101101101110",
18910 => "010000001110000000110110",
18911 => "001110001100101111000100",
18912 => "001110011111101001110000",
18913 => "001111001000101000011000",
18914 => "001101000001001100010000",
18915 => "001000100111100110110110",
18916 => "000100010110011110011001",
18917 => "000001000001010100101011",
18918 => "111101111011101011010000",
18919 => "111010101101001011000110",
18920 => "110111110100010000000110",
18921 => "110101001011001101001110",
18922 => "110010010000000111001010",
18923 => "101111000001101001110000",
18924 => "101011010010000100011010",
18925 => "100111100000101010011000",
18926 => "100100110100011001000101",
18927 => "100011000011100101000111",
18928 => "100010000000101011000001",
18929 => "100001110000100010011100",
18930 => "100001111010001011011110",
18931 => "100010100010000101110001",
18932 => "100011010010010110110101",
18933 => "100011101010001111101000",
18934 => "100100010001001101011011",
18935 => "100101001111010111110011",
18936 => "100110001011010101010111",
18937 => "100110111011000010010011",
18938 => "100111001001000010101110",
18939 => "100111000100010001111001",
18940 => "100110111101101010101111",
18941 => "100111001000010010100101",
18942 => "101001001000101000101000",
18943 => "101101101010100100011100",
18944 => "110011100010011000101100",
18945 => "111001111110000001111011",
18946 => "000000111000010110001110",
18947 => "001000000110010101000111",
18948 => "001110110011011001110010",
18949 => "010100000011101001100110",
18950 => "011000100000111111011110",
18951 => "011100011000001101010101",
18952 => "011110001010101011111000",
18953 => "011110100111000100011111",
18954 => "011110101101101100011110",
18955 => "011011111011111110101101",
18956 => "010101111110011101110000",
18957 => "010000011101111100100110",
18958 => "001100100111001111101010",
18959 => "001001110101111111011111",
18960 => "001000110001110110011000",
18961 => "001001011001101011011000",
18962 => "001010110110100011101010",
18963 => "001011111011111100011010",
18964 => "001011011000010111101110",
18965 => "001001101000000101110010",
18966 => "001000000011010110101000",
18967 => "000111001010011100110111",
18968 => "000111010001011001100010",
18969 => "001000101100111011111001",
18970 => "001011001010100110010110",
18971 => "001101110000001000000110",
18972 => "001110111010001110000100",
18973 => "001101100101100011010000",
18974 => "001010110101010000101101",
18975 => "001000110001101110101010",
18976 => "000111111000100110100001",
18977 => "000110100001111001001100",
18978 => "000011101110110001111010",
18979 => "000000010011100011011011",
18980 => "111100110101000001011000",
18981 => "111000111000011100101110",
18982 => "110100000100010000100111",
18983 => "101110101101101110000100",
18984 => "101001110010110001111000",
18985 => "100101011101010010111011",
18986 => "100001111001010011100101",
18987 => "100000101110110110111010",
18988 => "100001011011011001010111",
18989 => "100001100010101100010111",
18990 => "100001100111110010001111",
18991 => "100010011111111110100101",
18992 => "100011011111111111101111",
18993 => "100110110010110000101111",
18994 => "101110011011110001011110",
18995 => "111000000011100111000100",
18996 => "000000101011001100110010",
18997 => "000111000011100110011001",
18998 => "001011010001111001010001",
18999 => "001110011010111111111100",
19000 => "010000001101001001101110",
19001 => "001111100011000100010100",
19002 => "001101011001000000110000",
19003 => "001011001111011110110101",
19004 => "001001010110011101101000",
19005 => "000111101001111001101011",
19006 => "000110000111111111001011",
19007 => "000100100110111011111010",
19008 => "000011010001010111000110",
19009 => "000010011010100011101110",
19010 => "000001110011010111001100",
19011 => "000000110110000100101001",
19012 => "111111010001000000001000",
19013 => "111101011001001100011010",
19014 => "111011110011000101111110",
19015 => "111010110000001100001011",
19016 => "111010111011011011101111",
19017 => "111101110100101010101110",
19018 => "000011011011010101001100",
19019 => "001000101110001000100000",
19020 => "001011011001100101111000",
19021 => "001101001110001001111100",
19022 => "001111011010111001001100",
19023 => "001110100111101110010110",
19024 => "001000110100110011111001",
19025 => "000001011111101011010110",
19026 => "111011001101110110110101",
19027 => "110100101100111011000010",
19028 => "101110010101001000000110",
19029 => "101011000100001011000000",
19030 => "101010111010010101110010",
19031 => "101011001100110011111000",
19032 => "101100001000010010000010",
19033 => "101111111000011110010010",
19034 => "110101100110110011100010",
19035 => "111010110111101111010101",
19036 => "111111100111101110111100",
19037 => "000100100001101111101000",
19038 => "001001001000001001101101",
19039 => "001101010011100111010010",
19040 => "010001000010110001101010",
19041 => "010011001101001001111110",
19042 => "010010101011101000100000",
19043 => "010000011010100010011100",
19044 => "001111000111000010011000",
19045 => "001111101001000111110110",
19046 => "010000010001111110101010",
19047 => "010000011000101011110000",
19048 => "010000011011010110010000",
19049 => "001111100001000101000000",
19050 => "001101011010011110101100",
19051 => "001011011011001010100000",
19052 => "001001000101110110000100",
19053 => "000101101010111011100011",
19054 => "000011011110000110011100",
19055 => "000100000010001000010010",
19056 => "000101100110100100111110",
19057 => "000110011000101000000111",
19058 => "000110000011010110000100",
19059 => "000101011100101110111000",
19060 => "000101010110011100000001",
19061 => "000100111001111110111110",
19062 => "000011100000101000011101",
19063 => "000010100111110011111010",
19064 => "000011010100011001111111",
19065 => "000011100010000000000000",
19066 => "000000111110001111100001",
19067 => "111101000010001010111110",
19068 => "111001000111000011101011",
19069 => "110100000101101101000010",
19070 => "101110101111111111111100",
19071 => "101011000101111100110100",
19072 => "101000001101100110101110",
19073 => "100101010101100111100000",
19074 => "100100001000000101100011",
19075 => "100100101010110100100100",
19076 => "100101011001001000101010",
19077 => "100101101110110011101001",
19078 => "100101100100110000011111",
19079 => "100110110101110110000001",
19080 => "101100010101000111001110",
19081 => "110011101110111100111010",
19082 => "111000011111010010010101",
19083 => "111010011101000101010100",
19084 => "111100001101001101100011",
19085 => "111111001010010000010110",
19086 => "000010011101001001011010",
19087 => "000100100111101010001110",
19088 => "000111001111001101011000",
19089 => "001100111111001011111010",
19090 => "010011010011011111110100",
19091 => "010110000011000000011100",
19092 => "010111100100011000001100",
19093 => "011010100110100001111001",
19094 => "011011111001110011010111",
19095 => "011010011100100101111111",
19096 => "011001010111011001000110",
19097 => "011000000111110111011111",
19098 => "010100011010011001110110",
19099 => "001111010111101011101000",
19100 => "001010101101001011001111",
19101 => "000111011110101101101111",
19102 => "000111000101011101011110",
19103 => "001000000011011000110010",
19104 => "001000101101101100001101",
19105 => "001011011110111110100100",
19106 => "010000010100100100100010",
19107 => "010011011110010000010010",
19108 => "010100011110000110011100",
19109 => "010100110110110110110010",
19110 => "010100110111000011111000",
19111 => "010011110110111110100110",
19112 => "010001100011111000011110",
19113 => "001111101101101010101100",
19114 => "001111000100100010110110",
19115 => "001100101010011100011110",
19116 => "000110011011101110000010",
19117 => "111110001111011101000111",
19118 => "110110110110000111110100",
19119 => "110000011011101101100010",
19120 => "101001100111001110001100",
19121 => "100011100001111101001001",
19122 => "100000110011001111011011",
19123 => "100000110011010001110101",
19124 => "100001001001101011001011",
19125 => "100001010111110010000100",
19126 => "100001101101001000101011",
19127 => "100001110101010110000100",
19128 => "100001100111110110001101",
19129 => "100001100010100011011101",
19130 => "100010001001110111110010",
19131 => "100010111000110011111001",
19132 => "100011011010001011111001",
19133 => "100101011100100101110100",
19134 => "101010001101101110010100",
19135 => "110000100100001001011110",
19136 => "110110011100110111011100",
19137 => "111010110010100011001000",
19138 => "111110010001111010001110",
19139 => "000001101000110000110010",
19140 => "000011101001111010101101",
19141 => "000010111010011110100101",
19142 => "000000100001001101010101",
19143 => "111110001111100100010101",
19144 => "111011100000000100100011",
19145 => "111000000010101110000111",
19146 => "110101111111101011001101",
19147 => "110110011100110111011110",
19148 => "110111111101010111011010",
19149 => "111001100110011011101111",
19150 => "111100100110110010101010",
19151 => "000001100100110111010011",
19152 => "000111011100010000101110",
19153 => "001101000110001110011000",
19154 => "010001110011011001111000",
19155 => "010101111100010110001100",
19156 => "011001010100010001001001",
19157 => "011010010101111001001100",
19158 => "011001101011110101110100",
19159 => "011000111110011011001111",
19160 => "011000011110000111010010",
19161 => "010111111000111111101000",
19162 => "010110001010111000000100",
19163 => "010011011110110010001000",
19164 => "010001000001001011000110",
19165 => "001110100101011100110100",
19166 => "001011100000001011101001",
19167 => "000111010111001001111100",
19168 => "000011100010111001101100",
19169 => "000001001111110110001101",
19170 => "111110100111101101010101",
19171 => "111011101101001100110000",
19172 => "111010111001001011101011",
19173 => "111100100111100000101110",
19174 => "111111110001001100000011",
19175 => "000010001010100111100010",
19176 => "000010111001001010111111",
19177 => "000011110110001001000100",
19178 => "000101110010010111001100",
19179 => "000111100100001010011111",
19180 => "001001001010110011010000",
19181 => "001011010011101000101000",
19182 => "001100100111101100101000",
19183 => "001010111110101100101100",
19184 => "000110011111001101000110",
19185 => "111111110000101110001110",
19186 => "110110110010011000010101",
19187 => "101101000111011111100100",
19188 => "100101110010001000100101",
19189 => "100010110111000001011011",
19190 => "100011101011000001100111",
19191 => "100101110001011001100101",
19192 => "101000001100011011100000",
19193 => "101100000110001100010010",
19194 => "110001011111111101100000",
19195 => "110110011110010011101100",
19196 => "111010011100001011001011",
19197 => "111110100101010010010000",
19198 => "000011100100000011001101",
19199 => "001000110000000000101101",
19200 => "001100000000000110101110",
19201 => "001011100001111011000100",
19202 => "001000001100110111000110",
19203 => "000011101001001010110110",
19204 => "111110100011110010110110",
19205 => "111010010011011001001011",
19206 => "111000000100111000101100",
19207 => "110111001100111111111110",
19208 => "110111000011010100110010",
19209 => "110110111101000010100001",
19210 => "110101100111100001101100",
19211 => "110100000000001011011101",
19212 => "110011100110111110101110",
19213 => "110011100111011101110100",
19214 => "110011010011100011111000",
19215 => "110011011110110001100000",
19216 => "110100101001100110001010",
19217 => "110100110100101001010110",
19218 => "110010101011010100001010",
19219 => "110001011101001000101000",
19220 => "110011110101110010001110",
19221 => "111000100100100101010100",
19222 => "111110011111111010111001",
19223 => "000110010000101010111010",
19224 => "001110101010100111011110",
19225 => "010011001100001101110110",
19226 => "010010101100011000011110",
19227 => "010000111001111101100100",
19228 => "001111010001000110010110",
19229 => "001100111100110100100110",
19230 => "001001111010101110111001",
19231 => "000111101011111001110001",
19232 => "001000101011011111011011",
19233 => "001100001101100000000100",
19234 => "001111100001101010000110",
19235 => "010010000101100111001000",
19236 => "010101001110111010011000",
19237 => "011000100010110111110001",
19238 => "011001001011101011101011",
19239 => "011000000111111111011001",
19240 => "011000011100110001010001",
19241 => "011000101001101001101111",
19242 => "010111101101000111101010",
19243 => "010101110101101101101000",
19244 => "010001110100101010001000",
19245 => "001101100101101000000010",
19246 => "001010011011100100100000",
19247 => "000110110001111011001110",
19248 => "000101000001100000000101",
19249 => "000110011000010010110011",
19250 => "000110100000011110100010",
19251 => "000100010000111000100010",
19252 => "000001100011001001011111",
19253 => "111110010011100011100100",
19254 => "111010100111100001110000",
19255 => "110110001011000110010101",
19256 => "110001111111110010000110",
19257 => "101111101011110000101000",
19258 => "101010111101011110011000",
19259 => "100011011110101100100011",
19260 => "100000100011000011000010",
19261 => "100001011010000011001110",
19262 => "100001100111110011011111",
19263 => "100010011110010011001011",
19264 => "100011010010100110001001",
19265 => "100011110111010100001100",
19266 => "100111100000110100100011",
19267 => "101101011100000000111110",
19268 => "110010110101001011111000",
19269 => "110111010100100010011011",
19270 => "111010010011011110110000",
19271 => "111011011111111001010010",
19272 => "111011100001011101101100",
19273 => "111010001000101101000110",
19274 => "110111101111110100110011",
19275 => "110101000110111111001110",
19276 => "110001111010001010010110",
19277 => "101110111110010111111110",
19278 => "101101101000110010001010",
19279 => "101101100110110011111100",
19280 => "101110010110100010100110",
19281 => "110000111000111111010000",
19282 => "110110000101010001011000",
19283 => "111010101001010001000100",
19284 => "111011011110010100010100",
19285 => "111011011111111000110100",
19286 => "111101100110110100111111",
19287 => "000001000101111011101110",
19288 => "000100010110101110110111",
19289 => "000110001001001111101100",
19290 => "001000100001010100100110",
19291 => "001101110001010000101100",
19292 => "010010110110010010010100",
19293 => "010100100111011100001010",
19294 => "010101000010001111010110",
19295 => "010110110101010110011010",
19296 => "011001000010110000000001",
19297 => "011001000100110010111111",
19298 => "010101101111001111111100",
19299 => "001111111001101111101110",
19300 => "001010001110110111101110",
19301 => "000110010000110111001010",
19302 => "000011001001000001100000",
19303 => "000000101010010011000000",
19304 => "000000000101000011110100",
19305 => "000001011100111000100100",
19306 => "000010111000000101110110",
19307 => "000011011110101111100100",
19308 => "000100001100110111110110",
19309 => "000101110101000110010000",
19310 => "000111101111100010000110",
19311 => "001000001001110110110110",
19312 => "001000000100011010111001",
19313 => "001001100100101101011110",
19314 => "001011001001001111111000",
19315 => "001100011100000010010110",
19316 => "001101110101001110111110",
19317 => "001101000101011010011000",
19318 => "001010101010011001101010",
19319 => "001000011011110101000111",
19320 => "000101011010101011000011",
19321 => "000000100010001001001001",
19322 => "111011100110011011100000",
19323 => "111001101101101100110110",
19324 => "111010001110101011011000",
19325 => "111010101101100111000010",
19326 => "111011010001111000101001",
19327 => "111100011111000111011111",
19328 => "111110011011011011111100",
19329 => "000000011100001101101100",
19330 => "000001111100010101100111",
19331 => "000011011110000110100100",
19332 => "000100111001000110000010",
19333 => "000110111101010010000000",
19334 => "001001011111001001010110",
19335 => "001010000000111100111100",
19336 => "001001011100001000110010",
19337 => "001001011100000010101000",
19338 => "001000101000001011111100",
19339 => "000110011101101101001010",
19340 => "000100000110110001000100",
19341 => "000011000001010001001001",
19342 => "000011011001110101111111",
19343 => "000011101010001111011010",
19344 => "000010001110011100000111",
19345 => "111101111001111101001110",
19346 => "110111000001000101100000",
19347 => "101111110000010010000010",
19348 => "101001100110011101110010",
19349 => "100101011011110010100111",
19350 => "100100011100110101101111",
19351 => "100110011000101000110111",
19352 => "101001100101110110100100",
19353 => "101101001111001000100110",
19354 => "110001011111100110110100",
19355 => "110110101011101100101011",
19356 => "111100000101010011001001",
19357 => "000000000000111100100001",
19358 => "000010010101101001001101",
19359 => "000011001011001011100111",
19360 => "000000111110000111110000",
19361 => "111100000011111111000001",
19362 => "110111011111110000110110",
19363 => "110100111001001100001110",
19364 => "110011011110111110101010",
19365 => "110011001111000101000100",
19366 => "110101101011010010010101",
19367 => "111010100110111100101000",
19368 => "111110111101111111101100",
19369 => "000000101100001100001000",
19370 => "000001111001111100100100",
19371 => "000101001010101001111111",
19372 => "001001010100110101000111",
19373 => "001100010010100110001010",
19374 => "001110000100010010101000",
19375 => "010001101101101001111000",
19376 => "011000010000010000111001",
19377 => "011100000011011100111100",
19378 => "011011010000100111110010",
19379 => "011010010100000011111000",
19380 => "011001111101000010011000",
19381 => "011001010000110000111011",
19382 => "011000010111001001110110",
19383 => "010111011000110011111110",
19384 => "010111000000001011101000",
19385 => "010110101011100100010100",
19386 => "010110010001101101001100",
19387 => "010011101010001101010000",
19388 => "001011100100010011101001",
19389 => "000001000100001010100100",
19390 => "110111110011100111100000",
19391 => "110000010011001010000110",
19392 => "101010101110111110001100",
19393 => "100101100110000000100011",
19394 => "100001111011111101101111",
19395 => "100001011011100000001011",
19396 => "100010001010110001101001",
19397 => "100101000001000111110101",
19398 => "101011010100100101101000",
19399 => "110011000010010011010010",
19400 => "111011000000011111110011",
19401 => "000001011101110100111101",
19402 => "000011011101011110111010",
19403 => "000001101001100110000001",
19404 => "111110101000101110010011",
19405 => "111010111100101100111100",
19406 => "110110101111110101001111",
19407 => "110010001100101001010110",
19408 => "101101000000000100011110",
19409 => "101000101001001100101000",
19410 => "100101110101111010101010",
19411 => "100011110101010100010011",
19412 => "100011011111101000011011",
19413 => "100100100110011100010010",
19414 => "100101111111110001101111",
19415 => "100111101111110010000001",
19416 => "101000110100000000100100",
19417 => "101000101101110110101100",
19418 => "101000100110010111101010",
19419 => "101000101001111111011010",
19420 => "101001011001101110000110",
19421 => "101100100010101110110010",
19422 => "110010001100110110110110",
19423 => "111000110000011111011100",
19424 => "000000010111010010000111",
19425 => "001001111101110010011110",
19426 => "010010111010100000111000",
19427 => "011000001110101111001011",
19428 => "011011100100001100101001",
19429 => "011110001111001101101011",
19430 => "011110101000011101111100",
19431 => "011110010000111011011011",
19432 => "011110110001011011001001",
19433 => "011100111010111011000011",
19434 => "011000000100110111100111",
19435 => "010011000111111010101000",
19436 => "001110100010000111011100",
19437 => "001010001101111100100110",
19438 => "000110111101111101001111",
19439 => "000101001111101011010010",
19440 => "000100001000100111100111",
19441 => "000001111111000110101011",
19442 => "111111010001110010110110",
19443 => "111101011011011101110111",
19444 => "111101000111111000011001",
19445 => "111110000010110110110001",
19446 => "111111011110111111101100",
19447 => "000001111111100111011101",
19448 => "000100010000100010011101",
19449 => "000100010010101100001001",
19450 => "000011011011101000111101",
19451 => "000010010101111010010101",
19452 => "000000100110101001000001",
19453 => "111110110011100000111111",
19454 => "111100101011010101100110",
19455 => "111001001010010001110010",
19456 => "110011111010101100001110",
19457 => "101111000101110110100110",
19458 => "101100101110111111100110",
19459 => "101011110000100100111000",
19460 => "101011101000010011001010",
19461 => "101100110001111101111100",
19462 => "101110000011011001100100",
19463 => "101110100101101000011100",
19464 => "101111010111100000111100",
19465 => "110000110010001011000110",
19466 => "110001101001000001111010",
19467 => "110010110001001101101100",
19468 => "110101111010101101011001",
19469 => "111001111111001010101011",
19470 => "111101100011110010110100",
19471 => "000000110010011101101110",
19472 => "000100000110110110110111",
19473 => "000111000010010110011110",
19474 => "001001101010000111001100",
19475 => "001101101101101101110000",
19476 => "010010001111000010001000",
19477 => "010100110001101101010010",
19478 => "010101111011001011000110",
19479 => "010110011010110000011000",
19480 => "010101100111001101001100",
19481 => "010011001010011110100100",
19482 => "010000101010001111100000",
19483 => "001111110101010101010100",
19484 => "001111101010001001111010",
19485 => "010000001110001101011100",
19486 => "010010010111011010111010",
19487 => "010100011010001011001000",
19488 => "010101100011111111100010",
19489 => "010110001011000101101000",
19490 => "010110010101100000101110",
19491 => "010101111100111101101100",
19492 => "010100111000000101101000",
19493 => "010100111101011010001110",
19494 => "010110111000000100111000",
19495 => "010111110111111011011000",
19496 => "010110100000111101011010",
19497 => "010011110101111010011000",
19498 => "010000111001010111110010",
19499 => "001110001001000010010000",
19500 => "001011101011000001000100",
19501 => "001000010001101010101100",
19502 => "000010101101111111000111",
19503 => "111100100000011100101000",
19504 => "110111010110010001011100",
19505 => "110011001011010001000010",
19506 => "101111110110111110011000",
19507 => "101101010000001001000010",
19508 => "101011011111010010011010",
19509 => "101010110110110101111100",
19510 => "101011011001100101101010",
19511 => "101101001111001111011010",
19512 => "110000000001000111010010",
19513 => "110011110101101001000100",
19514 => "111001000000101110111011",
19515 => "111110011111000001000010",
19516 => "000011100011001101001011",
19517 => "001000101110111110111001",
19518 => "001110001000111011011110",
19519 => "010011001001110001111010",
19520 => "010110100101110010100110",
19521 => "010111011001100100000110",
19522 => "010110101010111111000110",
19523 => "010101001010101001001000",
19524 => "010000111101000000001100",
19525 => "001001110001101101101100",
19526 => "000000110010010010111001",
19527 => "110110011101000011101001",
19528 => "101101001011111110100100",
19529 => "100110101101100001011101",
19530 => "100010111100010111101110",
19531 => "100010010100011101011001",
19532 => "100100001110011101101011",
19533 => "100111100110001010011011",
19534 => "101011110110011011011010",
19535 => "110000110110110000111010",
19536 => "110110001111001100100000",
19537 => "111010001100111111000110",
19538 => "111100111100001001001101",
19539 => "000000000100011001111100",
19540 => "000011110101011101000100",
19541 => "001000011001100010101110",
19542 => "001101010010001010110010",
19543 => "010001101010101010000000",
19544 => "010011001101010110111100",
19545 => "001111111111110100010110",
19546 => "001011110110111000011000",
19547 => "001001011100001110000100",
19548 => "000110000001011010111000",
19549 => "111111101011100000100010",
19550 => "110111100000010110111000",
19551 => "101111101101100100010110",
19552 => "101000001000100010001110",
19553 => "100010001100101101100101",
19554 => "100001011111110110100001",
19555 => "100010110011111010101110",
19556 => "100011011101111101111101",
19557 => "100111000001101101111110",
19558 => "101110001000011010011100",
19559 => "110111001110011010010000",
19560 => "000000000001101010110101",
19561 => "000101110010010010110010",
19562 => "001010001001101111010111",
19563 => "001111000100100101010000",
19564 => "010011000000011000111110",
19565 => "010100010001001100010100",
19566 => "010010011010110100100000",
19567 => "001110101110111010010100",
19568 => "001011011011110100000011",
19569 => "001000010100000001110010",
19570 => "000011001011001111010001",
19571 => "111101100101011010110101",
19572 => "111011101101111001110010",
19573 => "111101001000011011001101",
19574 => "111110100010111000101011",
19575 => "111111001001011101000001",
19576 => "000000000110011101000001",
19577 => "000010001101101010011010",
19578 => "000100000111000100011010",
19579 => "000011111110000111101111",
19580 => "000010111111010000001001",
19581 => "000010111100101010110010",
19582 => "000010110011101011101111",
19583 => "000001101011110011000001",
19584 => "000000101000111100011111",
19585 => "111111100011001110001100",
19586 => "111101101001010111110101",
19587 => "111100011011010001011110",
19588 => "111101100100010101110111",
19589 => "111111010110101011010011",
19590 => "111111101010110010110000",
19591 => "000000000000100001110111",
19592 => "000000111000001101111100",
19593 => "000000001100001110001101",
19594 => "111110001000100000010011",
19595 => "111011110010000011110111",
19596 => "111000100100000011110101",
19597 => "110011011110000101000010",
19598 => "101101001101000011011110",
19599 => "101000000010000111001010",
19600 => "100100010111111000011011",
19601 => "100010101010100100001101",
19602 => "100011100001100111010011",
19603 => "100100101111011101011001",
19604 => "100110000010100010110111",
19605 => "101000110101000011110010",
19606 => "101100010000111110011000",
19607 => "101111001110100010100100",
19608 => "110001010001100111111000",
19609 => "110011011110000010101010",
19610 => "110110000110101101000101",
19611 => "111000001100101011110001",
19612 => "111010101011100010011001",
19613 => "111100101101100100000111",
19614 => "111100110001001101101011",
19615 => "111100001001001111110100",
19616 => "111011101001110110110100",
19617 => "111100000011000100011111",
19618 => "111101100101110100001110",
19619 => "111111110110111000001110",
19620 => "000011001011101101000110",
19621 => "000110010000001101101000",
19622 => "001000110101111111010100",
19623 => "001100001100100010000100",
19624 => "001110101011000100000010",
19625 => "001111110000001010001110",
19626 => "010001111010011010100010",
19627 => "010101001011100000000000",
19628 => "010110101101110011100010",
19629 => "010110001110100111010100",
19630 => "010101111100100100000100",
19631 => "010101101011100000010010",
19632 => "010100011111111110111110",
19633 => "010011100000110101101000",
19634 => "010011011001000101001010",
19635 => "010011100010101001111000",
19636 => "010100000001100111101010",
19637 => "010101110110110011101100",
19638 => "011000000101100001000100",
19639 => "011000101101010110101111",
19640 => "010111111010100110101110",
19641 => "010110000100100101010010",
19642 => "010011101111000001110000",
19643 => "010001111110001111110010",
19644 => "001111011000101101101110",
19645 => "001010011001010100000011",
19646 => "000100010011101110101010",
19647 => "111111101101000100010110",
19648 => "111101100111011010011000",
19649 => "111100111011100001001011",
19650 => "111100110010100111011100",
19651 => "111101101001110011111100",
19652 => "111111111111101000011100",
19653 => "000010010000100010010100",
19654 => "000010100000110100111110",
19655 => "000010010000011111100000",
19656 => "000010101010000010001101",
19657 => "000001101011000101111001",
19658 => "111110101010110110010000",
19659 => "111011011101001110000110",
19660 => "111001010111001011100000",
19661 => "110111110101000110101010",
19662 => "110101100010100100001001",
19663 => "110010111000101001001010",
19664 => "110010011011001101101110",
19665 => "110101011100100000111010",
19666 => "111001011111111101111110",
19667 => "111100011111111000001001",
19668 => "111101110010001101110000",
19669 => "111011001101100101011111",
19670 => "110101000100100100110100",
19671 => "101110111101100110111110",
19672 => "101010011011100101100110",
19673 => "100111000000010010111001",
19674 => "100101001001100000101100",
19675 => "100110000111000110111101",
19676 => "101001100110001010000000",
19677 => "101110001011110010111100",
19678 => "110010111011001000010110",
19679 => "110110110000100011100101",
19680 => "111001111110000111111010",
19681 => "111101101101110110010010",
19682 => "000001011010101111000111",
19683 => "000100011101001001101000",
19684 => "000111011111101101000101",
19685 => "001010010111111000011100",
19686 => "001010100011001101011000",
19687 => "000110001100000110101001",
19688 => "111111011011110111101011",
19689 => "111010010101000010011010",
19690 => "111001100001010110111010",
19691 => "111011100000000001001011",
19692 => "111100111101001010000000",
19693 => "111110011001100011110001",
19694 => "000001001001011110101110",
19695 => "000011100100011100001011",
19696 => "000100011010000001011101",
19697 => "000101000011101010101101",
19698 => "000110010010001111000001",
19699 => "000110010100110000101000",
19700 => "000101111000010000101001",
19701 => "000110110111101010011011",
19702 => "000111111100110010001100",
19703 => "001000010110101111000101",
19704 => "001000000110101000101010",
19705 => "000111111000001001101111",
19706 => "001001110101001001000011",
19707 => "001101010011101111001000",
19708 => "010001001001001010010110",
19709 => "010100110100110100101110",
19710 => "010110011100001111101110",
19711 => "010110000100110011110010",
19712 => "010100001101100011001100",
19713 => "010000010100100110011000",
19714 => "001011010110011101010111",
19715 => "000111000011100001111010",
19716 => "000100111100101111111000",
19717 => "000100010110001110000100",
19718 => "000100010001111111111011",
19719 => "000101100010010100101010",
19720 => "000111001001100100010011",
19721 => "001000000111101111010000",
19722 => "001001000100010011011000",
19723 => "001001110110101101110111",
19724 => "001010001100000110100001",
19725 => "001001001101111001001100",
19726 => "000101110101010010110111",
19727 => "000000001110011010011000",
19728 => "111001011001010001100000",
19729 => "110011001011000110101110",
19730 => "101110111001001100101110",
19731 => "101100000011010000100000",
19732 => "101010000001100101111110",
19733 => "101001000111011110101000",
19734 => "101001011100000110111100",
19735 => "101010100111101010111010",
19736 => "101100101011110001100110",
19737 => "101111011000100100001100",
19738 => "110001110111000001110100",
19739 => "110011110001111000110000",
19740 => "110100100110100101011100",
19741 => "110011000111100000011000",
19742 => "101111101000001100001100",
19743 => "101100001010111000011110",
19744 => "101001011010100110001100",
19745 => "100110110100110000010110",
19746 => "100101010100100100010001",
19747 => "100101100111110000101110",
19748 => "100110010101000100111101",
19749 => "100110111001001100111011",
19750 => "101001100110001100010000",
19751 => "101111011000110010011110",
19752 => "110101111000001100001100",
19753 => "111100100110001000101111",
19754 => "000100010011000000000010",
19755 => "001011011011000101101100",
19756 => "010001001000101010010110",
19757 => "010100111111001100100100",
19758 => "010110011010011001110110",
19759 => "010110001111011100010000",
19760 => "010101010001101100101100",
19761 => "010100110000010100101010",
19762 => "010100001101011001010110",
19763 => "010001110011011001011010",
19764 => "001110111000111010010110",
19765 => "001100011010000100000010",
19766 => "001001110101100010101100",
19767 => "000111111010001001000010",
19768 => "000110111001101100111111",
19769 => "000111000010011001001011",
19770 => "001000010110110010111000",
19771 => "001010100101010000001011",
19772 => "001100111100100000011010",
19773 => "001101101011001000001110",
19774 => "001101011100001111110100",
19775 => "001101101101001010011100",
19776 => "001110010010010110000000",
19777 => "001111010010101101101110",
19778 => "010000011100000011110110",
19779 => "010010000101000100110000",
19780 => "010011100111011100110000",
19781 => "010010100001101001000110",
19782 => "001111011100101010100010",
19783 => "001100000110010110111000",
19784 => "001000100111110011110101",
19785 => "000101000001011010011111",
19786 => "000000001011011011011100",
19787 => "111001010001011010010011",
19788 => "110000000101001101001010",
19789 => "100110011011011001010100",
19790 => "100001011101011101111110",
19791 => "100001100010110010110111",
19792 => "100001110000110101110011",
19793 => "100001000110001101011010",
19794 => "100001001100110100100111",
19795 => "100010000101010111011010",
19796 => "100011011011000111111111",
19797 => "100100010001110011010100",
19798 => "100100101110110100000110",
19799 => "101000000100110101110110",
19800 => "101110100110110010110000",
19801 => "110100110010001111011111",
19802 => "111011001001110001100000",
19803 => "000011000101011111101111",
19804 => "001001111001101010101100",
19805 => "001110010010001100101000",
19806 => "010001000010001001010000",
19807 => "010010011111101010100110",
19808 => "010100001000000010000010",
19809 => "010110011001100100011000",
19810 => "010110010010011010110100",
19811 => "010010011101101101101100",
19812 => "001101110111101000001100",
19813 => "001001101000011011010010",
19814 => "000100001000100000100110",
19815 => "111110001000000011001011",
19816 => "111001111101010110100100",
19817 => "111000000100110101000110",
19818 => "111000000101001001110100",
19819 => "111010010000000011111100",
19820 => "111101001001110010100010",
19821 => "111101111011101001111101",
19822 => "111100101111011001111000",
19823 => "111101001000101110001000",
19824 => "000010001101101000001010",
19825 => "001001110100010000011101",
19826 => "001111010010010110011000",
19827 => "010011111110011111110100",
19828 => "011010000101101011101110",
19829 => "011101000001100000110110",
19830 => "011000111110001001010101",
19831 => "010000111110001011111110",
19832 => "001001110111101100010110",
19833 => "000011110111100100100001",
19834 => "111100100000110110111001",
19835 => "110100010110011101111100",
19836 => "101101011100111111001000",
19837 => "101001000101010010010000",
19838 => "100110100101000000110101",
19839 => "100100000010110111110011",
19840 => "100011100011011100001011",
19841 => "101000000001000000100010",
19842 => "101110111000001001110100",
19843 => "110100010011110100111000",
19844 => "111000001000011110111010",
19845 => "111100001110110100111111",
19846 => "000000110010010000110100",
19847 => "000100001101010000010111",
19848 => "000110001000011111011101",
19849 => "000111101010011111110100",
19850 => "001001100000000110110110",
19851 => "001011000100001000001010",
19852 => "001100010010110111001010",
19853 => "001101111001100110011110",
19854 => "001110101100011010010010",
19855 => "001101000110010111101110",
19856 => "001001110110101001001110",
19857 => "000110110010100000000110",
19858 => "000100000010100000001010",
19859 => "000000010100101101011000",
19860 => "111100011111100011101110",
19861 => "111010000000111001010010",
19862 => "111000100100101010111011",
19863 => "111000011110101000010010",
19864 => "111010011101100111001100",
19865 => "111110010001011111010000",
19866 => "000010100100101111101101",
19867 => "000101110110000111110100",
19868 => "000111110011111111110101",
19869 => "000111111010110010111100",
19870 => "000101111111011110010000",
19871 => "000011101010001111100011",
19872 => "000001111011101011011001",
19873 => "000000110110011101100100",
19874 => "111111111100010010010101",
19875 => "111110000110100111101100",
19876 => "111010101110010110101111",
19877 => "110110100101101101101100",
19878 => "110011010111100100011000",
19879 => "110000110111100011111100",
19880 => "101110010010011000001110",
19881 => "101100111001100001100100",
19882 => "101100111100000000011100",
19883 => "101101011101101111010010",
19884 => "101110011010100001111100",
19885 => "101111100001100110011100",
19886 => "110001001000101100110110",
19887 => "110011101111000011110100",
19888 => "110110001100010110011001",
19889 => "110111100101110101010101",
19890 => "111000101001100000011011",
19891 => "111010000111101110111111",
19892 => "111011100111011101110001",
19893 => "111100110011001101010000",
19894 => "111110011111111100100111",
19895 => "000001101011001101010011",
19896 => "000101101110101110101110",
19897 => "001001010010111011011010",
19898 => "001100011010111010111010",
19899 => "001111010011100110110110",
19900 => "010000111111000000011110",
19901 => "010001010100100110000000",
19902 => "010001001111110100111100",
19903 => "010001000001010100001000",
19904 => "010000000001011101010100",
19905 => "001110001111100100101100",
19906 => "001100111010000101111110",
19907 => "001100101110011110101110",
19908 => "001100111111000001100110",
19909 => "001100111010011000111010",
19910 => "001101010011010110001010",
19911 => "001111101111001101110110",
19912 => "010100000110001010001100",
19913 => "011000010011110110001110",
19914 => "011010010001011001111011",
19915 => "011010000100000000110111",
19916 => "011001011011111110101011",
19917 => "011001000110001000011001",
19918 => "011000110000001100111111",
19919 => "011000000010101110111001",
19920 => "010111010101101000111110",
19921 => "010110101111011100001010",
19922 => "010011110001101011110100",
19923 => "001101011011101011111110",
19924 => "000101011110011000110010",
19925 => "111100100100000100000000",
19926 => "110011100010010100010110",
19927 => "101011001100110011011000",
19928 => "100100011111000110111111",
19929 => "100001101101101111001100",
19930 => "100001110100100010111111",
19931 => "100001101010011100010011",
19932 => "100001010100101001011111",
19933 => "100001110010001011100001",
19934 => "100010101101111101100000",
19935 => "100011100110101111110011",
19936 => "100100001001000101101111",
19937 => "100011111000001110001111",
19938 => "100100011010111010100101",
19939 => "101001000010010001100000",
19940 => "110000010011010001010100",
19941 => "110110010110001010111111",
19942 => "111010101110011110001010",
19943 => "111101010111110110001000",
19944 => "111110010111101100011010",
19945 => "111111100100001101101000",
19946 => "000001100011100100110111",
19947 => "000010111110000111110000",
19948 => "000010100110101111001101",
19949 => "000001100111010001100100",
19950 => "000010001111011101000001",
19951 => "000100010011001101111101",
19952 => "000101011010100011101111",
19953 => "000011101000000110001010",
19954 => "000000000001110001001011",
19955 => "111101100000000011110000",
19956 => "111100011100100001010100",
19957 => "111100010110101001100000",
19958 => "111110001100111011011011",
19959 => "000001100100010100111000",
19960 => "000100011111011110101100",
19961 => "000111000001111100011000",
19962 => "001011010010110100011111",
19963 => "010001001100001100011100",
19964 => "010101010001010111010000",
19965 => "010110100101000110101000",
19966 => "011000001110010110101010",
19967 => "011010110111111110011110",
19968 => "011100010011001000110111",
19969 => "011011110110010010000101",
19970 => "011010101001110001110101",
19971 => "011010001010011110011111",
19972 => "011001000100011001010111",
19973 => "010100101001010111000100",
19974 => "001111000100111110111000",
19975 => "001011010111111111100110",
19976 => "001000010101000001100000",
19977 => "000101010110101000001010",
19978 => "000010101001110011001110",
19979 => "111111000101001101011100",
19980 => "111010111000101001011001",
19981 => "110111010000001001110100",
19982 => "110100100001101011100001",
19983 => "110011010111001010011000",
19984 => "110100101111101101000001",
19985 => "111000011000101101101110",
19986 => "111100100011001100101010",
19987 => "111111111110111111111111",
19988 => "000011000101111100101010",
19989 => "000101011111000000010000",
19990 => "000101011010101110011100",
19991 => "000011111110001000011101",
19992 => "000010010110110010001111",
19993 => "111110001010110011100110",
19994 => "110111011001011110111010",
19995 => "101111101111011111011010",
19996 => "100111100110101001011001",
19997 => "100010100010000101001111",
19998 => "100001111010110011101101",
19999 => "100010000111101111001111",
20000 => "100001111100101111101110",
20001 => "100001100000010000101100",
20002 => "100001110101000000110001",
20003 => "100101111011001000010011",
20004 => "101100100110111110111000",
20005 => "110010111101100100100010",
20006 => "111001000111111001010111",
20007 => "111110111100010000101011",
20008 => "000011111001111100010010",
20009 => "000111110111100001111000",
20010 => "001001011010100001010010",
20011 => "000111110100101010000011",
20012 => "000011100101110011100101",
20013 => "111101000110101011100100",
20014 => "110110110100111111001000",
20015 => "110100000011101101110011",
20016 => "110011110110110010011100",
20017 => "110011000011001011100110",
20018 => "110001010111011011100100",
20019 => "110000101010100110010000",
20020 => "110001011110101101011100",
20021 => "110010100011000011101110",
20022 => "110011011001000000111010",
20023 => "110100101111110111001100",
20024 => "110110111011010010001110",
20025 => "111010001110101001111110",
20026 => "111111000000011000010001",
20027 => "000100010101110100011101",
20028 => "001000011110110001011010",
20029 => "001011100001101000001110",
20030 => "001111011010000100010000",
20031 => "010011011001101010111110",
20032 => "010101001000010101111100",
20033 => "010101001111100010001110",
20034 => "010100111101111011101100",
20035 => "010011101101011111100100",
20036 => "010001010101101101101110",
20037 => "001110110011001001001000",
20038 => "001100110111100011001100",
20039 => "001011001100010101010111",
20040 => "001001011000010101011100",
20041 => "001000010000001001110011",
20042 => "001000010001011110100110",
20043 => "001001000010001110001011",
20044 => "001010011111011100101111",
20045 => "001101001110111110010010",
20046 => "010001110101010011101110",
20047 => "010110110101001111110010",
20048 => "011001011000100101100101",
20049 => "011001010111011110111011",
20050 => "011000101100111101001001",
20051 => "011000000110111010000101",
20052 => "010111010111110100000100",
20053 => "010101010111111001100010",
20054 => "010001111011001010000110",
20055 => "001111000001011110101000",
20056 => "001011110001001101000100",
20057 => "000110001011000111110001",
20058 => "000000110001000001010111",
20059 => "111101001001001110010001",
20060 => "111010001100110000111010",
20061 => "110111110000000110111000",
20062 => "110100010001011010011110",
20063 => "101111101011001111001110",
20064 => "101100100010001010000010",
20065 => "101001010101000100011000",
20066 => "100100111001110110010101",
20067 => "100010111001011010100001",
20068 => "100011001001000110110000",
20069 => "100010101010010001111111",
20070 => "100010011101100111111111",
20071 => "100011001100110101001111",
20072 => "100011101110111001011111",
20073 => "100100011101110110101101",
20074 => "100101100011001111011111",
20075 => "100110011100000001000010",
20076 => "100110101101110001110000",
20077 => "100110110100010110010001",
20078 => "101001011110110100000000",
20079 => "101111001000011111101000",
20080 => "110100000110100011101001",
20081 => "110111000111111111111000",
20082 => "111000111101000000011010",
20083 => "111000101111000011011000",
20084 => "110111010111010011001010",
20085 => "110111001000100111000110",
20086 => "110111001010011101100010",
20087 => "110110010110101111111110",
20088 => "110110101101100111110100",
20089 => "111000101000100001011000",
20090 => "111001111111001100001101",
20091 => "111010111110010100110111",
20092 => "111101110100110110000011",
20093 => "000011100100010000110101",
20094 => "001010011000001110111101",
20095 => "001110101010011011101100",
20096 => "001111111111111011110110",
20097 => "010001011010101010101000",
20098 => "010011011011011101101000",
20099 => "010011111110110010100110",
20100 => "010010111100011110111110",
20101 => "010001100100001011011110",
20102 => "010000101011111111110000",
20103 => "010001000111000101101010",
20104 => "010001110011110101010110",
20105 => "010000001111000111100010",
20106 => "001101000011111101011010",
20107 => "001011000011110111110000",
20108 => "001001110001100111000101",
20109 => "000111111111101000111111",
20110 => "000111101101100110010111",
20111 => "001001110111001011111011",
20112 => "001011101010010001100001",
20113 => "001011010110000001111000",
20114 => "001010001000011011111010",
20115 => "001001000000011000010110",
20116 => "000111100110101110010000",
20117 => "000110001010101110000110",
20118 => "000101111100001100011001",
20119 => "000111000101011111111100",
20120 => "001000000010101101110010",
20121 => "000111100100001110001110",
20122 => "000101111110110011011000",
20123 => "000100000010110111011100",
20124 => "000001100010011000110111",
20125 => "111110010000111111110101",
20126 => "111011010010100100001111",
20127 => "111001001010001000111000",
20128 => "110111000100101110001110",
20129 => "110101000000100011111111",
20130 => "110011110001110011111000",
20131 => "110011011101011001001100",
20132 => "110011111111001100101010",
20133 => "110101110000000000111100",
20134 => "111000101000001001011011",
20135 => "111011111100001010101110",
20136 => "111111011011100001000110",
20137 => "000010111101101000101110",
20138 => "000101010001100010100111",
20139 => "000101000100111001100000",
20140 => "000011010011000111101101",
20141 => "000001101110001111010101",
20142 => "000000101000100000010111",
20143 => "111111110001000001110001",
20144 => "111111011010010001000111",
20145 => "111111111100010111110100",
20146 => "000001100111100110001001",
20147 => "000011110010110000111101",
20148 => "000101001010111011111101",
20149 => "000101111100101010111111",
20150 => "000111001001000111110100",
20151 => "001000100111001101101100",
20152 => "001001101110100000001000",
20153 => "001001101101100010011000",
20154 => "000111011100101111001110",
20155 => "000010101001000110111001",
20156 => "111100010010101001001010",
20157 => "110101011100110001011111",
20158 => "101111001001001000001000",
20159 => "101011010010001111101000",
20160 => "101010101001000010110100",
20161 => "101011101000111101101110",
20162 => "101101011101010111101100",
20163 => "110000110110110110100110",
20164 => "110101101110100010001000",
20165 => "111010101011100000001110",
20166 => "111111001001110010011001",
20167 => "000011110010111000011010",
20168 => "001000001000100001101001",
20169 => "001011000000011001011111",
20170 => "001101000111101100100100",
20171 => "001111101101110010100110",
20172 => "010001101111011100100110",
20173 => "010001010101010010111110",
20174 => "001110100001011111111110",
20175 => "001010100111101110101111",
20176 => "000111010011000110001010",
20177 => "000101100000001101111000",
20178 => "000100100111111100000111",
20179 => "000100011010111110001100",
20180 => "000101000011110001111001",
20181 => "000110011100010100001101",
20182 => "001000101101110100100010",
20183 => "001011100100100000111011",
20184 => "001111000010111010001010",
20185 => "010010011001111111010000",
20186 => "010011110010110111010100",
20187 => "010100100101000110010010",
20188 => "010110011001000011111000",
20189 => "010111000110001000111100",
20190 => "010110011001100011001100",
20191 => "010110000111101000001110",
20192 => "010101110001111111001100",
20193 => "010101010111111000010110",
20194 => "010100010000111010100100",
20195 => "001111000011010011100000",
20196 => "000111011110011100011100",
20197 => "000010101110001000001001",
20198 => "111111010100001011101101",
20199 => "111001110011010000000100",
20200 => "110010011011111110001110",
20201 => "101010110011101000011110",
20202 => "100101100001000101011001",
20203 => "100011100110011111000101",
20204 => "100011101110011101001011",
20205 => "100101111101011001111010",
20206 => "101010010010011110010010",
20207 => "101111010101011001000010",
20208 => "110100101111000011001000",
20209 => "111010000000001110111111",
20210 => "111101000000101111111011",
20211 => "111100001001011010011001",
20212 => "111000110110111101001100",
20213 => "110110000100100100101101",
20214 => "110010010111010111101100",
20215 => "101010011110011001110100",
20216 => "100010111111110110111111",
20217 => "100001101111000100011100",
20218 => "100010110111101110101001",
20219 => "100010100100001111000011",
20220 => "100010101110011101100001",
20221 => "100011011100110111100011",
20222 => "100100000110001000110011",
20223 => "100101001000001000001110",
20224 => "100101111011000100100010",
20225 => "101000000111110111100100",
20226 => "101101111100000101110110",
20227 => "110101001000011111010000",
20228 => "111011011011101011010000",
20229 => "000001000110111011010111",
20230 => "000101101001000011011100",
20231 => "001001100000100010100110",
20232 => "001101111101111000000110",
20233 => "010001010000001011001100",
20234 => "010010011100011001011000",
20235 => "010011110100000001000110",
20236 => "010110100101111110111010",
20237 => "011001011110001001100110",
20238 => "011001101000110001001001",
20239 => "010110110001011110100110",
20240 => "010100001000011011100000",
20241 => "010010100111101110000010",
20242 => "010000110100011111111010",
20243 => "001110110111010000001110",
20244 => "001101011100001001100010",
20245 => "001101000000101100101010",
20246 => "001101101101010010100100",
20247 => "001110001010010001100010",
20248 => "001100101100011011000100",
20249 => "001010000000101101001101",
20250 => "000111011010111110110010",
20251 => "000100111001111100101101",
20252 => "000011010111001000110011",
20253 => "000011011110001010011110",
20254 => "000100100111011110000000",
20255 => "000110011001000000110110",
20256 => "000111011100111000000000",
20257 => "000110010110010001111010",
20258 => "000011001000111000111110",
20259 => "111111000111110000100110",
20260 => "111011110011011000000011",
20261 => "111000110110101111011001",
20262 => "110101010010001111011100",
20263 => "110001000111001011111010",
20264 => "101101001110100110101000",
20265 => "101010001011110100110100",
20266 => "100110101101000011001101",
20267 => "100011000111000000100111",
20268 => "100001111001011001111100",
20269 => "100010110101101100111000",
20270 => "100011110011110011001100",
20271 => "100100011011101101100001",
20272 => "100101100011101001000001",
20273 => "100110011111010111001101",
20274 => "100110010011100010111101",
20275 => "100110011100110100011111",
20276 => "100111110000111001101111",
20277 => "101001110100010010111110",
20278 => "101101001111001111101110",
20279 => "110001111001110111100010",
20280 => "110110100100000001010000",
20281 => "111010110000100001110101",
20282 => "111110001010101000111100",
20283 => "000000000010000011100101",
20284 => "000000110110001011010101",
20285 => "000010000001011011010001",
20286 => "000011011010011100010111",
20287 => "000100001110000000101010",
20288 => "000100110011100010001100",
20289 => "000101101100000111100101",
20290 => "000111000111000111110110",
20291 => "001000111000101110111111",
20292 => "001010010100000001100011",
20293 => "001100000001100111111110",
20294 => "001111010100000010001100",
20295 => "010011010110010010010010",
20296 => "010101110101111000111100",
20297 => "010101111001111100110110",
20298 => "010101011000011101100110",
20299 => "010101110111111101011100",
20300 => "010110010001111010000100",
20301 => "010101101100000011000000",
20302 => "010100101001000001011000",
20303 => "010011100111001001011100",
20304 => "010010101101101000101100",
20305 => "010001110001100100111000",
20306 => "010000101101101101110010",
20307 => "001111111001101100000010",
20308 => "010000000000100001001000",
20309 => "010000100001111010100100",
20310 => "010000100011011001011010",
20311 => "010000110001001110000000",
20312 => "010000011110101101101110",
20313 => "001110010011111010000100",
20314 => "001100000011001101110100",
20315 => "001011011111100001100100",
20316 => "001100000110111011100010",
20317 => "001100101010110001000110",
20318 => "001100001101011101110010",
20319 => "001010110110011111011110",
20320 => "001000101100001001110110",
20321 => "000100000111100110101110",
20322 => "111101000011100110100011",
20323 => "110111000101010110111110",
20324 => "110011110010100000010110",
20325 => "110001101011011011110110",
20326 => "110000110101110110011010",
20327 => "110001101011010010110110",
20328 => "110010111100000101100010",
20329 => "110011010010100010000010",
20330 => "110011011001000110111010",
20331 => "110100110001000010101111",
20332 => "110110110010110110001100",
20333 => "111000100110110000000000",
20334 => "111010001100000000000110",
20335 => "111010111010110000011001",
20336 => "111010100000110000010111",
20337 => "111010010000011001001000",
20338 => "111011000001010011011000",
20339 => "111011000101001000101100",
20340 => "111010011111110000101000",
20341 => "111011101000000011011011",
20342 => "111101101011000111001101",
20343 => "111110100110100101010011",
20344 => "111110101101010100011111",
20345 => "111111011011010111101011",
20346 => "111111111000011001111001",
20347 => "111110100011111011100010",
20348 => "111101001011010010101100",
20349 => "111100101000000001001010",
20350 => "111100100111010010010000",
20351 => "111101000111100000000001",
20352 => "111101100001101110000110",
20353 => "111110101111001111101011",
20354 => "111111111111101100111111",
20355 => "111111011010000101110010",
20356 => "111101110001111111000111",
20357 => "111011101010001000011101",
20358 => "111000011011000101110001",
20359 => "110011111000010111110000",
20360 => "101111111100101000101010",
20361 => "101110101101100010101000",
20362 => "101111111110011010000010",
20363 => "110011010101110111110110",
20364 => "110111001110000000000111",
20365 => "111001111101011011000100",
20366 => "111100100000000011010000",
20367 => "000000000100000001010000",
20368 => "000011101100011000010100",
20369 => "000101111100010110100000",
20370 => "001000100100001110000000",
20371 => "001100001110010111001100",
20372 => "001111001110100000001100",
20373 => "010010101100011000100100",
20374 => "010110011100100110001110",
20375 => "011000000000101101111111",
20376 => "010111100100110110101100",
20377 => "010111001111011010110110",
20378 => "010111111001110000000000",
20379 => "011000001111011100011100",
20380 => "010110001101100101101100",
20381 => "010000101101110111100100",
20382 => "001010000100111100000010",
20383 => "000101000001101111111110",
20384 => "000000101011010101100100",
20385 => "111101011111011001111001",
20386 => "111100011100111001011001",
20387 => "111011100001011000001100",
20388 => "111010110110000010111111",
20389 => "111110000010011100101100",
20390 => "000100101001011011010011",
20391 => "001000111001000010001100",
20392 => "001000111011100011110110",
20393 => "000110100011000100101100",
20394 => "000010110110000100100111",
20395 => "111111111110000010001010",
20396 => "111101110110011001111110",
20397 => "111011010101001100110101",
20398 => "111000101110000010111001",
20399 => "110101111101110000100010",
20400 => "110011101011000011101000",
20401 => "110001110100011011011100",
20402 => "110000110111001010101110",
20403 => "110001110011011100101000",
20404 => "110011011111011001001110",
20405 => "110101001111100110101100",
20406 => "110111000011000110001001",
20407 => "110111110001000101001001",
20408 => "110101010101111011110010",
20409 => "101111110011011100001000",
20410 => "101010101110010110111110",
20411 => "101000011011000011100110",
20412 => "101000001000100010010010",
20413 => "100111010100001001111101",
20414 => "100101010110100000011111",
20415 => "100100110101001101010001",
20416 => "100110001001110010001011",
20417 => "101000001001111101100000",
20418 => "101010011001001001010100",
20419 => "101100101101110111011100",
20420 => "101111111111110011111010",
20421 => "110100001000100111111111",
20422 => "111000000001001111011101",
20423 => "111011001010100111100100",
20424 => "111101001000100111011101",
20425 => "111101010001100100111010",
20426 => "111011111110111001011011",
20427 => "111011010000100000110110",
20428 => "111100011110100101010110",
20429 => "111111000110111011111011",
20430 => "000001111101000000010000",
20431 => "000100111111101100100001",
20432 => "001000011101100111001001",
20433 => "001011100110010010100100",
20434 => "001101111101000010100010",
20435 => "001110110100100111100100",
20436 => "001110001100001101011000",
20437 => "001101100001011000010010",
20438 => "001101110101110001111110",
20439 => "001110011001111101111100",
20440 => "001100110001111010010000",
20441 => "001001100101110110011110",
20442 => "000111100011000110100101",
20443 => "000111001011001010101100",
20444 => "001000110101101010010001",
20445 => "001011101001100011110111",
20446 => "001110001000100010101000",
20447 => "001111100010101101110100",
20448 => "001111011110111110110100",
20449 => "001111100111111101101010",
20450 => "010000011011000000110100",
20451 => "010000111010001100001010",
20452 => "010000111101011001001010",
20453 => "010000110000000100010010",
20454 => "010000011100110011010010",
20455 => "001111000100011101111000",
20456 => "001100110100000001100110",
20457 => "001010101000000001001110",
20458 => "001001010010001111100100",
20459 => "001001110110101000111101",
20460 => "001010100111000001101010",
20461 => "001010011111000011101100",
20462 => "001001111010001111111010",
20463 => "001000101000110010010000",
20464 => "000110111011000111101111",
20465 => "000011011111010011101111",
20466 => "111110010001110100100100",
20467 => "111001001000001011001110",
20468 => "110100110010011101001010",
20469 => "110001100101001101111100",
20470 => "101110010101101111011010",
20471 => "101011000110001010110010",
20472 => "101010100100100111011110",
20473 => "101101111000010010011010",
20474 => "110011000100110010000000",
20475 => "111000101101111011100000",
20476 => "111111001111111110101100",
20477 => "000101001101001001100110",
20478 => "001001001111100000111001",
20479 => "001011110000101111011010",
20480 => "001101000011111111110000",
20481 => "001110000010111010111100",
20482 => "001101111101101010111100",
20483 => "001011110111011000101111",
20484 => "000111001100011111111010",
20485 => "111111011110010011110101",
20486 => "110111010010110110010110",
20487 => "101111110100001001101010",
20488 => "101000110000011100001100",
20489 => "100100000001100111110101",
20490 => "100010110011011100111011",
20491 => "100011110010000000100111",
20492 => "100101001100110010100111",
20493 => "101000101011001010011010",
20494 => "101110111100011101110000",
20495 => "110101010000111000000001",
20496 => "111010000110011010001100",
20497 => "111110000100111101100011",
20498 => "000100000100110011101101",
20499 => "001010101101011110100000",
20500 => "001100010010100111111100",
20501 => "001000111101000010001001",
20502 => "000011111100101010000110",
20503 => "111110101000000101111100",
20504 => "111001001100110110101011",
20505 => "110101100010110111110101",
20506 => "110101110010011001101110",
20507 => "110111100001001011011001",
20508 => "111001000110000100111001",
20509 => "111010100000101000010000",
20510 => "111010111001101101011000",
20511 => "111011100100011101110111",
20512 => "111101100001100011010101",
20513 => "000000011011100111000010",
20514 => "000011100100111000001100",
20515 => "000111010101101110011101",
20516 => "001100110100001010001000",
20517 => "010001111000001001001110",
20518 => "010101100011000100100100",
20519 => "011001011101000110010101",
20520 => "011100100000000011111001",
20521 => "011100100111111000101001",
20522 => "011011000000101100001000",
20523 => "011010010010101101111001",
20524 => "011001111101111110010011",
20525 => "011000111011111000010100",
20526 => "011000010011011000101000",
20527 => "010111110011111101001100",
20528 => "010100101000110110000100",
20529 => "001100111001111110101010",
20530 => "000011110010011000101100",
20531 => "111101001000111101110000",
20532 => "111000000000010100111001",
20533 => "110011011110101011010000",
20534 => "110000111101011111001010",
20535 => "110000011001111100110100",
20536 => "110000100011111110011000",
20537 => "110010000001101010110010",
20538 => "110101011010000000110010",
20539 => "111001001101011100011100",
20540 => "111101000010100011011001",
20541 => "000000100001010000100010",
20542 => "000001011000010011100010",
20543 => "111110011100101111100110",
20544 => "111001000011110010111011",
20545 => "110011101101110111000100",
20546 => "101111011011110101100110",
20547 => "101100011010100101011100",
20548 => "101010100100100110110010",
20549 => "101000001001101100111000",
20550 => "100101001111010111110001",
20551 => "100011111111000001110001",
20552 => "100100101101001011000100",
20553 => "100110011010100000101001",
20554 => "101000100100100101100110",
20555 => "101011001110101001110110",
20556 => "101110000011111101100000",
20557 => "101111100110111001101110",
20558 => "101110010001101100010110",
20559 => "101011010110011101010000",
20560 => "101010000101001001100110",
20561 => "101010001100110001010110",
20562 => "101010011110101100100110",
20563 => "101101010011000001001100",
20564 => "110100010000111011010000",
20565 => "111110010001001001101111",
20566 => "001001000000110110011100",
20567 => "010001111010101100100000",
20568 => "011001000111110101101101",
20569 => "011110001001010000111111",
20570 => "011110110000111010110110",
20571 => "011110000011110110011011",
20572 => "011110100010110100010100",
20573 => "011110001010000010011110",
20574 => "011101111110010111110111",
20575 => "011101101111010111100101",
20576 => "011010000110111110111101",
20577 => "010100011101011101010000",
20578 => "010000011011100101010100",
20579 => "001110101001100101110100",
20580 => "001101111110110010001110",
20581 => "001110001000101100100010",
20582 => "001110000011000011000010",
20583 => "001100001110010101010010",
20584 => "001001110101000000101111",
20585 => "001000101111111111101010",
20586 => "001010010000011101101111",
20587 => "001101000110100101101110",
20588 => "001110101011101001110110",
20589 => "001111100010001101101000",
20590 => "010000011011100101000100",
20591 => "010000101100101000101110",
20592 => "001110101101000001000100",
20593 => "001010111110001110011110",
20594 => "001000110000010101100100",
20595 => "000110010111000111010011",
20596 => "000010001011100100011110",
20597 => "111101101101110000011110",
20598 => "111000010100000010010011",
20599 => "110011000010110001001100",
20600 => "101101010001011111011010",
20601 => "100110000000101001110011",
20602 => "100001110101011100000111",
20603 => "100001011001001000010001",
20604 => "100001010011011001011001",
20605 => "100001010010011100010111",
20606 => "100001110011101111010001",
20607 => "100010110110000001110111",
20608 => "100100001011100101110101",
20609 => "100100110010100101101001",
20610 => "100101111110011110100101",
20611 => "101100011100111000111010",
20612 => "110110101100100110111000",
20613 => "111110000011001100111110",
20614 => "000011101010011000101110",
20615 => "001010000110011001001011",
20616 => "001110101000100110010100",
20617 => "010000001101101100101000",
20618 => "010000000101111001101110",
20619 => "001111101111101111100110",
20620 => "001110110010110101101010",
20621 => "001100001110101101011000",
20622 => "001001100010010001000010",
20623 => "000110111100111101111100",
20624 => "000100101001001000100010",
20625 => "000101001010000001010111",
20626 => "001000100001000011111101",
20627 => "001010110110110111101011",
20628 => "001010000110011100111110",
20629 => "001001110011001000101010",
20630 => "001011111010110101000000",
20631 => "001100100100101111011010",
20632 => "001010110101000001100100",
20633 => "001011000001101000000100",
20634 => "001110111001010110111000",
20635 => "010010010010001111110100",
20636 => "010010111010011111011000",
20637 => "010100111110011001100010",
20638 => "011001001000110011000111",
20639 => "011010001010111001100111",
20640 => "010111010111111100000000",
20641 => "010100111110110001000110",
20642 => "010011110001100000011100",
20643 => "010000101010010100010000",
20644 => "001001111000100001101010",
20645 => "111111011011001000110000",
20646 => "110100010100110000110001",
20647 => "101100001010111000110110",
20648 => "100101101101010110011101",
20649 => "100001101110111110110111",
20650 => "100010000001000000000000",
20651 => "100010101011010001111111",
20652 => "100010000100001110010110",
20653 => "100010000000001000000010",
20654 => "100010101011000100001001",
20655 => "100011010101110110101111",
20656 => "100101000111001100010000",
20657 => "101010110110000100100010",
20658 => "110011101111110111111110",
20659 => "111101101001000110010011",
20660 => "000111110000010011101000",
20661 => "010000100100001100010000",
20662 => "010111011000011000001110",
20663 => "011010101111000000110110",
20664 => "011010001000100111001011",
20665 => "011000011010001100010111",
20666 => "010111100110001001111110",
20667 => "010101100111011011011010",
20668 => "001101101101010111011010",
20669 => "000001100110110111100011",
20670 => "110111000011011010100111",
20671 => "101111010011010000101100",
20672 => "101010101001101111110110",
20673 => "101000010110101011001010",
20674 => "101000010000000110011000",
20675 => "101011011001010100110010",
20676 => "110000000101101000000110",
20677 => "110100101011101011011000",
20678 => "110111011001101101101011",
20679 => "111000101110000101111010",
20680 => "111010111110010100000110",
20681 => "111101011011011111010101",
20682 => "000001000001011110011000",
20683 => "000110101011111011101000",
20684 => "001100100110001001001000",
20685 => "010001000001010001110000",
20686 => "010001110100010010100010",
20687 => "001111101111110101101110",
20688 => "001101010111100011111000",
20689 => "001010111010100101000010",
20690 => "001000001111010101101011",
20691 => "000101010100101010101101",
20692 => "000000111100111101000110",
20693 => "111001100011101011100100",
20694 => "110000001110110100000010",
20695 => "100111111000000010010001",
20696 => "100010111100011010001001",
20697 => "100010100110011100100101",
20698 => "100011111010111110110010",
20699 => "100100101011001011001011",
20700 => "100111111011111001110111",
20701 => "101110101000111010001000",
20702 => "110101010101111000010111",
20703 => "111010101010011101000101",
20704 => "111111101111100101001101",
20705 => "000100111000100000011111",
20706 => "001001001011011000101010",
20707 => "001100001100010101011000",
20708 => "001110110001011111000010",
20709 => "010000010000010010011110",
20710 => "001111001101111011100110",
20711 => "001100101100110111101000",
20712 => "001001110100001101110100",
20713 => "000111100000000000001010",
20714 => "000110011110111011101001",
20715 => "000110101110011101011110",
20716 => "001000101010111110100100",
20717 => "001010111111010100000100",
20718 => "001100110111101011100110",
20719 => "001110101000011011000100",
20720 => "001111001111111011111000",
20721 => "001110111011010111100000",
20722 => "001101110010010011001110",
20723 => "001100011100011100011100",
20724 => "001011101001000100100111",
20725 => "001001111100010011100110",
20726 => "000111100010000010011010",
20727 => "000100111101101001011011",
20728 => "000011001001110111100110",
20729 => "000011110100111011011111",
20730 => "000101110101001001100000",
20731 => "000111111001100111100111",
20732 => "001010001001000110000110",
20733 => "001100100010011000010110",
20734 => "001101111101111111001100",
20735 => "001100101110110111011110",
20736 => "001000000010001001011011",
20737 => "000000101000111011000100",
20738 => "111001101010100101011110",
20739 => "110010001110111001010100",
20740 => "101000011011000001111010",
20741 => "100001111110011011001001",
20742 => "100001010000110010010100",
20743 => "100001110000100010001000",
20744 => "100001110101001011001001",
20745 => "100010011000011010000110",
20746 => "100011011011111100000110",
20747 => "100100010010101011011111",
20748 => "100101000000101100011111",
20749 => "100111001001111110001111",
20750 => "101100100011010110111110",
20751 => "110011010011001101011010",
20752 => "110111111110100000100010",
20753 => "111011100000110101111101",
20754 => "111110010101010100010000",
20755 => "111111011101101000010010",
20756 => "111111110101101001000001",
20757 => "111111110010001010111011",
20758 => "111111000000100000100110",
20759 => "111101001110110000101111",
20760 => "111011110001111010000100",
20761 => "111011110001011010110101",
20762 => "111011101111101001100111",
20763 => "111011100101100101010100",
20764 => "111011111110001111100000",
20765 => "111100011001001010110101",
20766 => "111100000111000100111010",
20767 => "111100010101101001101110",
20768 => "111111010101000011001111",
20769 => "000100010110010001001001",
20770 => "001001100110111000110110",
20771 => "001101100011010111000100",
20772 => "010000111101101111101010",
20773 => "010110010111101101100110",
20774 => "011011101011100010111111",
20775 => "011110001101000111100111",
20776 => "011110011100001100000001",
20777 => "011101110100100110110000",
20778 => "011101001110011010001011",
20779 => "011100011000010000011111",
20780 => "011011110001011111101001",
20781 => "011011000010001001111101",
20782 => "011001100110011011110110",
20783 => "010110110011011011000000",
20784 => "010001000101100101011000",
20785 => "001011001111001001001010",
20786 => "001000010010100011100110",
20787 => "000101111011100000010101",
20788 => "000000101010001100011111",
20789 => "111001001001011000101111",
20790 => "110011100000110100111000",
20791 => "110001001111101000001100",
20792 => "110001011101000100100000",
20793 => "110011010000011000110000",
20794 => "110111010110011101000000",
20795 => "111101110001110111110000",
20796 => "000010110011000110011101",
20797 => "000101111110111011101101",
20798 => "001000011001100001011101",
20799 => "001001011101001001000110",
20800 => "001010100010001001101000",
20801 => "001011100100001111111111",
20802 => "001100001001101011101100",
20803 => "001011110100011000000111",
20804 => "001010101011010000110001",
20805 => "001010010100111110110110",
20806 => "001001100101000101000000",
20807 => "001000000011100101000111",
20808 => "000110011010001111100110",
20809 => "000101010010000000100110",
20810 => "000100101011111111000100",
20811 => "000001111100001100101010",
20812 => "111011011011011101101110",
20813 => "101111100000100011101000",
20814 => "100011111001111001001011",
20815 => "100001010000011101110000",
20816 => "100010000011110001110111",
20817 => "100001010100111001010111",
20818 => "100001011100000011100001",
20819 => "100010100000010010010001",
20820 => "100011110001110001011000",
20821 => "100101001101110100100111",
20822 => "101010010011001011110010",
20823 => "110011010001111010111010",
20824 => "111011100111111010011000",
20825 => "000010011101011100101000",
20826 => "001000100011001101001010",
20827 => "001110110000101001100000",
20828 => "010010110001111010010100",
20829 => "010001101111110000110010",
20830 => "001100110111001100111100",
20831 => "000100111001111001111001",
20832 => "111100011111000110100101",
20833 => "110101110111111110011011",
20834 => "110001010011111011111000",
20835 => "101111010100101011000000",
20836 => "101110001111101001100000",
20837 => "101110100000101100101100",
20838 => "110000010111010110111010",
20839 => "110010001010000110001100",
20840 => "110101011110001010100101",
20841 => "111010011111011100010111",
20842 => "111111110111110001100010",
20843 => "000101001110001101010000",
20844 => "001010000011111000000011",
20845 => "001110010100011011100000",
20846 => "010000101010011010110110",
20847 => "010001000001011110011010",
20848 => "010010001010010101001010",
20849 => "010101011101001100111110",
20850 => "011001000110010001011110",
20851 => "011010010001010111101101",
20852 => "011001010101100111111111",
20853 => "011000010100001001000010",
20854 => "010111001110010111101010",
20855 => "010110010111100100000010",
20856 => "010101100011100010010110",
20857 => "010010101111100011111010",
20858 => "001110001110010010110010",
20859 => "001001101110000101000001",
20860 => "000101100010000010101111",
20861 => "000010000010100111111001",
20862 => "111111011101011110110000",
20863 => "111110010100101110011111",
20864 => "111111110000010110101010",
20865 => "000011001111100000100111",
20866 => "000110101010001001001000",
20867 => "001000100111001110000011",
20868 => "001001011010001000101010",
20869 => "001000011011000011110111",
20870 => "000100110000101110010010",
20871 => "111110010100111010001000",
20872 => "110101011101101101111111",
20873 => "101101011000100110000010",
20874 => "100111010000100110111011",
20875 => "100010011111110001100000",
20876 => "100001000111111010011001",
20877 => "100001100011000110101001",
20878 => "100001100011101011000011",
20879 => "100001101100010000111101",
20880 => "100001100111000010000001",
20881 => "100001111010111011100001",
20882 => "100010101011101111011001",
20883 => "100011011101100010011001",
20884 => "100100001000101100111011",
20885 => "100100011110011110001111",
20886 => "100101011010000001110011",
20887 => "100110001110110100000100",
20888 => "100110010101100110101110",
20889 => "100111000010101111100001",
20890 => "101000111000101101100000",
20891 => "101010100101011000001100",
20892 => "101011101011111110101000",
20893 => "101110111101111010111110",
20894 => "110100000010011000010001",
20895 => "111000110010000010110000",
20896 => "111110001100010100101111",
20897 => "000011110011011110010101",
20898 => "001001001011101111101101",
20899 => "001101001101110001101110",
20900 => "001110100101100100110010",
20901 => "001110101111001101000100",
20902 => "001101100000010100010000",
20903 => "001011011001000100000000",
20904 => "001010000100010101011110",
20905 => "001010000010000101100111",
20906 => "001010111101111111110011",
20907 => "001011010010001111101000",
20908 => "001100000101000100000000",
20909 => "001110101011001001110000",
20910 => "010010100010111000001100",
20911 => "010111000011100100111110",
20912 => "011010011101010010001110",
20913 => "011101000000111111000010",
20914 => "011110010101101110011101",
20915 => "011101110100101100111110",
20916 => "011100011011000001111111",
20917 => "011000000011100100110101",
20918 => "010010000100011110011000",
20919 => "001101110001010001010000",
20920 => "001010000100001100000100",
20921 => "000111000011010010011101",
20922 => "000100110010100011010010",
20923 => "000010111110011000100000",
20924 => "000010001000001110000100",
20925 => "000000001111010001010110",
20926 => "111100100110100001010001",
20927 => "111001101000010100001010",
20928 => "110111110110100001111100",
20929 => "110101011101000111000001",
20930 => "110010111111100100000010",
20931 => "110001110101011011010100",
20932 => "101111110010001100011100",
20933 => "101011100101110011010100",
20934 => "100110110011001110111110",
20935 => "100011010111110110110011",
20936 => "100011110001101001100110",
20937 => "100111100010001110001110",
20938 => "101100000010011010100110",
20939 => "110000011010100100010000",
20940 => "110011011100000000101000",
20941 => "110100011110101100001010",
20942 => "110100111011111100000011",
20943 => "110101110100101100000010",
20944 => "110111111001011101000010",
20945 => "111011000001000110100101",
20946 => "111110000010010101111011",
20947 => "000000110110010010110000",
20948 => "000100000101101010011110",
20949 => "000111100010001001111010",
20950 => "001001100010010111011100",
20951 => "001010001001111010001110",
20952 => "001011001011010000000101",
20953 => "001100110111001110001100",
20954 => "001111001111101111111000",
20955 => "010000101110011101111010",
20956 => "001111010100111111111100",
20957 => "001100011111110101100000",
20958 => "001001110101111001100010",
20959 => "001000001011011010011011",
20960 => "000111000000100000100000",
20961 => "000110000000010011011100",
20962 => "000111000010100101101111",
20963 => "001001001110011001110100",
20964 => "001011001010110111001000",
20965 => "001100110111100100010000",
20966 => "001101001011111111101000",
20967 => "001100010111111001101100",
20968 => "001010110111011001111100",
20969 => "001010010001110100001110",
20970 => "001100011010011010111110",
20971 => "001111001011001000110100",
20972 => "010001100100001000011100",
20973 => "010011100111010010011100",
20974 => "010011000101001110010100",
20975 => "001110110110111101010100",
20976 => "001000100100100000100010",
20977 => "000010000011011101101000",
20978 => "111011000001110111011001",
20979 => "110011110000110111110000",
20980 => "101101011101000100110110",
20981 => "101000011110011101110010",
20982 => "100110010000110001110100",
20983 => "100111000101101000010011",
20984 => "101001011100011110011110",
20985 => "101101010010101110110110",
20986 => "110011011011100001000010",
20987 => "111011011111000010100001",
20988 => "000010111111111100011011",
20989 => "001000000100101110011001",
20990 => "001011001001001110111010",
20991 => "001100110000111010000100",
20992 => "001101101011000011001010",
20993 => "001110111010010101110010",
20994 => "010000011000001011001110",
20995 => "010001101010110010011000",
20996 => "010011001010101000110100",
20997 => "010100011111001000111100",
20998 => "010100010001111011000010",
20999 => "010010010001010010010010",
21000 => "001111000110001111111000",
21001 => "001100000110011011001010",
21002 => "001010011110001100001000",
21003 => "001001010111111100111100",
21004 => "001000001110111101011111",
21005 => "000111110010001000101100",
21006 => "000111100110100000100100",
21007 => "000110110010011101000010",
21008 => "000101011111000000110011",
21009 => "000100100001101001011101",
21010 => "000100101010110110001001",
21011 => "000100110111011101001001",
21012 => "000011000101011101000110",
21013 => "111111111011001110010001",
21014 => "111100110101100010010100",
21015 => "111001011101001000100101",
21016 => "110111001110111101010000",
21017 => "111000010000011111101100",
21018 => "111010001010110000110110",
21019 => "111001111111000111101000",
21020 => "111000001101111011001001",
21021 => "110110011010000010100011",
21022 => "110101011011111111100010",
21023 => "110011111011110001110010",
21024 => "101111110101110001010100",
21025 => "101010111111001111010010",
21026 => "100111010010000100011101",
21027 => "100011111111011001100111",
21028 => "100010000001010110001100",
21029 => "100001111101111010010001",
21030 => "100010100111000100001100",
21031 => "100100000000000000110101",
21032 => "100110100011101110111101",
21033 => "101001110111000000001100",
21034 => "101100100001011111101110",
21035 => "101101110100101101001100",
21036 => "101111100000110101011000",
21037 => "110010000011011010111110",
21038 => "110011100010011001111010",
21039 => "110011111011011000000100",
21040 => "110101000000011100001000",
21041 => "110111111101111000011000",
21042 => "111100110110010001110001",
21043 => "000001110110010011101100",
21044 => "000101001110111110001100",
21045 => "001000101101101111100110",
21046 => "001101101001100011011000",
21047 => "010001100111110001110010",
21048 => "010011010111110101001100",
21049 => "010011011100111100011100",
21050 => "010010001110011010000100",
21051 => "010001000010011001110010",
21052 => "001111001001010101001000",
21053 => "001010111111001101110110",
21054 => "000111001010111101101101",
21055 => "000110101001001001100001",
21056 => "001001000001001010011011",
21057 => "001100110010111000110010",
21058 => "010001100110110011000100",
21059 => "010110101000111001111010",
21060 => "011001100101011111100101",
21061 => "011010100001001101100010",
21062 => "011010110101100010011011",
21063 => "011010100011110110111001",
21064 => "011010001000010000101110",
21065 => "011000101111111000101111",
21066 => "010100110001111000010010",
21067 => "010000000110011101001110",
21068 => "001101100000001111001100",
21069 => "001010100101011000101010",
21070 => "000100111110110011100010",
21071 => "111111001100010110010010",
21072 => "111001011000001100001100",
21073 => "110100000100010101000111",
21074 => "101111110101100111110100",
21075 => "101000011101100101111000",
21076 => "100001110110101000000011",
21077 => "100001001110001010101101",
21078 => "100001100100111000101101",
21079 => "100001011001110111001111",
21080 => "100001100001001010110111",
21081 => "100001011110101101110101",
21082 => "100010100110110110001011",
21083 => "100011101000000001100000",
21084 => "100100100001110100101111",
21085 => "100110011111111100000011",
21086 => "101000010010010111001000",
21087 => "101001001101100001011100",
21088 => "101010011111011111001000",
21089 => "101101001111111100110000",
21090 => "101111110111100000101010",
21091 => "110010010011101110110000",
21092 => "110101010100011011101011",
21093 => "110111000000100011011000",
21094 => "110111101100011011001111",
21095 => "111000000101000010111110",
21096 => "111000101100110110111010",
21097 => "111010100110101111110101",
21098 => "111100110111110111111001",
21099 => "111110101010010100100000",
21100 => "111110101011101001000000",
21101 => "111101101101001110110111",
21102 => "111101111011000010001011",
21103 => "111110110001110011111011",
21104 => "000000100101011110010001",
21105 => "000011111000010010000100",
21106 => "001000100110000000111011",
21107 => "001110010000010000000100",
21108 => "010011100011011000011010",
21109 => "011000010000110010100110",
21110 => "011011001010001110100111",
21111 => "011100011111010101000000",
21112 => "011101110100000010000111",
21113 => "011110011111101010001001",
21114 => "011110101101001110110101",
21115 => "011110100000000011111111",
21116 => "011110001100110000011011",
21117 => "011110000110110011010101",
21118 => "011100011110101000110101",
21119 => "011001000100011001000110",
21120 => "010100110110111100000110",
21121 => "010001101101110011100100",
21122 => "010000111010000000100000",
21123 => "010000011111100101101110",
21124 => "001110110001010010000110",
21125 => "001011101011001101010011",
21126 => "001000100110100010111000",
21127 => "000110011000010010101000",
21128 => "000100011011100110101011",
21129 => "000011100100011111001011",
21130 => "000100000101101011110110",
21131 => "000101011110111011100100",
21132 => "000111100011101110010010",
21133 => "001000110000100001011010",
21134 => "000111100101001111010110",
21135 => "000100110010001110000101",
21136 => "000010100101000001000010",
21137 => "000010001101011000110010",
21138 => "000011010010110100100000",
21139 => "000100001010101010000110",
21140 => "000011110000100000010011",
21141 => "000010000110010111101110",
21142 => "111101100000111011100010",
21143 => "110101110100000010100001",
21144 => "101101010000111010100010",
21145 => "100101100100111110100010",
21146 => "100001100010010001000101",
21147 => "100001010101110100111101",
21148 => "100001101001000010111101",
21149 => "100001011101101101100111",
21150 => "100001100010011110110011",
21151 => "100010000010000000110101",
21152 => "100011011110110100101000",
21153 => "100111010101101111001001",
21154 => "101110000010100111110100",
21155 => "110110001001110000110000",
21156 => "111110010010101100000011",
21157 => "000100011000001011110010",
21158 => "000110001100101011100100",
21159 => "000100101001000110101001",
21160 => "000010010000011111001110",
21161 => "111111100001101101101001",
21162 => "111100011011110100101100",
21163 => "111010010111101100101011",
21164 => "111000111100110100011000",
21165 => "110111010000000011100001",
21166 => "110110001001100100001001",
21167 => "110101101001000100000000",
21168 => "110101010111101111000010",
21169 => "110101100001010000001000",
21170 => "110101111011011100111110",
21171 => "110110011011101111001111",
21172 => "110111001100100001001010",
21173 => "111000111000011000111011",
21174 => "111011101001001100010110",
21175 => "111111000100111001110101",
21176 => "000010110001100000010101",
21177 => "000110100111011100011010",
21178 => "001010110010110110101000",
21179 => "001110110111011111101000",
21180 => "010010101101010001011010",
21181 => "010110010101001001110000",
21182 => "011001101000100011100111",
21183 => "011100001000000110110101",
21184 => "011011111101100011111011",
21185 => "011001111110100000110011",
21186 => "010111101101011011010110",
21187 => "010011011011000001110110",
21188 => "001101001110010110100000",
21189 => "000110110011000011101001",
21190 => "000001101011000100111110",
21191 => "111111100010111110001100",
21192 => "111111001010011111101000",
21193 => "111111000110011010011110",
21194 => "000000100000010001010000",
21195 => "000100001000001100001110",
21196 => "001000001001100110010010",
21197 => "001001110110111100010100",
21198 => "001001111010000100010111",
21199 => "001010101100101000111110",
21200 => "001100011000100100010110",
21201 => "001101010100110111110010",
21202 => "001100010001000101010100",
21203 => "001010100100111101100010",
21204 => "001001100011101111000000",
21205 => "000111110111000001100100",
21206 => "000101000101010101110010",
21207 => "000011010000100011011001",
21208 => "000011111101001001110010",
21209 => "000101100101110000011101",
21210 => "000101111001100101010011",
21211 => "000101010110101011000000",
21212 => "000011101100010100110010",
21213 => "111111010001011111110011",
21214 => "111001000001111110011010",
21215 => "110010101101111110110010",
21216 => "101100100011011111011010",
21217 => "100111001001111110111001",
21218 => "100011100101111000111000",
21219 => "100001110010000111101111",
21220 => "100001010111010110111000",
21221 => "100001111011010100111010",
21222 => "100010110111111011011101",
21223 => "100100000111010001111011",
21224 => "100101010001011010110111",
21225 => "101000011011101011001110",
21226 => "110000011100000110101000",
21227 => "111001100101000010000010",
21228 => "111111101111010101011011",
21229 => "000011010110000010100101",
21230 => "000100010000110111100010",
21231 => "000100000011000001110010",
21232 => "000100011111111110111110",
21233 => "000100001011001011001100",
21234 => "000010110000010110101010",
21235 => "000000110111110110000000",
21236 => "111110100111011011010110",
21237 => "111011101111100111110010",
21238 => "110111101100011101100111",
21239 => "110100001000101010000000",
21240 => "110011101101111011011110",
21241 => "110111000000111000111100",
21242 => "111011101110101111100101",
21243 => "111110100110001110010010",
21244 => "111111101011111011111100",
21245 => "000001001010110000111111",
21246 => "000011001001001011010111",
21247 => "000100001110110100110100",
21248 => "000100110101001000100100",
21249 => "000111010011100110110111",
21250 => "001011011001110100101110",
21251 => "001110011010000000011110",
21252 => "010000010000110010110100",
21253 => "010001100111001000111100",
21254 => "010000010000001100001100",
21255 => "001011010101111011010010",
21256 => "000110011011001110110010",
21257 => "000100110001000011110101",
21258 => "000101001000000100010110",
21259 => "000100100011000110000111",
21260 => "000010100111110011010000",
21261 => "000000101001001101101011",
21262 => "111111101011111001010110",
21263 => "111111100010100111110010",
21264 => "111110100100110000001000",
21265 => "111110000010100010010011",
21266 => "000001000101011001101010",
21267 => "000110010001000111011110",
21268 => "001010010111111100101110",
21269 => "001100100000100100001010",
21270 => "001101000000110101011000",
21271 => "001101000110010011011110",
21272 => "001101000100101101111000",
21273 => "001100111010010100001110",
21274 => "001101101000110011000010",
21275 => "001110000011111010000110",
21276 => "001011110110000110111111",
21277 => "001000000100111100100110",
21278 => "000101001100001010101011",
21279 => "000011011001000111000011",
21280 => "000001011101100111101001",
21281 => "111111001110100110001111",
21282 => "111110101101101101100011",
21283 => "000000100011001000110000",
21284 => "000001110111101001000111",
21285 => "000000001011101101111000",
21286 => "111011010111100100111000",
21287 => "110101101001000101011111",
21288 => "110000100111110000010010",
21289 => "101011111010101000010000",
21290 => "101001100011001000111100",
21291 => "101010100001001110010000",
21292 => "101100111111011101000110",
21293 => "110001010000011110110110",
21294 => "110110011010000000111111",
21295 => "111011000100110100111000",
21296 => "000000100110001110011010",
21297 => "000110101110101001010111",
21298 => "001011100111110010111110",
21299 => "001110000111100001001000",
21300 => "001110010111100000010010",
21301 => "001100011111001001011100",
21302 => "000111110010011010100010",
21303 => "000001110000110000111110",
21304 => "111100010101000011111001",
21305 => "110110011011011001111001",
21306 => "101110010111100100100010",
21307 => "100110010111110101110101",
21308 => "100010110001010101001001",
21309 => "100011001111010101000011",
21310 => "100100100101111010010100",
21311 => "100101011111101000010111",
21312 => "100110011011101010110010",
21313 => "100111101001111101101000",
21314 => "101000100101000110100000",
21315 => "101011111001001101000000",
21316 => "110011001101110000100100",
21317 => "111010101100111001000011",
21318 => "000001010101011111101110",
21319 => "001001000011111001100011",
21320 => "010001010001011110001100",
21321 => "010111100011110000001000",
21322 => "011010101001000000110011",
21323 => "011011111011100100111101",
21324 => "011011010100000101100101",
21325 => "010111001010101101111110",
21326 => "010000111101001001100000",
21327 => "001011101100110000011011",
21328 => "001000010101101111111010",
21329 => "000101010101000110101011",
21330 => "000010001000111000100000",
21331 => "111111101111101011110011",
21332 => "111110111000000100101100",
21333 => "111111101011010011001111",
21334 => "000000111001101101100001",
21335 => "000010111001110010011001",
21336 => "000110111100011111110011",
21337 => "001100010001010100100100",
21338 => "010001110101001010100010",
21339 => "010110001011111001010010",
21340 => "011001010111001111110101",
21341 => "011011011100111101100111",
21342 => "011010110010110001000110",
21343 => "011001001100001111101101",
21344 => "011000100010101100110111",
21345 => "010111101111101111000000",
21346 => "010110101110001010101010",
21347 => "010101111101111100100000",
21348 => "010101001110101010111000",
21349 => "010001011110100010010100",
21350 => "001000001101101000010101",
21351 => "111101001010111011111001",
21352 => "110100011101101001000000",
21353 => "101101101101010111110000",
21354 => "101000011100000011010110",
21355 => "100101100011010111110101",
21356 => "100011110010000101011101",
21357 => "100010000110010110010001",
21358 => "100010011101100010001101",
21359 => "100100000110101110111011",
21360 => "100101001011110011000111",
21361 => "100111001111000001111101",
21362 => "101001010011100111110010",
21363 => "101000010101101011011100",
21364 => "100101111100000001100110",
21365 => "100101100100110100101111",
21366 => "100110010101110011011111",
21367 => "100110001110111111000110",
21368 => "100110011010011100110000",
21369 => "100111000010011001110111",
21370 => "100111010011010011011001",
21371 => "101000110111001110000100",
21372 => "101100011001111010110100",
21373 => "110000001111011111110110",
21374 => "110100011101110001010101",
21375 => "111010000110100100010001",
21376 => "111110101111100010101010",
21377 => "000000100001010000000011",
21378 => "000001011111100100010010",
21379 => "000010010110010001001111",
21380 => "000010000011001100101111",
21381 => "000000100000011000100010",
21382 => "111111001101111111010010",
21383 => "000001010101001011100001",
21384 => "000110111000101011110001",
21385 => "001101000011110101101010",
21386 => "010010111001100010000110",
21387 => "011000000100011110011100",
21388 => "011011110110101110110001",
21389 => "011101110101000000111010",
21390 => "011110010010110000110011",
21391 => "011110011101101010000010",
21392 => "011110010111001000110100",
21393 => "011101011010110000000010",
21394 => "011100011010100011101000",
21395 => "011011111011111010010011",
21396 => "011011100101011010101011",
21397 => "011001011101101110111111",
21398 => "010011001010010111000110",
21399 => "001011011011100011100000",
21400 => "000111001110001110100001",
21401 => "000101010101001000100100",
21402 => "000011010011001100110101",
21403 => "000010001111010011000011",
21404 => "000010011000101110110010",
21405 => "000010000101111010111001",
21406 => "000000010001110110111111",
21407 => "111110100111101001000011",
21408 => "111111011111010101110001",
21409 => "000001110110101000110010",
21410 => "000010111000010111011101",
21411 => "000001100011001101100110",
21412 => "111111100010001001001110",
21413 => "111101100000000000001010",
21414 => "111010001001111011001001",
21415 => "110110110100101100011110",
21416 => "110101001001101111011011",
21417 => "110011110101011001101110",
21418 => "110001101110101010010010",
21419 => "101111010010111111111010",
21420 => "101100101011010101010100",
21421 => "101000100001000011100100",
21422 => "100011110001010110011010",
21423 => "100001101101010110110011",
21424 => "100001110111001010101111",
21425 => "100010010000111010010001",
21426 => "100011001000110101001011",
21427 => "100100000100000101101101",
21428 => "100101001101110001011000",
21429 => "101001001110100001011110",
21430 => "110000001011011010011110",
21431 => "110111011000000011100110",
21432 => "111110010111101110101101",
21433 => "000100110111100101001111",
21434 => "001010010101111101100010",
21435 => "001111001110101000100110",
21436 => "010001111011001011110010",
21437 => "010010101111110001111100",
21438 => "010011111111111000110010",
21439 => "010100011110001111100000",
21440 => "010011011111000100011100",
21441 => "010011001001101101010010",
21442 => "010100101000101100100010",
21443 => "010110000010001100011010",
21444 => "010100110000000110100010",
21445 => "010001011101110010001010",
21446 => "001101110010000011111110",
21447 => "001010001111100010110001",
21448 => "000110100010111100100100",
21449 => "000001111000110010101101",
21450 => "111101011011100110011110",
21451 => "111010001001100010000100",
21452 => "111000001011010001001101",
21453 => "111001001101110000001011",
21454 => "111101000000011101001101",
21455 => "000000010101111000001101",
21456 => "000010101010001011110110",
21457 => "000111001000110010110011",
21458 => "001101011110001101011110",
21459 => "010001101101000001010010",
21460 => "010011110110010011110000",
21461 => "010101011101101110010100",
21462 => "010101110111101100110000",
21463 => "010100110011101000011110",
21464 => "010010001001110111111100",
21465 => "001101010010110001000100",
21466 => "000110101010110000000101",
21467 => "000000001011000000000001",
21468 => "111010101001101011010000",
21469 => "110101010010000111100100",
21470 => "101111001101100110110000",
21471 => "100111111111101010111001",
21472 => "100010100100100110011011",
21473 => "100001100010010000100111",
21474 => "100001011011111010101001",
21475 => "100000110011000111000101",
21476 => "100010011010100011101000",
21477 => "100111001011101010100100",
21478 => "101111111111010111110000",
21479 => "111100101111011111110101",
21480 => "001001111001011010000111",
21481 => "010101000001110010101110",
21482 => "011100001011110000111011",
21483 => "011101001100000011100111",
21484 => "011011001110101010010101",
21485 => "011001111100001011110001",
21486 => "011000011001001101111111",
21487 => "010111000001011100111110",
21488 => "010100101001001011010100",
21489 => "001110000111000000101110",
21490 => "000110011001101000100110",
21491 => "000000001101000001000010",
21492 => "111001110101101110011001",
21493 => "110100001111101010100110",
21494 => "110001000100001100101110",
21495 => "101111101110011111101110",
21496 => "101111111111010100011110",
21497 => "110001100001100101110010",
21498 => "110011000111001001010100",
21499 => "110100000110100110000000",
21500 => "110100101101010100111010",
21501 => "110101100100101001110011",
21502 => "110111101110011010000010",
21503 => "111011001000101111110101",
21504 => "111110010001110101011010",
21505 => "111111110001111111011101",
21506 => "111111010101011010100101",
21507 => "111100111001011001100110",
21508 => "111000001001110000010010",
21509 => "110011000111100011101010",
21510 => "110001100010000111100000",
21511 => "110011000100011110100010",
21512 => "110100010100101111001000",
21513 => "110100011001110111111001",
21514 => "110011100100001110101100",
21515 => "110000100011011000010010",
21516 => "101011111001101100010010",
21517 => "101000001100101011011010",
21518 => "100110110000101101100111",
21519 => "101000010010011101001010",
21520 => "101100010011011011010010",
21521 => "110001110010010001111010",
21522 => "111000110000001100001101",
21523 => "111111110101011000010111",
21524 => "000110011010000010100011",
21525 => "001100110110010100000100",
21526 => "010010000010110011100000",
21527 => "010110010010000110100110",
21528 => "011001000101010011100001",
21529 => "011000100100000101001110",
21530 => "010101100110011110000010",
21531 => "010001100100101101111010",
21532 => "001100110110000001001100",
21533 => "000111100111010111111111",
21534 => "000010110110101100100000",
21535 => "000000110101000010010000",
21536 => "000010010000011110001100",
21537 => "000101101000001011111110",
21538 => "001001010110101110010010",
21539 => "001101001010110110101100",
21540 => "010000011010000110011010",
21541 => "010000011001111111001010",
21542 => "001100110000110100100110",
21543 => "001001000110100000111110",
21544 => "001000000000111101110100",
21545 => "001000011011001010110001",
21546 => "001000111011101111010110",
21547 => "001001010101010011100100",
21548 => "001001000000110001101110",
21549 => "001000001110111111100111",
21550 => "000111011011010110111110",
21551 => "000110111010000000111011",
21552 => "001000001000110110101100",
21553 => "001010100101100001001100",
21554 => "001100100001110011101010",
21555 => "001100111111000001001000",
21556 => "001011001110001110100011",
21557 => "000111001111001111001000",
21558 => "000000011001111110001010",
21559 => "110111110001011011010110",
21560 => "101110111011010101011100",
21561 => "100110011001100101000111",
21562 => "100001111000011111010100",
21563 => "100001101010010100111111",
21564 => "100001110000001000100111",
21565 => "100010000001101010101101",
21566 => "100010100101010010011011",
21567 => "100011010011001101110011",
21568 => "100100011011111111111101",
21569 => "100101000110011100000001",
21570 => "101000100000110110101110",
21571 => "110001001110100100111100",
21572 => "111010110110100011101111",
21573 => "000001011100110001011111",
21574 => "000100101111110011000111",
21575 => "000101000011011100111001",
21576 => "000011110100011011001110",
21577 => "000001110100101111010101",
21578 => "111110011000110111100100",
21579 => "111011100100000101000111",
21580 => "111010011001101100110011",
21581 => "111000111011111111100110",
21582 => "111000000111101101011111",
21583 => "111000001011011111110110",
21584 => "110111011110010011000100",
21585 => "110111100011100111101100",
21586 => "111001100101100010000001",
21587 => "111011110101100011000010",
21588 => "111011101000001110000101",
21589 => "111001000001001001101100",
21590 => "111000000010110010011101",
21591 => "111010010111000001010100",
21592 => "111101100001010001110110",
21593 => "111111101011000010000000",
21594 => "000010111000111101100110",
21595 => "001001111001011001010111",
21596 => "010001101010000001010000",
21597 => "010110001011101011011100",
21598 => "011000001111011000010011",
21599 => "011001101101100010010001",
21600 => "011010110111011010110000",
21601 => "011001111001111010001110",
21602 => "010101101000001001110010",
21603 => "001111110101100001001000",
21604 => "001011000001100000100001",
21605 => "001000011001101111111010",
21606 => "000111000000001101001000",
21607 => "000101011010101011100111",
21608 => "000100011010010011111100",
21609 => "000101001101001000101000",
21610 => "000110101010000111100000",
21611 => "000110100110111111011011",
21612 => "000110011010101101101001",
21613 => "001000110111011011100010",
21614 => "001100010101001100100110",
21615 => "001110000001100001100100",
21616 => "001110011010111011100000",
21617 => "001111000011011101101010",
21618 => "010000001100101111010000",
21619 => "010001010000010011111110",
21620 => "010001110100001011011110",
21621 => "010001110011111100001000",
21622 => "010001111010100011110010",
21623 => "010011000010110101000000",
21624 => "010100001110011000010010",
21625 => "010011011001010111100000",
21626 => "010000000111011100100100",
21627 => "001100000001001111100100",
21628 => "001000100011001010101111",
21629 => "000101010001101001010011",
21630 => "000001111101110011110100",
21631 => "111111101010100110001001",
21632 => "111110110010101100000100",
21633 => "111101110010000101111100",
21634 => "111010000101111010100011",
21635 => "110011101011101100000000",
21636 => "101100101101111011100110",
21637 => "100110110100101101101001",
21638 => "100011010001000001011001",
21639 => "100001110100010100111101",
21640 => "100010010110001101101001",
21641 => "100110001100111101111011",
21642 => "101011110100111110111010",
21643 => "110001000001001100011000",
21644 => "110101111101111101100000",
21645 => "111010010000101000010100",
21646 => "111101110000000110010100",
21647 => "000000100110000111001001",
21648 => "000010001111000011110001",
21649 => "000001110011001001111010",
21650 => "111101011111110000000001",
21651 => "110110010000011000000101",
21652 => "101111100010100001001110",
21653 => "101010010100010000110000",
21654 => "100111001000001111000010",
21655 => "100111110101110010001111",
21656 => "101100011001011011100000",
21657 => "110010011010011010111100",
21658 => "110111100010111010011010",
21659 => "111010001111101111001000",
21660 => "111010011001010011001101",
21661 => "111010010011011000001000",
21662 => "111100100010010010001101",
21663 => "000000110101001101110010",
21664 => "000100010111100011000111",
21665 => "000110111000000010100111",
21666 => "001011011101101001011011",
21667 => "010001111000011000011110",
21668 => "010111111010010111100100",
21669 => "011100010010111000011010",
21670 => "011101000110110011110001",
21671 => "011011100101101111100100",
21672 => "011010011010000101000111",
21673 => "011001101010111111100001",
21674 => "011001000001011000011110",
21675 => "011000010110010000000111",
21676 => "010111110101000111001010",
21677 => "010100101010011000000100",
21678 => "001100111001110010001000",
21679 => "000101010011101000010001",
21680 => "111111111110011001000001",
21681 => "111011101000100001000111",
21682 => "111001000011001110001100",
21683 => "110111101110111110110000",
21684 => "111000001010001101011110",
21685 => "111010101001110100010101",
21686 => "111101000000000110000000",
21687 => "111111101100111101001000",
21688 => "000100001100101010101000",
21689 => "001001100001001101000110",
21690 => "001110011011110100101110",
21691 => "010001010000011110100110",
21692 => "001111101101100011110110",
21693 => "001001011001100011011101",
21694 => "000000011000100010001101",
21695 => "111000000110110110001011",
21696 => "110001101111000100000010",
21697 => "101010010100111001100100",
21698 => "100011011001000011000010",
21699 => "100001100001010011011101",
21700 => "100001101111100000110011",
21701 => "100001010100110111010001",
21702 => "100001100000010111110011",
21703 => "100001011100001101010101",
21704 => "100001110011111001111011",
21705 => "100010101101000110010011",
21706 => "100011010100110001100000",
21707 => "100101101101110000100101",
21708 => "101000110010101100010110",
21709 => "101010001110110101101010",
21710 => "101100000111100111010100",
21711 => "110000000001000001100110",
21712 => "110011111110000111011010",
21713 => "110111101001000111001100",
21714 => "111101000111010101101000",
21715 => "000010110010101111010101",
21716 => "000110101010001001001000",
21717 => "001001101111000000100010",
21718 => "001011100110101000010110",
21719 => "001100101110011010100100",
21720 => "001110000010110000100000",
21721 => "001110001100111011100100",
21722 => "001101000010010010010000",
21723 => "001010111101010111000011",
21724 => "001000010010011011101101",
21725 => "000101010110110100111101",
21726 => "000001100100011000000011",
21727 => "111101101011100111001101",
21728 => "111011100111101000001000",
21729 => "111100010111011111100010",
21730 => "111110100011101111000110",
21731 => "111111110100000110000010",
21732 => "000000100011111010100011",
21733 => "000010001010000100110100",
21734 => "000011110011001110110010",
21735 => "000101000010101100000011",
21736 => "000111010100010100100000",
21737 => "001010001000110011000000",
21738 => "001010111100001011000000",
21739 => "001001101011110110011001",
21740 => "000111010000001000001100",
21741 => "000011111000001011110011",
21742 => "000000001000011010001111",
21743 => "111011110001101101010010",
21744 => "110111100011101110101010",
21745 => "110100011000000100011101",
21746 => "110010000000110001111000",
21747 => "110000100010110011010110",
21748 => "101111001100100001111000",
21749 => "101110110010111010100000",
21750 => "110000101000000011010110",
21751 => "110010110111011011010100",
21752 => "110100101100111001011100",
21753 => "110110011110111100110001",
21754 => "111001000001001010100010",
21755 => "111101011111001011111010",
21756 => "000010000001110111000100",
21757 => "000101100010001110101110",
21758 => "001001001011110010101001",
21759 => "001100100010000011100000",
21760 => "001110101110101100111110",
21761 => "001111010100010001110000",
21762 => "001110001101001110101000",
21763 => "001011110110010101100010",
21764 => "001001000000000010110011",
21765 => "000111100011000100001100",
21766 => "000111110001010110111000",
21767 => "000111101110100110001100",
21768 => "000111011101111110011001",
21769 => "001000001000111100010001",
21770 => "001000110111011010111010",
21771 => "001000110100010000110011",
21772 => "001001000000001110100000",
21773 => "001010010001111110001000",
21774 => "001100100011101110011010",
21775 => "001111000000000000110010",
21776 => "010000010010110111000010",
21777 => "001111111101111110110000",
21778 => "001110011010010000110110",
21779 => "001100011110001101100010",
21780 => "001001111010101011111111",
21781 => "000110011101110111110111",
21782 => "000100111101100000001111",
21783 => "000101110010010000011100",
21784 => "000110001110000011111100",
21785 => "000110110111111100101111",
21786 => "000111001111111001010101",
21787 => "000101101100101011010110",
21788 => "000011110100111111101001",
21789 => "000001101111111011001100",
21790 => "111110011111011010100011",
21791 => "111010011111000110011101",
21792 => "110101011110110000110001",
21793 => "101111000001100011000100",
21794 => "101000010011101001011000",
21795 => "100100100011010100001001",
21796 => "100100100000101111101101",
21797 => "100101111110001001000000",
21798 => "101000111101101010101110",
21799 => "101100111110101101111010",
21800 => "101111101101100010111000",
21801 => "110000110000110101100110",
21802 => "110000011110001011010000",
21803 => "110000000010001111101110",
21804 => "110001101011110001111110",
21805 => "110101001100110100000110",
21806 => "111000110000010011110010",
21807 => "111101001111010110010101",
21808 => "000100100001000101111001",
21809 => "001100101101111001110100",
21810 => "010011000011100100010110",
21811 => "010111111110001001001000",
21812 => "011100001000110110000010",
21813 => "011101111011001100010111",
21814 => "011101000110110101100001",
21815 => "011011111010110110011101",
21816 => "011011000001011010010001",
21817 => "011010010001100010011100",
21818 => "011000011100101101111001",
21819 => "010011010000011011110000",
21820 => "001101110011110101000110",
21821 => "001011010011101111101011",
21822 => "001001111000001110110000",
21823 => "001001111111000101010001",
21824 => "001011100011011100101100",
21825 => "001011110111111010100101",
21826 => "001011001011011101110100",
21827 => "001010001001000000111111",
21828 => "001001000001010011010111",
21829 => "001000111011100011101001",
21830 => "001010001001011100010000",
21831 => "001100010011010110010110",
21832 => "001110110110010001010000",
21833 => "010001100001100011010100",
21834 => "010010001010101101100000",
21835 => "001101010011010100001010",
21836 => "000100110110010101111111",
21837 => "111110000111100110111001",
21838 => "111001101001110110010110",
21839 => "110100100000111100011111",
21840 => "101110000100111011110000",
21841 => "100111101110010111110101",
21842 => "100011001010010101110111",
21843 => "100001100111010001000011",
21844 => "100001100011011011000101",
21845 => "100001100100001111111101",
21846 => "100010001101000111100001",
21847 => "100010111001011110010100",
21848 => "100100010001010111010111",
21849 => "100111111000000111111101",
21850 => "101011111100101111100000",
21851 => "101110101110101100111010",
21852 => "110001110110000111010000",
21853 => "110110110100111010100111",
21854 => "111100001001001101100100",
21855 => "000000011010100001000000",
21856 => "000100001101100111101000",
21857 => "000110111111101000111101",
21858 => "000111101001101001001100",
21859 => "000110001110000101110100",
21860 => "000011010111001000001000",
21861 => "000000001001110111110001",
21862 => "111101101011100000010100",
21863 => "111100010101101000011101",
21864 => "111010110111101111001010",
21865 => "111001100100011101001010",
21866 => "111011011001110010011111",
21867 => "111111111110110100111000",
21868 => "000100010101001001001101",
21869 => "000110110101101110000001",
21870 => "001000001000101111100000",
21871 => "001010101100110101100111",
21872 => "001101010000001101010100",
21873 => "001100111001111101011110",
21874 => "001011001010001111000101",
21875 => "001001000111101001101011",
21876 => "000110000100100000110111",
21877 => "000010100100001011010110",
21878 => "000000000110110101000001",
21879 => "000000001011110111111100",
21880 => "000010010110111101011011",
21881 => "000101000000100100111101",
21882 => "000111010010100101010100",
21883 => "001001001000000111111110",
21884 => "001011000100101111101100",
21885 => "001100101000100001110000",
21886 => "001011111001111110011010",
21887 => "001000100100000010110110",
21888 => "000100011001111110001110",
21889 => "111111110011111010011101",
21890 => "111010001100011000111110",
21891 => "110100101000010100010011",
21892 => "101111110010111011110000",
21893 => "101100110001110111100000",
21894 => "101101001100010011000010",
21895 => "110000001011101010110000",
21896 => "110100001100010000111000",
21897 => "110111000111010111100000",
21898 => "111000100011001100100100",
21899 => "111011010011011000011101",
21900 => "111110010111011100011111",
21901 => "111111000011101001011001",
21902 => "111110101001101100010110",
21903 => "111110010111001011111001",
21904 => "111101001011011000100000",
21905 => "111001101100010101110011",
21906 => "110100111111000101000100",
21907 => "110001111011110010110110",
21908 => "110000111110101011011010",
21909 => "110000111100010101110010",
21910 => "110001011111110011111000",
21911 => "110011001001001110100010",
21912 => "110101101010111110101100",
21913 => "110111011011000011100010",
21914 => "110111101100011010011111",
21915 => "110111110000100011101110",
21916 => "111001011010000000011100",
21917 => "111100110110110001111110",
21918 => "000000001010010010011011",
21919 => "000001111011111000000101",
21920 => "000011000100001010100111",
21921 => "000100100111100011000110",
21922 => "000101100101111010011010",
21923 => "000101100100101110100110",
21924 => "000110010101001011001100",
21925 => "000111111100001001111000",
21926 => "001001000000001011101000",
21927 => "001000110110110011111010",
21928 => "000111101000100100111100",
21929 => "000110101011100001011100",
21930 => "000101111001100111011000",
21931 => "000100001110001011011111",
21932 => "000011000010000000110000",
21933 => "000011011111101000110110",
21934 => "000011100111110001010001",
21935 => "000000111010000001101111",
21936 => "111100011111000001001010",
21937 => "111000110000001100001000",
21938 => "110110001001100100001011",
21939 => "110101111000100110011010",
21940 => "110111110011000000101010",
21941 => "111010110100111111111100",
21942 => "000000100001101110100100",
21943 => "000110101001110101011001",
21944 => "001001100110100101111111",
21945 => "001011011010111110011000",
21946 => "001101101100001101110010",
21947 => "001111011100101010101010",
21948 => "010000010110111001111110",
21949 => "010000100110011101011100",
21950 => "010001001110010111110100",
21951 => "010011000001010001001010",
21952 => "010101001000101001000110",
21953 => "010110010100100111000110",
21954 => "010110101010010111110110",
21955 => "010110111100110011110110",
21956 => "010111101000010101001000",
21957 => "011000011000110001110000",
21958 => "011000001000010011111101",
21959 => "010110110100110110001100",
21960 => "010100100001011111000010",
21961 => "010000111001011101000110",
21962 => "001100011111000100110010",
21963 => "000110010001110101000101",
21964 => "111110000101000000011001",
21965 => "110110010110011110000111",
21966 => "110000111011111110000110",
21967 => "101110101011100001111000",
21968 => "101110011011011000011000",
21969 => "101110101000001010000110",
21970 => "101111100001111111110100",
21971 => "110001010111000110110000",
21972 => "110100000001010001100000",
21973 => "110110011000101101011111",
21974 => "111000000000110100010101",
21975 => "111010000000100011110110",
21976 => "111011100110110001110110",
21977 => "111010110011101000100000",
21978 => "110110101100111000001010",
21979 => "110001100011110111010100",
21980 => "101111000000000011010000",
21981 => "101110110110000110111110",
21982 => "101111000010000000000000",
21983 => "101110111111101001001110",
21984 => "101111001100101111000010",
21985 => "101111011110111001110000",
21986 => "101111111011011110010010",
21987 => "110001111010111011101100",
21988 => "110100000011000011000100",
21989 => "110100000010000100101001",
21990 => "110011011110010110110010",
21991 => "110100000101010011101110",
21992 => "110101010001101111000010",
21993 => "110101111110110111110010",
21994 => "110110100100100101111101",
21995 => "111000110001011000000010",
21996 => "111101001100110100000101",
21997 => "000010110111111100111000",
21998 => "001000010010000000101000",
21999 => "001100110100011000111100",
22000 => "010000110011010000011110",
22001 => "010100000100101100110100",
22002 => "010101011010110111000110",
22003 => "010011011110010101001010",
22004 => "001111100001011100011100",
22005 => "001011111001110000000011",
22006 => "001000010111111011000010",
22007 => "000100010111101111110001",
22008 => "000001000110010001011001",
22009 => "111111111101100000000001",
22010 => "000000110010111100100011",
22011 => "000010011000000100001010",
22012 => "000100010010011110000011",
22013 => "000110100110001100011100",
22014 => "001001001100010010001100",
22015 => "001011110011010111011010",
22016 => "001101001101100000011010",
22017 => "001100011001111110111000",
22018 => "001010001100001111010010",
22019 => "000111101100010010111100",
22020 => "000101101001110111011010",
22021 => "000100011000000111110110",
22022 => "000010100111110100111011",
22023 => "111111101110000100011110",
22024 => "111100010111110011000100",
22025 => "111001001000110101101000",
22026 => "110110100001011010001010",
22027 => "110100010011000111011000",
22028 => "110011000000000011000010",
22029 => "110011100101011110111000",
22030 => "110100110100010010000110",
22031 => "110110010011011001000011",
22032 => "111001000001011011100110",
22033 => "111100010100011000010101",
22034 => "111110101010001101100001",
22035 => "111111101010010011101011",
22036 => "111111101100111010101101",
22037 => "111110000010111100111010",
22038 => "111011000111001100000100",
22039 => "111000110000111000111110",
22040 => "110110100110110000110000",
22041 => "110100010001011011010000",
22042 => "110011010111101011111000",
22043 => "110100011101101111000011",
22044 => "110110101000001110111111",
22045 => "111001111001011001111101",
22046 => "111110010100100001000010",
22047 => "000010000110100111111000",
22048 => "000100100011101100011001",
22049 => "000110100111000001000110",
22050 => "001000101100000111011000",
22051 => "001010010011111000000111",
22052 => "001010100000111010111101",
22053 => "001001110100001100111011",
22054 => "001000010111011101101001",
22055 => "000101101101111011100101",
22056 => "000010111100101011011001",
22057 => "000000011100100100000011",
22058 => "111110111011111100010110",
22059 => "111111100011101011010010",
22060 => "000010000001010101000111",
22061 => "000101001000101011101101",
22062 => "000110101101010001000110",
22063 => "000110100001110011100011",
22064 => "000101110101010001111101",
22065 => "000100110101110100000000",
22066 => "000011101111000000001110",
22067 => "000010000101111110110000",
22068 => "000000111010011110010001",
22069 => "000001001010011100001010",
22070 => "000001100011001100010100",
22071 => "000001110100011010010000",
22072 => "000001111000010100011011",
22073 => "000001101010000100111011",
22074 => "000001010100110100100111",
22075 => "000000011010110010011111",
22076 => "111111010001000100101110",
22077 => "111100101110010110001100",
22078 => "110110001000011011110110",
22079 => "101011111011101000001000",
22080 => "100100001110000001001010",
22081 => "100011010111011111110011",
22082 => "100100011010011111011111",
22083 => "100100110111001110000111",
22084 => "101000011100100011111010",
22085 => "101110001001000101110000",
22086 => "110100010010011011001010",
22087 => "111010111110011101010101",
22088 => "000000101010110000101001",
22089 => "000110001011011110001110",
22090 => "001100001011101100011010",
22091 => "010000101111001001000010",
22092 => "010011101101001110101110",
22093 => "010110100001100100100110",
22094 => "011001010000011111111111",
22095 => "011010110000001101101001",
22096 => "011010101100101011101101",
22097 => "011010010000100111000111",
22098 => "011010000001010000101011",
22099 => "011001011111000101110011",
22100 => "011001001010011000101111",
22101 => "011000100010100000101110",
22102 => "010101000110101101111100",
22103 => "010000101001010010111000",
22104 => "001110111010000001001100",
22105 => "001110000000001110100110",
22106 => "001100000100010111001110",
22107 => "001011001111001011001011",
22108 => "001100000010100100111100",
22109 => "001101000111100110011100",
22110 => "001101100111000000010000",
22111 => "001011110101010110010110",
22112 => "000110100010010001101110",
22113 => "111111100000001111001111",
22114 => "111001011101100000010101",
22115 => "110101010111100110101110",
22116 => "110001101011110110010010",
22117 => "101101010010111101011110",
22118 => "101011100111110100011000",
22119 => "101101110010111100010100",
22120 => "101111110110000011111110",
22121 => "110001011111110101111110",
22122 => "110011111001001011000100",
22123 => "110110100100001110001100",
22124 => "111010101100101110111001",
22125 => "111111101010100001110010",
22126 => "000010001011111011110101",
22127 => "111111110001110011001101",
22128 => "111010001100000001000111",
22129 => "110100110011000011011010",
22130 => "101110001000101010010100",
22131 => "100110010010101111001101",
22132 => "100001101001111001110110",
22133 => "100000111101111100100011",
22134 => "100001101110011000111001",
22135 => "100010011011100000110100",
22136 => "100011101001011001100011",
22137 => "100100100011000111011011",
22138 => "100101001111001110001111",
22139 => "101010111101010100111010",
22140 => "110101000001111010100111",
22141 => "111101000111000101110111",
22142 => "000011101001011110001010",
22143 => "001011000110100110000110",
22144 => "010010000111010100111010",
22145 => "010101110111001110100000",
22146 => "010100111010101011010110",
22147 => "010010000101111001111010",
22148 => "010000010111101010011000",
22149 => "001110011000000000010000",
22150 => "001011000000000000101010",
22151 => "001000110001011101101110",
22152 => "001000110110100001110010",
22153 => "001001100001011100010010",
22154 => "001001111000010011111100",
22155 => "001001001011001001011011",
22156 => "000111111001000001100100",
22157 => "001000010101101010000010",
22158 => "001001101111001100101110",
22159 => "001001011100110011111011",
22160 => "000111110100110010001000",
22161 => "000111010001011011111111",
22162 => "001000101011001001010111",
22163 => "001010011101000111111011",
22164 => "001011101011110010001110",
22165 => "001101001010101111110000",
22166 => "001110101110001100110110",
22167 => "001111011010001000111010",
22168 => "001111001100011111110110",
22169 => "001101111010010001110010",
22170 => "001011011000111111110010",
22171 => "000111110010111010000100",
22172 => "000011000011010101001111",
22173 => "111101100111101010110010",
22174 => "110110111011101010111101",
22175 => "101110101101010111101000",
22176 => "100111111011011100110111",
22177 => "100100001010100011101111",
22178 => "100010001101111101101111",
22179 => "100001101000010111100101",
22180 => "100010111110000000110110",
22181 => "100111000100000001110101",
22182 => "101100010000111001101100",
22183 => "110000010000000010001010",
22184 => "110011101100001110110100",
22185 => "110111001010011011011001",
22186 => "111010011001101011110011",
22187 => "111100010100001010110100",
22188 => "111011010110100111111011",
22189 => "111000111001010010100001",
22190 => "110110011010001110010100",
22191 => "110011110000001101101110",
22192 => "110001010001100110111110",
22193 => "101111101000010111101100",
22194 => "110000111000010011011000",
22195 => "110101001110000110100111",
22196 => "111001110110101011011001",
22197 => "111110100101100001000010",
22198 => "000011100110100110111110",
22199 => "000111010001111110000000",
22200 => "001001010010111111010000",
22201 => "001010001110100100101110",
22202 => "001010110000000100011101",
22203 => "001010010000000110111010",
22204 => "000111111001000001110101",
22205 => "000101011001101101011111",
22206 => "000011111001000101011010",
22207 => "000010001111010011101110",
22208 => "000000010011111010000110",
22209 => "000000111000010000011111",
22210 => "000101110001011000001100",
22211 => "001011110101010011001101",
22212 => "010000110001111110101110",
22213 => "010101100001010000001110",
22214 => "011001010110001000011110",
22215 => "011011010010101001000101",
22216 => "011010001101110011011011",
22217 => "010101001010001010100110",
22218 => "001110101100001011110000",
22219 => "001000010000001111101011",
22220 => "111111010111100110010010",
22221 => "110011011100100100100010",
22222 => "101000011111010000100010",
22223 => "100010111001001100111111",
22224 => "100010010101001010000101",
22225 => "100100011010011100100011",
22226 => "101001000010111111111110",
22227 => "101111001100001110100110",
22228 => "110100111010011000000110",
22229 => "111010011000101110100010",
22230 => "111111011110010100000000",
22231 => "000011010100000111010100",
22232 => "000110000011101010001011",
22233 => "001000010100010011011100",
22234 => "001010001001001011110100",
22235 => "001011100101010000011000",
22236 => "001101010010000101100010",
22237 => "001110000111100110001110",
22238 => "001101011110010100111110",
22239 => "001101011000101101100010",
22240 => "001101111011111100000110",
22241 => "001110001101110011110010",
22242 => "001101011001011101101010",
22243 => "001010110110101000001011",
22244 => "001000001110111111010101",
22245 => "000100011000010011111101",
22246 => "111110000000010001111100",
22247 => "111001011000100110011101",
22248 => "111000011010010011100010",
22249 => "110111100101101000101101",
22250 => "110100101101001111001011",
22251 => "110010010101010011101100",
22252 => "110010111111011011110100",
22253 => "110100001011011100101100",
22254 => "110011011101111110100110",
22255 => "110001111100101111001110",
22256 => "110001001011110011100010",
22257 => "110010101011001010010110",
22258 => "110110111110000000101001",
22259 => "111100001100110010011100",
22260 => "000001110101010111100111",
22261 => "001000010010101010100000",
22262 => "001100010010100110001100",
22263 => "001100111101100001001000",
22264 => "001101110100000110000000",
22265 => "001111100100110101100000",
22266 => "010001001100000110011110",
22267 => "010001100100101110000010",
22268 => "010000001100111001001000",
22269 => "001100110110101010110110",
22270 => "000111100010010001101111",
22271 => "000011011100010010010001",
22272 => "000001101110000100011110",
22273 => "000000100011100000111100",
22274 => "111111110111001101010001",
22275 => "111110111100001111100010",
22276 => "111101100000110111011010",
22277 => "111100011110001011100110",
22278 => "111011111011011011001011",
22279 => "111010111101100111011111",
22280 => "111010000110101010000100",
22281 => "111100000111010101010000",
22282 => "000000100000001110000000",
22283 => "000110010000111000101100",
22284 => "001101001111010010000000",
22285 => "010011010101001010110010",
22286 => "011000001110110100110100",
22287 => "011010101010100000111111",
22288 => "011010000001011111000100",
22289 => "011000010001101101101011",
22290 => "010100110111111011010000",
22291 => "010000011000100001100100",
22292 => "001100001001000010000010",
22293 => "000111100100100100100110",
22294 => "000001000101100000010100",
22295 => "111000000001111100010101",
22296 => "101111110110000000001110",
22297 => "101010100011001001110100",
22298 => "101000010001010100111010",
22299 => "101001110110001010011100",
22300 => "101101101001101000011000",
22301 => "110001011111110111111010",
22302 => "110100010001001000111100",
22303 => "110110111111111101000111",
22304 => "111010110101110010001111",
22305 => "111111001000110001110101",
22306 => "000011100100000001011010",
22307 => "000110100101001000111111",
22308 => "001000101010011111001010",
22309 => "001011010001110110110100",
22310 => "001100010010100101110110",
22311 => "001010001100100101010100",
22312 => "000101110000100110000000",
22313 => "000000111111000100010111",
22314 => "111100010000111110100110",
22315 => "110111001100100001010000",
22316 => "110010111100000010101110",
22317 => "101111000101111000111100",
22318 => "101100010110101001010000",
22319 => "101011001101101001011010",
22320 => "101010000011010111100100",
22321 => "101001011011001111100000",
22322 => "101010001100110000110000",
22323 => "101100001110100100000010",
22324 => "101110011111101110101110",
22325 => "110001010100110100011010",
22326 => "110101110100011111110000",
22327 => "111010001010101001111001",
22328 => "111101110111111110100010",
22329 => "000001010000010010001011",
22330 => "000100011101110011100100",
22331 => "000111111100001100101100",
22332 => "001001110000011110010000",
22333 => "001010101011110100100100",
22334 => "001100001100001101010000",
22335 => "001100011110101000111010",
22336 => "001010011100000010010010",
22337 => "000110010110001001011001",
22338 => "000010010100110100111011",
22339 => "111111101101010000111111",
22340 => "111101011110000001001110",
22341 => "111010110000100001110101",
22342 => "110111111000101001101011",
22343 => "110110101010100111010001",
22344 => "110111111100111010010000",
22345 => "111011000011011110101111",
22346 => "111110101100000100111111",
22347 => "000010111100110001010000",
22348 => "001000101011000110010001",
22349 => "001101000100000011101000",
22350 => "001111010011001111000110",
22351 => "010001110001111111101110",
22352 => "010100000110001000011000",
22353 => "010100111101011101101010",
22354 => "010011011100100110100100",
22355 => "001111100111011101101010",
22356 => "001010001010011000001100",
22357 => "000011100100010110011101",
22358 => "111101001000110110001111",
22359 => "110111101001000110010101",
22360 => "110100001010000101110011",
22361 => "110010011110000010010100",
22362 => "110000000111011011100010",
22363 => "101100101011110010011100",
22364 => "101001101101111010001000",
22365 => "101000010100010000100110",
22366 => "101000011100100010011010",
22367 => "101010011010000101001110",
22368 => "101110001110110010111010",
22369 => "110010010001111000110000",
22370 => "110101101010000110010010",
22371 => "111000011100001000010000",
22372 => "111011100111011000110000",
22373 => "111111110101101101101111",
22374 => "000100010100111101111110",
22375 => "001000110100011111010011",
22376 => "001101001100101011000110",
22377 => "010001111111011010100100",
22378 => "010110100010101010001010",
22379 => "011000111100100011111011",
22380 => "011001110101000110001011",
22381 => "011001010011111010001000",
22382 => "010111001111111001011110",
22383 => "010101001110110101011000",
22384 => "010010111000101000101100",
22385 => "001110011011110011011110",
22386 => "000111111101101110001100",
22387 => "000000110011010100100011",
22388 => "111001010111110010111001",
22389 => "110001111111100011100010",
22390 => "101011001100001010000000",
22391 => "100101111101100011010110",
22392 => "100011101110111011100111",
22393 => "100011011000001111110101",
22394 => "100100000000000000110001",
22395 => "100101100111010100100011",
22396 => "100111010000100100010001",
22397 => "101001110001000001111100",
22398 => "101101011111011001010100",
22399 => "110010100110110011010010",
22400 => "111001101000110111000000",
22401 => "000000010011011110011001",
22402 => "000101100000010001001110",
22403 => "001001101100110101010010",
22404 => "001011010011000101010101",
22405 => "001000101001111100010001",
22406 => "000011100011000101101001",
22407 => "111110110101111110010011",
22408 => "111010011110001001010110",
22409 => "110110110100111111100010",
22410 => "110100010011011000101011",
22411 => "110001000101111011000010",
22412 => "101101111100011111001110",
22413 => "101100110010110101100110",
22414 => "101101000101010000100010",
22415 => "101101111110110010001010",
22416 => "101111101001000110110110",
22417 => "110001111110011110001010",
22418 => "110101000010111111100001",
22419 => "111000010011001100100110",
22420 => "111010011110001110010011",
22421 => "111100110101010111001110",
22422 => "000000101011101100011010",
22423 => "000101110010100000100100",
22424 => "001011101000010110010100",
22425 => "010001110101101101100010",
22426 => "011001010100000100101001",
22427 => "011110001001000000111001",
22428 => "011110000000010110101011",
22429 => "011101111011001011110110",
22430 => "011101101001010000101011",
22431 => "011100110011110001011001",
22432 => "011100011000011110001001",
22433 => "011000011010011110010101",
22434 => "010010100101001010010000",
22435 => "001110011100101101111100",
22436 => "001011101011111110000111",
22437 => "001010001110010011010101",
22438 => "001001100000001111101001",
22439 => "001010001111000101010011",
22440 => "001100011001101110001110",
22441 => "001110100101101000110010",
22442 => "010000100000001001101010",
22443 => "010001101111001101100000",
22444 => "010001111110101100010010",
22445 => "010000011110000111111010",
22446 => "001101101001000001100000",
22447 => "001011101010010101010011",
22448 => "001010110110011111111110",
22449 => "001010011110010001011011",
22450 => "001010101001100101110000",
22451 => "001010010011110001011100",
22452 => "000111111101000010010110",
22453 => "000100100011101001111100",
22454 => "000000110001111101011111",
22455 => "111100111111001111000111",
22456 => "111001000000011010110111",
22457 => "110011110101100110000110",
22458 => "101110111001110100111010",
22459 => "101000010110000111111000",
22460 => "100001101010100100100111",
22461 => "100001000000111000010011",
22462 => "100001101101011100110011",
22463 => "100001010011110100101101",
22464 => "100010100110100111101000",
22465 => "100011001111111100001111",
22466 => "100100010001010100010000",
22467 => "100101011011110110010111",
22468 => "100111010010000011011111",
22469 => "101101100110110111110100",
22470 => "110101101100110010010101",
22471 => "111101011000010010000000",
22472 => "000100100000000011111001",
22473 => "001010101110110011000011",
22474 => "010000000001011101101100",
22475 => "010010010000011001100010",
22476 => "010010011000000000101100",
22477 => "010001011110001110101110",
22478 => "001110101111000001101000",
22479 => "001010110111000001001010",
22480 => "000110100101110001010101",
22481 => "000011011000100010000011",
22482 => "000001100111011011000000",
22483 => "000001001110010100101100",
22484 => "000010010011111000110110",
22485 => "000011010100000011001101",
22486 => "000101011110011110101111",
22487 => "001010110111011011111110",
22488 => "010000111000110000010100",
22489 => "010101101110011111101100",
22490 => "011010011100001000000111",
22491 => "011100110000010011011001",
22492 => "011011111011110100100000",
22493 => "011011001001010000110001",
22494 => "011010010011110001101001",
22495 => "011001100010100000100011",
22496 => "011000110110101001010101",
22497 => "010111111011110001011110",
22498 => "010110111000100010110100",
22499 => "010001110011110101111100",
22500 => "001010010101111000101010",
22501 => "000011100100100010011111",
22502 => "111100001001100111001110",
22503 => "110101011100110011011110",
22504 => "101100010110101101100000",
22505 => "100011000110111011001101",
22506 => "100001001001110101010011",
22507 => "100001101001110100001000",
22508 => "100001101010100010110001",
22509 => "100001101110000010010011",
22510 => "100010000000010111010111",
22511 => "101001000111010010000110",
22512 => "110101001110010111100001",
22513 => "111101111000110110110110",
22514 => "000010101000001011101011",
22515 => "000110011001011100000001",
22516 => "001010011101010010101100",
22517 => "001101001010100110011000",
22518 => "001011101011001111110100",
22519 => "000110101101101110110101",
22520 => "000000111110010001010010",
22521 => "111011110011010010000010",
22522 => "111001010000110111101010",
22523 => "111000111010011110011110",
22524 => "110111101011011011100000",
22525 => "110111011111001000010100",
22526 => "111001100111010101011110",
22527 => "111011111101011011100001",
22528 => "111101110111100100000110",
22529 => "111101100101001100110001",
22530 => "111010100011111111001010",
22531 => "110110010010001010110111",
22532 => "110001101010001111111000",
22533 => "101101000010010101101110",
22534 => "101000100010101101110000",
22535 => "100110001100101100111011",
22536 => "100110100101000001100111",
22537 => "101000111101110100001010",
22538 => "101101101100100010010000",
22539 => "110011011110000011100110",
22540 => "111001100000011110100101",
22541 => "111111111110010001001101",
22542 => "000111000110111001001100",
22543 => "001110010110101110011010",
22544 => "010011110001101101100010",
22545 => "010111010010100101000010",
22546 => "010111111010111100110000",
22547 => "010100000011100011001010",
22548 => "001101110010100011000110",
22549 => "001000001101000000010011",
22550 => "000011010110110101111110",
22551 => "111100111111111111101010",
22552 => "110110000101010110111000",
22553 => "110000011011010110100110",
22554 => "101011000110000000110000",
22555 => "100110111100111011111110",
22556 => "100101000001100011101000",
22557 => "100101001100010111011011",
22558 => "100111010011101100100101",
22559 => "101010001110011100110010",
22560 => "101110010010011111111010",
22561 => "110011101110000100010100",
22562 => "111000100100011111001111",
22563 => "111011110100101001111010",
22564 => "111110111101000100000010",
22565 => "000011000110011101110000",
22566 => "000110101100001000000011",
22567 => "001001000101011010100010",
22568 => "001011100001011011101110",
22569 => "001101101100010000101110",
22570 => "001110001001101110101110",
22571 => "001100010001101100010000",
22572 => "001000101111010010000111",
22573 => "000100100010001011011001",
22574 => "000000011000000001010111",
22575 => "111100101100011111100000",
22576 => "111001111100000101010010",
22577 => "111000101110111011001111",
22578 => "111000110001001001100011",
22579 => "111001100000010110101001",
22580 => "111011000101000101000011",
22581 => "111101101011100000011111",
22582 => "000001010100010100110110",
22583 => "000101101000111111101000",
22584 => "001001110100110000010100",
22585 => "001100111101011101111010",
22586 => "001111011001001010000010",
22587 => "010001000110001110001000",
22588 => "010000110110101001011110",
22589 => "001111100110011010001100",
22590 => "001110101110001101000010",
22591 => "001101110111010011011100",
22592 => "001100011101100001001010",
22593 => "001001110110111000111010",
22594 => "000101111010000001110111",
22595 => "000001011100010010000000",
22596 => "111101101001110000100010",
22597 => "111010101010011010000110",
22598 => "110111111001001110111111",
22599 => "110101101111000000111010",
22600 => "110100001110000000011101",
22601 => "110010110101100001110000",
22602 => "110001010110100100101110",
22603 => "110000011010000110110100",
22604 => "110001010101111010001000",
22605 => "110011100011101100100100",
22606 => "110101100001001000001001",
22607 => "110110111100111101110111",
22608 => "110111111001110010111111",
22609 => "111000011111010110111101",
22610 => "111001101001110010011101",
22611 => "111100001100110111101010",
22612 => "111111001000000001100000",
22613 => "000001100000011010001101",
22614 => "000100010010101100001100",
22615 => "001000000111100010010001",
22616 => "001010111001000011111101",
22617 => "001010011011100111001000",
22618 => "001001000011011010100010",
22619 => "001000101000101101011001",
22620 => "000111100111110011101010",
22621 => "000110011101000101010010",
22622 => "000110011000001101100110",
22623 => "000110111010000101011111",
22624 => "000110110000101010110110",
22625 => "000101011100111110111000",
22626 => "000011101110111111011011",
22627 => "000001001000101000001110",
22628 => "111110101101110110000100",
22629 => "111111100111011001101011",
22630 => "000011101111110010110100",
22631 => "001000101001110101010101",
22632 => "001100110000010101001000",
22633 => "001111010000111011010010",
22634 => "010000010010100010110000",
22635 => "010010001000001100101110",
22636 => "010101100110000100110010",
22637 => "011000000011011101110001",
22638 => "011000100100010001101111",
22639 => "011000001100100000100001",
22640 => "011000101000010001100111",
22641 => "011000111111010010000101",
22642 => "010100110010111110101110",
22643 => "001100101110000100001010",
22644 => "000101011000110000001000",
22645 => "000000010100001101111000",
22646 => "111011100111111010100101",
22647 => "110101000101100010101110",
22648 => "101110101110001011101110",
22649 => "101010101001001110010010",
22650 => "101000111111100110010000",
22651 => "101010100000110100110100",
22652 => "101110011001011001101100",
22653 => "110100110010110101010111",
22654 => "111100011101001111000010",
22655 => "000001000110100010100011",
22656 => "000011001111000111000110",
22657 => "000101111110010000110010",
22658 => "001001101111010000010011",
22659 => "001100111100110000010110",
22660 => "001101111111010110110000",
22661 => "001101111100011100110110",
22662 => "001101100100000110001110",
22663 => "001100001010010001111110",
22664 => "001011110110110110111000",
22665 => "001100110110001010010100",
22666 => "001011000101101011000110",
22667 => "000110010001101001110101",
22668 => "000000010001101110111111",
22669 => "111010001100111101000100",
22670 => "110100110101000001011001",
22671 => "101100111001110011111100",
22672 => "100100001110001111001011",
22673 => "100001011011110110101011",
22674 => "100001111010110100111011",
22675 => "100010001000111000111001",
22676 => "100011111010110101010111",
22677 => "101001010011000100010000",
22678 => "110011100011001010010110",
22679 => "111110100010101010010100",
22680 => "000110001100101010101100",
22681 => "001011011100011000011000",
22682 => "001110101010010111000000",
22683 => "010000001101110011110000",
22684 => "001111101110011010111100",
22685 => "001100010001111000101000",
22686 => "000111010111110100001111",
22687 => "000011010010011011001010",
22688 => "000000100011010000111110",
22689 => "111100011010110000011110",
22690 => "110110100100011010110000",
22691 => "110011101001110001000110",
22692 => "110100111001011011010000",
22693 => "110111010101001110110010",
22694 => "111010001100011101111101",
22695 => "111101110011000111111000",
22696 => "111111011111011000010101",
22697 => "111101111010001000001010",
22698 => "111100001111001010000100",
22699 => "111100101010111101000110",
22700 => "111110010100100110011100",
22701 => "111111101000000010100000",
22702 => "000000100000001011000000",
22703 => "000010101001010101110001",
22704 => "000110001101001001010010",
22705 => "001001100000010001000010",
22706 => "001011010010001111010010",
22707 => "001011100000111000000000",
22708 => "001011010010110100100101",
22709 => "001011010100010011001001",
22710 => "001011100110010011100110",
22711 => "001100000001101101010100",
22712 => "001011111011000100011000",
22713 => "001010010001100011110010",
22714 => "000110111001111111101101",
22715 => "000011001100110110010100",
22716 => "000000011100000010100110",
22717 => "111110001110101100110100",
22718 => "111100000101000100100000",
22719 => "111010101010010000100111",
22720 => "111010000111001011011001",
22721 => "111010010111001110010010",
22722 => "111100011000001110000001",
22723 => "111111000000111011001001",
22724 => "000000000000100000000101",
22725 => "000000000011001110100101",
22726 => "000001001101000101110100",
22727 => "000100001100100111001101",
22728 => "000101111100100101010100",
22729 => "000011001000101111011010",
22730 => "111101101110011011110111",
22731 => "111000000100111100111000",
22732 => "110011100000111011011010",
22733 => "110001000000101000101010",
22734 => "101110000010001010110010",
22735 => "101010000101000100000010",
22736 => "100111111001111111001111",
22737 => "100111110110110010011101",
22738 => "101000101110100111000100",
22739 => "101001001111100100100000",
22740 => "101001010110101110011100",
22741 => "101001101010100101111000",
22742 => "101001001100111111000100",
22743 => "100111110100001101101011",
22744 => "100110110101011000010001",
22745 => "100111000101010010000011",
22746 => "100111110111001100101101",
22747 => "101000001110111101010010",
22748 => "101001000100010100101010",
22749 => "101011011001010100100000",
22750 => "101111011100101000101110",
22751 => "110100001101011111001100",
22752 => "111000011111111100101101",
22753 => "111101101101010101110011",
22754 => "000011111101100010110001",
22755 => "001000110010110000100111",
22756 => "001011101100100001111101",
22757 => "001101110101100000101000",
22758 => "001111001101111000100010",
22759 => "001110101110011110010000",
22760 => "001101011110100111010000",
22761 => "001101100101010110010100",
22762 => "001110010011000011101110",
22763 => "001110111010111001110100",
22764 => "010000001010111010110100",
22765 => "010010011100000101110100",
22766 => "010101010011011011000000",
22767 => "010111110000110000000110",
22768 => "011010011100001010100111",
22769 => "011101011110011011111111",
22770 => "011110011011110000011011",
22771 => "011101001110111010100100",
22772 => "011100001111110111110000",
22773 => "011011110011110001001111",
22774 => "011011010100010101011001",
22775 => "011010111000110010111001",
22776 => "011010011001100110011001",
22777 => "011000111110001100010001",
22778 => "010101010111110000010100",
22779 => "010001110000000000110010",
22780 => "010000111100000000000100",
22781 => "010000000010001011011000",
22782 => "001101010101010011101010",
22783 => "001010110100000101100000",
22784 => "001000100000111011101100",
22785 => "000110100001001111000001",
22786 => "000100011011100001110000",
22787 => "000001101011101100001010",
22788 => "111110011001010110000110",
22789 => "111001010111100010001010",
22790 => "110010110100101111111110",
22791 => "101010110010110001001000",
22792 => "100011001011110011000001",
22793 => "100000110010000111110001",
22794 => "100001010100111000100100",
22795 => "100000111111111010011001",
22796 => "100001010111100101010111",
22797 => "100010111100001010001011",
22798 => "100110010101100001101111",
22799 => "101011111111101110100110",
22800 => "110001001100010011101110",
22801 => "110101100101000111100111",
22802 => "111011001001101101101100",
22803 => "000000111000010110111000",
22804 => "000101100000011101111101",
22805 => "001001000001001011101110",
22806 => "001010000001101010011100",
22807 => "001000010100011100000010",
22808 => "000100010101010100011100",
22809 => "111110110011100011001100",
22810 => "111010000111011011110111",
22811 => "110101001010001010000000",
22812 => "101110111010100101011010",
22813 => "101010011101000100010010",
22814 => "101000101010111000101010",
22815 => "101001000010001110001110",
22816 => "101011100011001001111000",
22817 => "110000001010001110010100",
22818 => "110110110011010011010100",
22819 => "111101001101111110010000",
22820 => "000010011100000000101000",
22821 => "001000000010000010111110",
22822 => "001101001110111111000010",
22823 => "010000110101100100000000",
22824 => "010011000111001101000110",
22825 => "010011000000010111011000",
22826 => "010000100110101010100100",
22827 => "001110110111110000001010",
22828 => "001110110101110111110110",
22829 => "001110110110000011011000",
22830 => "001110000101011100111100",
22831 => "001101100110011011100100",
22832 => "001100100100010010011100",
22833 => "001000001101001111100110",
22834 => "000010110100111111000111",
22835 => "111111011110100001110111",
22836 => "111011111101001100101001",
22837 => "110111101110100110010010",
22838 => "110100000000100000110001",
22839 => "110001111000011010101110",
22840 => "110010110111101011101010",
22841 => "110101100111010010100110",
22842 => "111001001111011100011010",
22843 => "111110110101010000101011",
22844 => "000101101011000000011011",
22845 => "001011101010001010111001",
22846 => "001111010001100100100010",
22847 => "010000111001010101010110",
22848 => "010000110001001000110100",
22849 => "001110100101100111110100",
22850 => "001010100010010100011110",
22851 => "000100100001100111110101",
22852 => "111110110000011011111101",
22853 => "111011011110111010110100",
22854 => "111001011100110000110011",
22855 => "111000000101001010110110",
22856 => "111000010010001011010110",
22857 => "111010000100011110010010",
22858 => "111100101101000000110000",
22859 => "111111000100111010110100",
22860 => "000001010001000110111111",
22861 => "000100100101100110001010",
22862 => "001000011011111011010011",
22863 => "001010001001010001001100",
22864 => "001001010011001000110110",
22865 => "001000100110010011101010",
22866 => "001000111110101111011100",
22867 => "001000101000110011101101",
22868 => "000111001100010101110001",
22869 => "000101011001111100101011",
22870 => "000011001010010111011111",
22871 => "000000100001011101100101",
22872 => "111101100000111001100000",
22873 => "111001111110111000011101",
22874 => "110110000110010000011110",
22875 => "110011011100010100011010",
22876 => "110011111111110000001000",
22877 => "110101100000011001101000",
22878 => "110101100100111000110001",
22879 => "110101100011001111100010",
22880 => "110101010010101011110100",
22881 => "110100010000001011010000",
22882 => "110010100011110101001010",
22883 => "101111110100011100001110",
22884 => "101100110110010010010110",
22885 => "101001100010010001001100",
22886 => "100110101000001101100010",
22887 => "100110010000111111000110",
22888 => "100111000110010000010001",
22889 => "100111110110011110010000",
22890 => "101001110111001001000010",
22891 => "101101011011010010100110",
22892 => "110001101011100001011010",
22893 => "110101111010010110011100",
22894 => "111001110010011101101100",
22895 => "111101000110110101111001",
22896 => "111111111010001001100111",
22897 => "000010000001100000100101",
22898 => "000010100001001010011001",
22899 => "000010010001101101110101",
22900 => "000011010110001011110010",
22901 => "000100011010101001001110",
22902 => "000011110001101001100010",
22903 => "000011011110101110001110",
22904 => "000101000110110110000011",
22905 => "000111100110011100010001",
22906 => "001010011110000000011111",
22907 => "001110010000011110100010",
22908 => "010010010001000100110110",
22909 => "010101010001100111100000",
22910 => "011000000111011001111111",
22911 => "011011000101000110111001",
22912 => "011100101101010100000101",
22913 => "011100111010000000100100",
22914 => "011100011010010110101000",
22915 => "011011111001100011001111",
22916 => "011011010101110111110111",
22917 => "011010011111100100000111",
22918 => "011001000001100101111000",
22919 => "010100101010111100011010",
22920 => "001111001101000001110100",
22921 => "001101011110000011011010",
22922 => "001101100110011110000010",
22923 => "001011111010011110110010",
22924 => "001001100011010111001001",
22925 => "001001011010001111010111",
22926 => "001011010100101100011101",
22927 => "001011100100011101010101",
22928 => "001001101011001001010010",
22929 => "001000111100010100011110",
22930 => "001001111011000000100010",
22931 => "001000111101110010001010",
22932 => "000011010001001111011011",
22933 => "111011101011110100010010",
22934 => "110110000000000110001101",
22935 => "110010111010100101011000",
22936 => "110010001000101101110110",
22937 => "110010100010011100100110",
22938 => "110100001110111000000101",
22939 => "110110111111101000010010",
22940 => "110111000010101000101010",
22941 => "110100000110001001001111",
22942 => "110011000111110001110110",
22943 => "110101101100011011111000",
22944 => "111000110101000101101001",
22945 => "111001111101001101000100",
22946 => "111001101011000000001000",
22947 => "111010010111001101110100",
22948 => "111011101101000011100011",
22949 => "111011110101100110000111",
22950 => "111010100010100000100000",
22951 => "111000001100101110101010",
22952 => "110110000010001111101000",
22953 => "110100110000100110111100",
22954 => "110100010100111101000111",
22955 => "110100011110101111001111",
22956 => "110011000000010111010000",
22957 => "110000000000010100000110",
22958 => "101101011100000000000000",
22959 => "101011001100110010001010",
22960 => "101010101100001000110100",
22961 => "101100010100001010000010",
22962 => "101110011000110001011100",
22963 => "110001111110001100010000",
22964 => "110111010011110101100010",
22965 => "111010111111100100010110",
22966 => "111100000000111111011010",
22967 => "111110100101101101011100",
22968 => "000011111101111111110110",
22969 => "001000101010110111101100",
22970 => "001100100101010000000000",
22971 => "010000011111011000010100",
22972 => "010010110111001001100110",
22973 => "010010100110100010010000",
22974 => "001110111000111111000100",
22975 => "001001001010110011010100",
22976 => "000011101100110001000001",
22977 => "111110110010100010010101",
22978 => "111011111010001100011100",
22979 => "111100010010000011011100",
22980 => "111101110010111000101110",
22981 => "111110001110011010000011",
22982 => "111110110000010001010001",
22983 => "000001101000111011010001",
22984 => "000110000001100111111010",
22985 => "001001101111100110110000",
22986 => "001100000000111001100010",
22987 => "001100001101000101001110",
22988 => "001010110011100010001101",
22989 => "001001011011001100000110",
22990 => "000111101110011011001110",
22991 => "000101010100010011100010",
22992 => "000011110000101100010010",
22993 => "000011111001010110001100",
22994 => "000101000010011111110011",
22995 => "000110100110010001000110",
22996 => "001001011000111110100011",
22997 => "001100111111011010111010",
22998 => "001101111001001100100110",
22999 => "001010110110010000101111",
23000 => "000110010101001000000001",
23001 => "000010101010010100100100",
23002 => "111111110011001010111011",
23003 => "111100001100101011110010",
23004 => "111001000101100011000010",
23005 => "111000100000010000111011",
23006 => "111001010111011110101000",
23007 => "111011000101111110101100",
23008 => "111110001100111011111100",
23009 => "000001101010011110011001",
23010 => "000011111010110000011000",
23011 => "000100111001100111100010",
23012 => "000100111101101111100111",
23013 => "000010111100001110000010",
23014 => "111110011100000110011011",
23015 => "111000010111101100010011",
23016 => "110001100011000110101100",
23017 => "101011010110011101100100",
23018 => "100110011001010001000011",
23019 => "100011011101100110110111",
23020 => "100011100001111001100000",
23021 => "100100101111101011101111",
23022 => "100101011111111010110100",
23023 => "100110000110010111000111",
23024 => "100110101101010101011011",
23025 => "101000000110111101010100",
23026 => "101010100010100110011110",
23027 => "101100111100001110110100",
23028 => "101110100110001000011010",
23029 => "101111101000000101001000",
23030 => "110000101100110100000100",
23031 => "110001100001010010100100",
23032 => "110010010001001101101010",
23033 => "110100000111001010100100",
23034 => "110101011000010100001010",
23035 => "110101000110001010111111",
23036 => "110101101010000110110100",
23037 => "110111100011101001101011",
23038 => "111010000011001011100100",
23039 => "111101000111011011110011",
23040 => "000000011110101111010011",
23041 => "000100100010001000111110",
23042 => "001001001000001011110001",
23043 => "001101100011010000100010",
23044 => "010001011111100010101100",
23045 => "010100011101001000010110",
23046 => "010110101111001000001110",
23047 => "011000010101010110111101",
23048 => "011000100011010010110101",
23049 => "011000001001100000101010",
23050 => "011000010010010111010000",
23051 => "011000100101110101110010",
23052 => "010111011100011101000100",
23053 => "010100101001010000100010",
23054 => "010010001100101110011000",
23055 => "010001100110000000001100",
23056 => "010011010101000110100110",
23057 => "010110010101111011111110",
23058 => "010111110000101111010010",
23059 => "010110101001101001111110",
23060 => "010100101010100000000000",
23061 => "010010101100101000011000",
23062 => "001111101000001111101110",
23063 => "001011001111110110011111",
23064 => "000111110100100101010011",
23065 => "000110010010110010100010",
23066 => "000101111101100111010101",
23067 => "000110001010011011111000",
23068 => "000101000000011101111000",
23069 => "000010011001110010101101",
23070 => "000000101011101011001001",
23071 => "000000000111110110100100",
23072 => "111110111101010000100001",
23073 => "111011010110010000110101",
23074 => "110101110000101010110111",
23075 => "110000011010101101101000",
23076 => "101011100000010111101010",
23077 => "100111010011010100011000",
23078 => "100101110000110001011001",
23079 => "100111110011100011001110",
23080 => "101011111001001110000000",
23081 => "101110110011110000110010",
23082 => "110000110100110111010110",
23083 => "110100011101010110000110",
23084 => "110111101011010100111010",
23085 => "111000011100100100110010",
23086 => "111000010100100001010101",
23087 => "110111101011011011010110",
23088 => "110110001011001000000011",
23089 => "110101001110100100101101",
23090 => "110101110011001100100110",
23091 => "110110010001000011110110",
23092 => "110101011111101000010010",
23093 => "110101101100100010110101",
23094 => "111001000101011101111010",
23095 => "111111001000001000100111",
23096 => "000101100111101000010000",
23097 => "001010011011000001111001",
23098 => "001101001001011001101000",
23099 => "001110110010111001100100",
23100 => "010000011100100111110100",
23101 => "010010010010010011000100",
23102 => "010010111010100110011000",
23103 => "010010000001110110010000",
23104 => "010001010011111110111100",
23105 => "010000100100010000101010",
23106 => "001110110001111010010000",
23107 => "001100100101101110110100",
23108 => "001010011000101010001000",
23109 => "001000110001111011110110",
23110 => "001000011001010100111001",
23111 => "001001001000100000111000",
23112 => "001010111111100010010100",
23113 => "001101000010011101101010",
23114 => "001111001110001111100100",
23115 => "010001001100000100010000",
23116 => "001111101100110110101110",
23117 => "001010111101101001101000",
23118 => "000111111110111100111010",
23119 => "001001101001110011011110",
23120 => "001101000000001000110110",
23121 => "001101010001100110010100",
23122 => "001011001001001001010111",
23123 => "001001010111110010011001",
23124 => "000111000001011100000011",
23125 => "000010100000011111110101",
23126 => "111101000100101100011011",
23127 => "111001011101101111111010",
23128 => "110111010100011001011010",
23129 => "110011111001010101110100",
23130 => "101110000110000010101110",
23131 => "100111011100100000000001",
23132 => "100100010001000101101011",
23133 => "100110000000101101001001",
23134 => "101001101100000010111110",
23135 => "101110011010101110110000",
23136 => "110100111110010010111101",
23137 => "111101001000111111100011",
23138 => "000100111111011110001001",
23139 => "001001111111100001010001",
23140 => "001100101110100001011110",
23141 => "001110010100011110000100",
23142 => "001101110010000110100010",
23143 => "001010111101100100101110",
23144 => "001000001000000010010110",
23145 => "000111011101011101001100",
23146 => "000110111000111011011111",
23147 => "000100000000110111000100",
23148 => "000001000100100001010100",
23149 => "111111001000111001100100",
23150 => "111100111101000001101100",
23151 => "111010110010010011001000",
23152 => "111000010110000100000111",
23153 => "110101110000000010000010",
23154 => "110100101111000111001100",
23155 => "110101011001010010110100",
23156 => "110110011100011011001100",
23157 => "110110011000001011010000",
23158 => "110101010001011000011111",
23159 => "110101100101010000011110",
23160 => "110111101000001111101000",
23161 => "111001100010000101111010",
23162 => "111011000101101000110001",
23163 => "111100000000101001101000",
23164 => "111001111100001011000110",
23165 => "110101000100101001000111",
23166 => "110000101010000100011110",
23167 => "101011111110011100101010",
23168 => "100110011110100001101001",
23169 => "100100011011000000011101",
23170 => "100101101110100100111011",
23171 => "100110011111001101100111",
23172 => "100110110010011100010101",
23173 => "101000111110101000110110",
23174 => "101101100110110111001110",
23175 => "110011000100110011111110",
23176 => "111000100111001101101000",
23177 => "111101101000010111100101",
23178 => "000000100000001001100011",
23179 => "000001101100100101011000",
23180 => "000010010000001001011100",
23181 => "000001110101000111010001",
23182 => "000000011000100011011010",
23183 => "111110101111100101010010",
23184 => "111110010111011000100100",
23185 => "111110111011100010100001",
23186 => "111110110101101001010111",
23187 => "111111001111111010011110",
23188 => "000001111010101000011010",
23189 => "000110011101110000010001",
23190 => "001100111010101010000110",
23191 => "010011110111101111111110",
23192 => "011000011111000100010001",
23193 => "011011011001000011000011",
23194 => "011101001011100010101111",
23195 => "011101000001100100010101",
23196 => "011011110000100100101111",
23197 => "011001011000111010000010",
23198 => "010110010001101000111110",
23199 => "010011011000010011111000",
23200 => "010000100000010101110010",
23201 => "001101101100011110100000",
23202 => "001010110101101111010101",
23203 => "001001000101010111110010",
23204 => "001001001100000100111011",
23205 => "001010001001100111111110",
23206 => "001100001111011011001110",
23207 => "001111001010000111100100",
23208 => "010001101000001000010100",
23209 => "010010111011010000011100",
23210 => "010011000101111010111000",
23211 => "010001111100100010000010",
23212 => "001110010100100010001010",
23213 => "001001001110010011011001",
23214 => "000011100010000000101110",
23215 => "111100101110100101111100",
23216 => "110100000011010110100010",
23217 => "101001000100010001110110",
23218 => "100001101110111111011001",
23219 => "100001001111010010001011",
23220 => "100001100110100011111011",
23221 => "100000111001111100101101",
23222 => "100000101001100101000101",
23223 => "100010001110110001110000",
23224 => "100110111110110101001011",
23225 => "101010101000011100100110",
23226 => "101010000001110011101000",
23227 => "101000111010101100010100",
23228 => "101001111100010110000000",
23229 => "101010000000011111101100",
23230 => "100111010001101011100101",
23231 => "100101101001010111001010",
23232 => "100110100111101111011001",
23233 => "100111001101011010000101",
23234 => "100111010101111011010011",
23235 => "101001100110011101011010",
23236 => "101110101000101110111110",
23237 => "110101101011111010101101",
23238 => "111101010000011000010101",
23239 => "000010011100011010100001",
23240 => "000100100001100001001111",
23241 => "000101110010011101111100",
23242 => "000110111110001100110110",
23243 => "000110110110001100010010",
23244 => "000110000011100111011010",
23245 => "000110100010100000101110",
23246 => "000111011101011011001110",
23247 => "001000011010100001111000",
23248 => "001010011101001110101101",
23249 => "001011111110000000010010",
23250 => "001011111101001101000100",
23251 => "001010101001001000110001",
23252 => "001001010011010001000110",
23253 => "001010101011000110101100",
23254 => "001101010100100110111000",
23255 => "001110011100111011110110",
23256 => "001110111010000101011000",
23257 => "010000010000110011100110",
23258 => "010001011000001110101100",
23259 => "010000111011111001000110",
23260 => "010001101010001111001010",
23261 => "010100101010101110011010",
23262 => "011000110110100111110000",
23263 => "011101010000010100101111",
23264 => "011110001110001010000011",
23265 => "011100010111100001001011",
23266 => "011011000111011111111101",
23267 => "011001110110100110011001",
23268 => "010111111000100011111000",
23269 => "010011111110000111010100",
23270 => "001101101000011010111000",
23271 => "000110101011001101001000",
23272 => "000000011001111101010011",
23273 => "111011100101111100111000",
23274 => "110110110110111010001010",
23275 => "110010001111001001110000",
23276 => "110001100001111101110110",
23277 => "110101110100111111011110",
23278 => "111100001100101100100001",
23279 => "000001011011101000010011",
23280 => "000101001100010100100001",
23281 => "001001100001000000100011",
23282 => "001101100011110100101010",
23283 => "001110000000011111111000",
23284 => "001011110011100001000011",
23285 => "001010101010100010101001",
23286 => "001010001101111001011000",
23287 => "000111110001111011011110",
23288 => "000010101111110100000001",
23289 => "111100101000011110100110",
23290 => "110110011011000111000010",
23291 => "101111100110010010000100",
23292 => "101001010010101010111010",
23293 => "100101001011010100010101",
23294 => "100011100010000110110000",
23295 => "100100011010100011001101",
23296 => "100110011110010001000011",
23297 => "101000001010111001101110",
23298 => "101001101000001100100100",
23299 => "101011111000000000110000",
23300 => "101111000001101101000110",
23301 => "110001111000001011011100",
23302 => "110101000010100000111010",
23303 => "111001000000000001010110",
23304 => "111011101100111100110101",
23305 => "111100101000001011110100",
23306 => "111100110001100101010100",
23307 => "111011111001010010100101",
23308 => "111001100001100011100111",
23309 => "110110110000111101101010",
23310 => "110101100111100110101100",
23311 => "110110000100101010100010",
23312 => "110110011111001011001100",
23313 => "110110111100101100100011",
23314 => "110111111100001001001100",
23315 => "111000100110101001010001",
23316 => "111001011111111101001101",
23317 => "111011100111111100110110",
23318 => "111101110011001010001100",
23319 => "111111000001001010101100",
23320 => "000000101101010000110001",
23321 => "000100011111000111110100",
23322 => "001000111011000111011100",
23323 => "001100110010110101110010",
23324 => "010001001111000011101000",
23325 => "010101100001101000101100",
23326 => "010111111011111101010000",
23327 => "011001010010010000111101",
23328 => "011011011001110000111000",
23329 => "011100110111110100100110",
23330 => "011100000000101110000111",
23331 => "011010111010101010001011",
23332 => "011001011010100011110001",
23333 => "010110110111010001101110",
23334 => "010100111101011001100000",
23335 => "010010101110000111001010",
23336 => "010000001111010010001000",
23337 => "001110101001100011011010",
23338 => "001101110010111111110010",
23339 => "001110001010111110110110",
23340 => "001110101000110100010100",
23341 => "001110000000111010000000",
23342 => "001100011111001111100010",
23343 => "001010111111111100011000",
23344 => "001010001000000110011100",
23345 => "001001000010011111111111",
23346 => "000111011111001111101100",
23347 => "000100011000010101011000",
23348 => "000000110111010111111000",
23349 => "000000000110010100101010",
23350 => "000000111011100000010000",
23351 => "000001010011001001101001",
23352 => "111111100111010010010000",
23353 => "111100101101010100011100",
23354 => "111100000010101110001110",
23355 => "111100111100111000000000",
23356 => "111100111010001101100001",
23357 => "111010000011010001001011",
23358 => "110100101010000000101011",
23359 => "101110101000110110000100",
23360 => "100111101100000011001001",
23361 => "100010010111101101101011",
23362 => "100001011001000011101011",
23363 => "100001100111011100011001",
23364 => "100001001011101111001110",
23365 => "100001010110010111111100",
23366 => "100001110000110000010010",
23367 => "100010000001110011011101",
23368 => "100010110101011111101100",
23369 => "100011010100110000001111",
23370 => "100100010101001001010100",
23371 => "100111111001101000001100",
23372 => "101100001101101010010110",
23373 => "101111111011000110010010",
23374 => "110011010110101001100110",
23375 => "110111000001101011110100",
23376 => "111011111000001110001110",
23377 => "000000101111101101000101",
23378 => "000100011010101000111101",
23379 => "000110001110111111101010",
23380 => "000111001011001111101000",
23381 => "001001011011000110011000",
23382 => "001010010000101011101001",
23383 => "000110011001101110110111",
23384 => "000000111010111100110101",
23385 => "111110010101111101001101",
23386 => "111101010000110000011000",
23387 => "111011111010110100011010",
23388 => "111100110010011000101100",
23389 => "111110110000011111111011",
23390 => "000000110001111000100100",
23391 => "000011110011000000010011",
23392 => "000101100100011110010101",
23393 => "000101011101010011110010",
23394 => "000100000010001100010110",
23395 => "000010111010000111110101",
23396 => "000011001000000101011011",
23397 => "000001111001000010111100",
23398 => "000000001100011010001101",
23399 => "000001010001100101010010",
23400 => "000100011000010100010010",
23401 => "000101110110100011010010",
23402 => "000100101111110010101000",
23403 => "000110000111101010111000",
23404 => "001010110010101011010100",
23405 => "001110000001000010110110",
23406 => "001110001101101101010100",
23407 => "001100110100110110010000",
23408 => "001010111100010101010001",
23409 => "000111010101011111000100",
23410 => "000001110111011111010110",
23411 => "111100010000010011011101",
23412 => "110111111000110101111010",
23413 => "110101010010010101010110",
23414 => "110010111101011101011110",
23415 => "110001110011011100100110",
23416 => "110010111100010111110110",
23417 => "110100111000010100010100",
23418 => "110111110101110100010001",
23419 => "111011000100100011010000",
23420 => "111101110010100100110000",
23421 => "000001010001011001001100",
23422 => "000101101010110110111000",
23423 => "001001101000001100001000",
23424 => "001011110011111101001110",
23425 => "001101111111000101010010",
23426 => "010000100111000100100110",
23427 => "010001001011111111101010",
23428 => "010000011000111011000100",
23429 => "001111011011011111010110",
23430 => "001110010011111000001110",
23431 => "001100101111001010101010",
23432 => "001010000111101010111111",
23433 => "000111100011100010101101",
23434 => "000101011110110110100101",
23435 => "000011010011011010111110",
23436 => "000001000001000001100101",
23437 => "111110010101000101100000",
23438 => "111011010010110010010010",
23439 => "111000101101000111111001",
23440 => "110110110100000000000100",
23441 => "110100100101011110111110",
23442 => "110010010100100101100010",
23443 => "110010000000111001000110",
23444 => "110011100111111111000010",
23445 => "110100111111101101010111",
23446 => "110100111010111010011110",
23447 => "110100011111111111010001",
23448 => "110100100101000001010000",
23449 => "110101010110000001000011",
23450 => "110111101011111100101110",
23451 => "111010001111100110111011",
23452 => "111011000100101000110011",
23453 => "111010110110111100010000",
23454 => "111001001100011001001100",
23455 => "110100011101011101011101",
23456 => "101101111111011100001010",
23457 => "101000111100100001011100",
23458 => "100110111101110110011001",
23459 => "100111010001000010110011",
23460 => "100111110110001111000001",
23461 => "101000110101000111011010",
23462 => "101011100111011000000000",
23463 => "110000000011001100000000",
23464 => "110110101000100111101111",
23465 => "111111010111100111110101",
23466 => "001000000001110000010111",
23467 => "001111101110011101110100",
23468 => "010110111110001001001010",
23469 => "011100011110011000111100",
23470 => "011110001110010011010111",
23471 => "011110000011101010011001",
23472 => "011110010000011011111011",
23473 => "011100101110100111111111",
23474 => "011001000011111000101111",
23475 => "010101101011111111111110",
23476 => "010011100000011011001100",
23477 => "010010100011100001110110",
23478 => "010010101000111110000000",
23479 => "010010111101100010010000",
23480 => "010010101001001001111010",
23481 => "010010101010000010000110",
23482 => "010100001101001110111010",
23483 => "010110001010000100101110",
23484 => "010111001011011011101110",
23485 => "010110111000010110110110",
23486 => "010110011011101101000010",
23487 => "010110110110101001011110",
23488 => "010111010010000000100110",
23489 => "010111001100011110000110",
23490 => "010110111100000010000010",
23491 => "010111000111101001100010",
23492 => "010110110100001001110010",
23493 => "010110000111110101111100",
23494 => "010101110111101110001010",
23495 => "010010101011110100101100",
23496 => "001100010110010100000000",
23497 => "000101001101101100101111",
23498 => "111100111110011110011110",
23499 => "110100011001001100101101",
23500 => "101010010001110011000010",
23501 => "100001111011111111011001",
23502 => "100000111010011010100011",
23503 => "100001110001001010100011",
23504 => "100001011010000110011111",
23505 => "100010000011100000111101",
23506 => "100001110010010110000011",
23507 => "100001110001100000001010",
23508 => "100100101110010010000111",
23509 => "101000001101001000011010",
23510 => "101001000001010111011110",
23511 => "101000111100101101111000",
23512 => "101001100011011111100110",
23513 => "100111101110100100010001",
23514 => "100100101010010011010111",
23515 => "100011101111111110001000",
23516 => "100100011110110100001101",
23517 => "100111010000100110111111",
23518 => "101011101100100011110100",
23519 => "110000100100110010011000",
23520 => "110111000100111010101100",
23521 => "000000001100001001000000",
23522 => "001010010101101111101010",
23523 => "010001110100000011000000",
23524 => "010101000011101011100010",
23525 => "010101100110101000011000",
23526 => "010100101110011100001110",
23527 => "010001110100011110001000",
23528 => "001100010011110001011110",
23529 => "000111101010111101010101",
23530 => "000110011011101001011110",
23531 => "000110001101101010000000",
23532 => "000101011101000001011000",
23533 => "000100010001100011110100",
23534 => "000011101000001001011100",
23535 => "000100100000111001110010",
23536 => "000110001100100110011010",
23537 => "001000101010011010010100",
23538 => "001100100001001100111010",
23539 => "010001001111010011111110",
23540 => "010101111111111100100100",
23541 => "011001101101001010110111",
23542 => "011010110110000001011101",
23543 => "011001010111001100101001",
23544 => "010111110000100111001110",
23545 => "010111011001010110000010",
23546 => "010110111110011010101110",
23547 => "010101010000001111101110",
23548 => "010001101100111001000100",
23549 => "001100101111110010001010",
23550 => "000110110010101101001111",
23551 => "111111001010010111001100",
23552 => "110101111101100100010100",
23553 => "101101001010101001101100",
23554 => "100111010111011111110010",
23555 => "100100111011110000110011",
23556 => "100011111011001010000000",
23557 => "100011010110001010010001",
23558 => "100011101110010111001011",
23559 => "100100111011100111101100",
23560 => "100101111110011101101111",
23561 => "100111011011011011100111",
23562 => "101011011000111010000000",
23563 => "110010010011101101101000",
23564 => "111001010101001010011010",
23565 => "111101111110110010111011",
23566 => "000001111010111111010010",
23567 => "000101110001000011001001",
23568 => "000111000010011011001100",
23569 => "000101101011000011111001",
23570 => "000011011100010110101011",
23571 => "000001000111110000001110",
23572 => "111110000011001100011010",
23573 => "111001110111010101111111",
23574 => "110101001011000000000100",
23575 => "101111101010111111010100",
23576 => "101011101110000010001000",
23577 => "101100000110101111011100",
23578 => "101110001101110101111100",
23579 => "110000000110110100100010",
23580 => "110010110011010010000000",
23581 => "110110011101110010111111",
23582 => "111001111111010111001011",
23583 => "111011100011110100010110",
23584 => "111011101011010000011100",
23585 => "111011110100010011100000",
23586 => "111011010010100000000001",
23587 => "111010101010011101011000",
23588 => "111011001100100001100000",
23589 => "111011100110111100101001",
23590 => "111011100100011000000100",
23591 => "111100100111011001110101",
23592 => "111110100101000110010111",
23593 => "000001000011101010111000",
23594 => "000100100000000101101010",
23595 => "000111001111001100011010",
23596 => "000111001101110000111100",
23597 => "000110000101110111101110",
23598 => "000110010011011011111100",
23599 => "000110010010001101000000",
23600 => "000100000001000000111101",
23601 => "000000111110110001010001",
23602 => "111110111001011011101011",
23603 => "111101011111010100001010",
23604 => "111100011100000010001100",
23605 => "111101000110010000001110",
23606 => "111111101110001011111000",
23607 => "000010101001001110010011",
23608 => "000110010111101011111100",
23609 => "001011011011010101011110",
23610 => "010000000000101011010100",
23611 => "010011000110000111001000",
23612 => "010101101101010100011110",
23613 => "011000100100000100000111",
23614 => "011001101101000100001011",
23615 => "011001011111111111110100",
23616 => "011010001100010111101011",
23617 => "011010000110110001110111",
23618 => "011000101011001000000001",
23619 => "010101111011000111010010",
23620 => "010000001010111001010000",
23621 => "001000101110011111111110",
23622 => "000001100011110111110111",
23623 => "111100001010110000111100",
23624 => "111001100000001100110000",
23625 => "111000110101101110011110",
23626 => "111010100111101000110100",
23627 => "111110000110000110011101",
23628 => "000000101100100111001110",
23629 => "000010110010100010000100",
23630 => "000110010100110000100000",
23631 => "001010100010110011100111",
23632 => "001101110001000010110000",
23633 => "010000100001001111111110",
23634 => "010011100001001000011000",
23635 => "010101111111011010110110",
23636 => "010101110000100101000010",
23637 => "010001101011100001101100",
23638 => "001011000111100011111001",
23639 => "000011010110111001101011",
23640 => "111100100101011000110110",
23641 => "110110010000111100111000",
23642 => "101100111000010110010110",
23643 => "100100010000011110000010",
23644 => "100001100100110011100000",
23645 => "100001110110110111111101",
23646 => "100001100011000100011101",
23647 => "100001100001001011111111",
23648 => "100010100011111101111111",
23649 => "100011100101010011001011",
23650 => "100101010001110100100011",
23651 => "100111110101110011011011",
23652 => "101001101001000100111000",
23653 => "101011110000010101011000",
23654 => "101101111111111110010110",
23655 => "101110100010001010000100",
23656 => "101111000011101010011110",
23657 => "110010001010111111101100",
23658 => "110111110111100110111010",
23659 => "111101101001011111110000",
23660 => "000010011011111011001100",
23661 => "000110100010100100010010",
23662 => "001001011111000001111000",
23663 => "001100110101111100011000",
23664 => "001111111111110110101010",
23665 => "001111100010000011010100",
23666 => "001100100011000000111100",
23667 => "001001001110111111010000",
23668 => "000101101110100100110011",
23669 => "000011001000011001100100",
23670 => "000010011100110110000010",
23671 => "000011001001000011001100",
23672 => "000100110101000011001110",
23673 => "001000000010100111101100",
23674 => "001010111110110001000100",
23675 => "001011101011111111100010",
23676 => "001100010010000111110000",
23677 => "001100100111111110110010",
23678 => "001001110010000001111011",
23679 => "000100101101110000000110",
23680 => "000000011110110101011000",
23681 => "111111110110111111111111",
23682 => "000010001101101000100100",
23683 => "000010111010001111011011",
23684 => "000001011110101100000000",
23685 => "000001101001111111111110",
23686 => "000100111010000110100111",
23687 => "001001101010111000111010",
23688 => "001110011000010011111010",
23689 => "010010111010100101010110",
23690 => "010101001101011111100100",
23691 => "010011000101000111101000",
23692 => "001101101111111101011010",
23693 => "000110101111001010101010",
23694 => "111111010110011011000010",
23695 => "111000011001100001011100",
23696 => "110001111111101111100000",
23697 => "101101001011001100011100",
23698 => "101010001111001010001110",
23699 => "101001000000010100010100",
23700 => "101001100001011101011110",
23701 => "101011010011010110100100",
23702 => "101110000000010000111010",
23703 => "110010010001010010111000",
23704 => "111001001110110111001010",
23705 => "000001000110100100101111",
23706 => "000110110001101000010100",
23707 => "001010101101110011011101",
23708 => "001110000000101100010000",
23709 => "001111101110100111000010",
23710 => "001111001011000011110110",
23711 => "001100011001100011010100",
23712 => "001000000001010011100001",
23713 => "000011010011110000100010",
23714 => "111110101100001100011011",
23715 => "111010000111010100011100",
23716 => "110101101101010001001010",
23717 => "110001000000111111000110",
23718 => "101101011100111001100010",
23719 => "101100100010100100001110",
23720 => "101101000100000100110100",
23721 => "101110101101010011101010",
23722 => "110001010111001001010100",
23723 => "110011101001000111111110",
23724 => "110100000001011010001011",
23725 => "110010001100000000101010",
23726 => "110000100001111010101010",
23727 => "101111110111010001110000",
23728 => "110000000100101000001100",
23729 => "110010000101110100110100",
23730 => "110100001111000111001000",
23731 => "110101100101011011110100",
23732 => "110111000010011110111100",
23733 => "111000010001011100000100",
23734 => "111001000111101000110001",
23735 => "111010011001100001111101",
23736 => "111100011100001111010101",
23737 => "111101010010111110111010",
23738 => "111100100001110111010101",
23739 => "111011110101111000100010",
23740 => "111010100101000011100110",
23741 => "111000001111111011100010",
23742 => "110110001001111111011101",
23743 => "110110001101001000010110",
23744 => "111000111011001000001010",
23745 => "111100001011110001100010",
23746 => "111111010110101001001011",
23747 => "000011011000101110100110",
23748 => "001000010010111100011000",
23749 => "001101100011111100000010",
23750 => "010010111101110111001000",
23751 => "011000100001100111010001",
23752 => "011100100111011100011001",
23753 => "011110001011011001000111",
23754 => "011110011011101010100101",
23755 => "011110001010011101100100",
23756 => "011101100001010000111000",
23757 => "011100101111001100101111",
23758 => "011011111010100110011111",
23759 => "011010110111000101101010",
23760 => "011001110001011101101100",
23761 => "011001010000101000011001",
23762 => "011001000101100011100111",
23763 => "011000110010100000010011",
23764 => "011000011110110011011101",
23765 => "010111000101110010001000",
23766 => "010011000001101110011000",
23767 => "001111100100100000010010",
23768 => "001111100001010110100000",
23769 => "001110110000000110101100",
23770 => "001011110110101111001110",
23771 => "001001100111111111100010",
23772 => "001010001000001101001001",
23773 => "001101000011001111000000",
23774 => "001110001101010111011010",
23775 => "001110010111111010010110",
23776 => "010000110110101011110010",
23777 => "010011100010100101001000",
23778 => "010100000001111100011010",
23779 => "010001001011101100110100",
23780 => "001100001111111111010110",
23781 => "000110010011110001000010",
23782 => "111111110101111011010001",
23783 => "111000110101111111011110",
23784 => "101101000100001101100010",
23785 => "100010011100001111001101",
23786 => "100001001111011001100111",
23787 => "100010000100101010001101",
23788 => "100001011010010111011101",
23789 => "100001110011110110010111",
23790 => "100001110010100101010011",
23791 => "100001101101111110101110",
23792 => "100001110101001010001001",
23793 => "100010010110101001000110",
23794 => "100010111110100101011011",
23795 => "100011010000101110011000",
23796 => "100101110100100011101000",
23797 => "101001110101111110101110",
23798 => "101101010111110100011010",
23799 => "110010110111100111111000",
23800 => "111010110110111110101111",
23801 => "000000111111101111010101",
23802 => "000011010010101000101011",
23803 => "000100101111000111110100",
23804 => "000110111000001000101010",
23805 => "001001111100001000110101",
23806 => "001101010110101001001000",
23807 => "001110101000001100010100",
23808 => "001101111001110001000110",
23809 => "001011110011101100011110",
23810 => "001000111111000100100010",
23811 => "000111100100001100011101",
23812 => "000110010011000001001110",
23813 => "000100011110101111100111",
23814 => "000100111100110101010110",
23815 => "001000000000100001000100",
23816 => "001011001011001001000001",
23817 => "001101000010010111011110",
23818 => "001110001101001101010100",
23819 => "001110101111011010000100",
23820 => "001101001100000011111010",
23821 => "001001111101010011010010",
23822 => "000111101111011100101010",
23823 => "001001001001110011110101",
23824 => "001110011100001000111100",
23825 => "010010111000010000111110",
23826 => "010010000010101110111000",
23827 => "001111000100010001011000",
23828 => "001101100101111011110010",
23829 => "001011111101110111010100",
23830 => "001001101111100010011111",
23831 => "000111100101110110010010",
23832 => "000011100110011001101100",
23833 => "111101010110100111111101",
23834 => "110111011001111111101000",
23835 => "110011010010010001101010",
23836 => "110000001100100111100110",
23837 => "101101011001011001100100",
23838 => "101011011100111111101010",
23839 => "101010111111110001011100",
23840 => "101011110011101000100000",
23841 => "101100111100100000011110",
23842 => "101101000010100010111110",
23843 => "101011001001110010110100",
23844 => "101000011100101010101000",
23845 => "100111110110001010110001",
23846 => "101010001101010001010010",
23847 => "101101100001101000100100",
23848 => "110001001010110010011110",
23849 => "110110010000110101101110",
23850 => "111100010010101001100100",
23851 => "000001010011111001100101",
23852 => "000100100001010101100000",
23853 => "000110101100001101000101",
23854 => "000111111000001110000010",
23855 => "000111100100100010101100",
23856 => "000101111011101011110100",
23857 => "000010001010010011100111",
23858 => "111100111110111110110110",
23859 => "111000111101110001111110",
23860 => "110101010111001100110100",
23861 => "110001001110111001000010",
23862 => "101110100110101101010010",
23863 => "101110100110101100111110",
23864 => "110000010110110100000010",
23865 => "110010010111000100110010",
23866 => "110011011110111100111010",
23867 => "110011011110101001111000",
23868 => "110011100101011001001100",
23869 => "110101010111100101111010",
23870 => "111000001010011010010110",
23871 => "111010010000001101000000",
23872 => "111011001000110101001100",
23873 => "111011110001001101111100",
23874 => "111100111010001101001101",
23875 => "111101101000111011111101",
23876 => "111101001110101010001101",
23877 => "111100011011110011111010",
23878 => "111011110110101101010000",
23879 => "111010011111010000101111",
23880 => "110111111001111011001010",
23881 => "110101010010011101001000",
23882 => "110010100010001001000100",
23883 => "101111110001000110010100",
23884 => "101110011011110010110100",
23885 => "101110110100101001010000",
23886 => "110000011111111010110000",
23887 => "110010101001110101101010",
23888 => "110101001000000111001001",
23889 => "111000010111111010011101",
23890 => "111100010011111100010011",
23891 => "000001100100001101100101",
23892 => "000111010001100011111110",
23893 => "001011001011011110000100",
23894 => "001101110011001011111000",
23895 => "010000011000000010001010",
23896 => "010010000000000011011000",
23897 => "010001111100100100010000",
23898 => "010001000110001100000100",
23899 => "010000010001111000010000",
23900 => "001111101101000000001000",
23901 => "001111011011110010100000",
23902 => "001111100111000010100010",
23903 => "010000101000000110110000",
23904 => "010010000001011011110110",
23905 => "010011001011000011110000",
23906 => "010011110011001110110110",
23907 => "010011011000000110110110",
23908 => "010011010100010001110100",
23909 => "010101010110000111011010",
23910 => "011000000000101010101110",
23911 => "011000100100000101010000",
23912 => "010110110000111010011100",
23913 => "010101100111000001010000",
23914 => "010101111011101100101010",
23915 => "010101001010100100111110",
23916 => "010011011011111001011010",
23917 => "010010101101101111110100",
23918 => "010011000000001111110000",
23919 => "010011010111111000001000",
23920 => "010010101100111101111000",
23921 => "010000011000000101000100",
23922 => "001101000111001110101010",
23923 => "001010001010110100001010",
23924 => "000111111110011000011100",
23925 => "000100100010010101001001",
23926 => "111101100000101111111001",
23927 => "110100101111011111111000",
23928 => "101101111110001110000000",
23929 => "101001100010001001100000",
23930 => "100101101110101100001100",
23931 => "100011000110100101101010",
23932 => "100011101101001000110000",
23933 => "100110100001010011001011",
23934 => "100111110010111010000001",
23935 => "100110001111001000010101",
23936 => "100100010011100010111110",
23937 => "100100101110100111101111",
23938 => "100111001010111010000011",
23939 => "101001111111111001101010",
23940 => "101101100101101000000110",
23941 => "110010100100000000011110",
23942 => "111000111001101111111101",
23943 => "000000101001011111101111",
23944 => "000111110000101100011101",
23945 => "001100101111111100110000",
23946 => "010001111111111110110000",
23947 => "010111110000111101101100",
23948 => "011010001111000001100111",
23949 => "010111101100100000111000",
23950 => "010001001011100111100110",
23951 => "001000011101101001110110",
23952 => "111111101100001110011111",
23953 => "111000111110101100000110",
23954 => "110101100100111110001111",
23955 => "110100100010101000100111",
23956 => "110101100110100100101010",
23957 => "111001100111010001100010",
23958 => "111110101001000110101110",
23959 => "000010010111000100011110",
23960 => "000101000010010101101101",
23961 => "000111111100011100100011",
23962 => "001011010001010110010001",
23963 => "001110001111011100010110",
23964 => "010000100001101110111100",
23965 => "010010110010010100000010",
23966 => "010110010110001001010110",
23967 => "011001000101111010001101",
23968 => "010111101000011110010110",
23969 => "010100000001011111101010",
23970 => "010001101110100101001110",
23971 => "010010000101000000111100",
23972 => "010011101001110100100000",
23973 => "010011001010100011011010",
23974 => "001111011001111101001110",
23975 => "000111011100100000010100",
23976 => "111100100010010011001011",
23977 => "110010110100001100100010",
23978 => "101100110000111101010110",
23979 => "101010100011100101001100",
23980 => "101001000000110111110100",
23981 => "100111111000100111010001",
23982 => "101001111010000011001000",
23983 => "101101000001010101110000",
23984 => "110000001000010101110000",
23985 => "110011001110001100110110",
23986 => "110101101011001111001110",
23987 => "111010000101000111001100",
23988 => "000000111000000110101001",
23989 => "000111111001101100100110",
23990 => "001101010100111100001100",
23991 => "010000000101101011101110",
23992 => "010000001111110000101000",
23993 => "001101001011011111010000",
23994 => "001000010011001110001100",
23995 => "000011010111110011101001",
23996 => "111101100001100010101001",
23997 => "110111010111101100101000",
23998 => "110001110101101110110000",
23999 => "101101000000100100011010",
24000 => "101010100000110001110110",
24001 => "101011100001011100111100",
24002 => "101110000100100001100110",
24003 => "101111101110011000000110",
24004 => "110010000011010101101010",
24005 => "110111011011010100101010",
24006 => "111101100010101000101000",
24007 => "111111111010000110011001",
24008 => "111101001100101000001001",
24009 => "110111100000000001100000",
24010 => "110001001111011110011000",
24011 => "101100010000111001001110",
24012 => "101001100010111110011010",
24013 => "101000010011110000111000",
24014 => "100111011110101010001101",
24015 => "101000001001000111101000",
24016 => "101011101101001001110010",
24017 => "110000110100101010011000",
24018 => "110110011111111010010010",
24019 => "111100110001100011000010",
24020 => "000001011010101000101100",
24021 => "000010111001001111100010",
24022 => "000010001001001010010001",
24023 => "111111011000010011111010",
24024 => "111010011011011001001111",
24025 => "110101001110111001110000",
24026 => "110001110000110001010100",
24027 => "101111011110011011100110",
24028 => "101110011101001011000000",
24029 => "101111100000110111011000",
24030 => "110010001111110111110110",
24031 => "110110101100100100001110",
24032 => "111100101011101000100100",
24033 => "000011100010001010010100",
24034 => "001010100001111010000101",
24035 => "010000110101001101100110",
24036 => "010110100000000011110000",
24037 => "011010101101101101011111",
24038 => "011011111001011001011111",
24039 => "011010011010111110000001",
24040 => "011000000001110110000011",
24041 => "010101101111100111000110",
24042 => "010011010110111001110100",
24043 => "010001000000111000001100",
24044 => "001110111010111001110110",
24045 => "001100100110110110111100",
24046 => "001010010001110010000010",
24047 => "001000100100100000011000",
24048 => "000111100001100001001011",
24049 => "000110011000101111110000",
24050 => "000101111011001001011000",
24051 => "001000011000101000110100",
24052 => "001011111111101000110000",
24053 => "001100110100000011100000",
24054 => "001011001110000111110011",
24055 => "001001101110000001000010",
24056 => "001000110001000000000000",
24057 => "000111111000011111010101",
24058 => "000111100001101110111010",
24059 => "001000010000111000010000",
24060 => "001001101011101101111010",
24061 => "001010111010010101111010",
24062 => "001010010011111000111011",
24063 => "000110001101011101011101",
24064 => "000000011101100010101110",
24065 => "111100011110011100100011",
24066 => "111001111000111101000100",
24067 => "110111000011111001010100",
24068 => "110010011010001101101010",
24069 => "101010010010010001001000",
24070 => "100011000100000100110001",
24071 => "100001111100100100101001",
24072 => "100011101000100011111111",
24073 => "100100001110101100111000",
24074 => "100100101110111100100100",
24075 => "100101011111001111011110",
24076 => "100110000001001100000101",
24077 => "100111001110011100001001",
24078 => "101000110110111100101100",
24079 => "101001010100111011111010",
24080 => "101001011100110010100100",
24081 => "101011100100001111111010",
24082 => "101111111100110001110100",
24083 => "110101111000001010100110",
24084 => "111101010110100011001000",
24085 => "000101101100010111000110",
24086 => "001100100101001000101110",
24087 => "010000111110100111111000",
24088 => "010101011001101111101010",
24089 => "011011000100000001111010",
24090 => "011110101011100100111101",
24091 => "011110110111111101111100",
24092 => "011110101100001001100110",
24093 => "011110011110001000011111",
24094 => "011011011100000111100111",
24095 => "010110000100100110001010",
24096 => "010000011001010001110000",
24097 => "001011001011000101111100",
24098 => "000111111000000111111110",
24099 => "000110110011010001011100",
24100 => "000111000101001000000110",
24101 => "001000111111011001011100",
24102 => "001010101100110010110000",
24103 => "001001111000001101011110",
24104 => "001000000001110000000100",
24105 => "000111000100001001011001",
24106 => "001000000101001111110110",
24107 => "001011101000010001010001",
24108 => "001111110000111010000110",
24109 => "010011000100110010011000",
24110 => "010101100100011000110100",
24111 => "010110000000011000111010",
24112 => "010011111010000000110010",
24113 => "010000011000111101001110",
24114 => "001100000001110001110100",
24115 => "000110111100101110100110",
24116 => "000000111010111001000110",
24117 => "111001000111000001111110",
24118 => "110000010111100101001110",
24119 => "101001100100100011011110",
24120 => "100101101010001011111110",
24121 => "100011000101110010111111",
24122 => "100001110110100100111001",
24123 => "100011111010010001000001",
24124 => "101001010000011100011010",
24125 => "101110111011010110001000",
24126 => "110010100111111101011000",
24127 => "110100110001011011100111",
24128 => "110111101001010000010001",
24129 => "111100011111101101100110",
24130 => "000000110011101111000110",
24131 => "000010010100010100101011",
24132 => "000011001101000000010010",
24133 => "000101100111000101000011",
24134 => "001000001101100010101000",
24135 => "001001010111011010100010",
24136 => "001001001100111010111101",
24137 => "000111110001000101010001",
24138 => "000100110001000000001010",
24139 => "000001100001011100000100",
24140 => "111111001000010101011011",
24141 => "111100010010000000101010",
24142 => "111000100011110110000100",
24143 => "110110000101000011110110",
24144 => "110101111111011110100110",
24145 => "110111100110011100000100",
24146 => "111010100011000101000011",
24147 => "111110011000111000011010",
24148 => "000001111111100010110100",
24149 => "000100100010000010000110",
24150 => "000101000011000010111001",
24151 => "000011000001010010011110",
24152 => "000000010111011000000110",
24153 => "111111100000101111110100",
24154 => "111111011101111011010110",
24155 => "111101101001111011101011",
24156 => "111010101001010010000011",
24157 => "111000100101100100011110",
24158 => "110111100100100101010101",
24159 => "110110111101000000001101",
24160 => "110111000100111111010101",
24161 => "111000010110010100010000",
24162 => "111010001011111010001010",
24163 => "111011101000100000000011",
24164 => "111100001101111010111110",
24165 => "111011100010111000011111",
24166 => "111010001111010101000010",
24167 => "111010001001011001111010",
24168 => "111011011010100110000101",
24169 => "111101000000011001101100",
24170 => "111110111000001110010111",
24171 => "000000000111001110100000",
24172 => "111111010011010111101001",
24173 => "111101011100001001000100",
24174 => "111100100011010111010100",
24175 => "111101010110010010110001",
24176 => "111111001010011001101000",
24177 => "000001000101100111011000",
24178 => "000011100110001110111001",
24179 => "000111011110001000001010",
24180 => "001011110000010010011101",
24181 => "001111010011010010000110",
24182 => "010010010011111000011000",
24183 => "010101001001010010110010",
24184 => "010111011011001110111110",
24185 => "011000101001001000000101",
24186 => "011000011000000010001011",
24187 => "010101100011100011100110",
24188 => "001111111100111100011010",
24189 => "001001111000101001001001",
24190 => "000101001001111100111101",
24191 => "000001100101011110001101",
24192 => "000000000010100111111110",
24193 => "000001000011100000111001",
24194 => "000010110100100111011110",
24195 => "000101001010100100110000",
24196 => "001001010110010111100000",
24197 => "001101101011010001000010",
24198 => "001111111110000101000100",
24199 => "010000110110111001101000",
24200 => "010001010100011010111000",
24201 => "010001111010001110001000",
24202 => "010011010001110001110000",
24203 => "010011101101001000011000",
24204 => "001111111001110100011010",
24205 => "000111110011011001110001",
24206 => "111110110101000011010100",
24207 => "110111110111000100000010",
24208 => "110010100101111011000110",
24209 => "101100101011101110111100",
24210 => "100110010100100111011101",
24211 => "100010101101100100010101",
24212 => "100010010110000111110001",
24213 => "100010011110101111010111",
24214 => "100010000010001111101011",
24215 => "100001110001010000011011",
24216 => "100010000011101011000011",
24217 => "100010110010100000101100",
24218 => "100011101000110011101011",
24219 => "100100100000110000100011",
24220 => "100101011010001111100011",
24221 => "100101111100011100100111",
24222 => "100110001011011101001001",
24223 => "100110100010101011010111",
24224 => "100111001110110101010111",
24225 => "101001000101111111010100",
24226 => "101101010001101110110100",
24227 => "110011100000100001111100",
24228 => "111001111100100000011000",
24229 => "111111010111000100000010",
24230 => "000100011101011111101001",
24231 => "001001011110000111010101",
24232 => "001101101100111111110000",
24233 => "010001101001000101110110",
24234 => "010011110110001000010100",
24235 => "010001010010101001100110",
24236 => "001100101000111101010100",
24237 => "001010110101001011101111",
24238 => "001010110000010001101110",
24239 => "001001100001110101101111",
24240 => "000111110100001010011111",
24241 => "000111011000011000100110",
24242 => "001000101011110001001100",
24243 => "001001111100000010011110",
24244 => "001001010101101001110010",
24245 => "000111111000010101011010",
24246 => "000110101000010111010001",
24247 => "000110010011111110010011",
24248 => "001001001111001101001011",
24249 => "001111001110010010011110",
24250 => "010101001111011110100100",
24251 => "011010001011110100011100",
24252 => "011101001010000101010101",
24253 => "011100110110110101010101",
24254 => "011011000011011000110110",
24255 => "011001101100001000101100",
24256 => "011000011100111110111011",
24257 => "010111001111000010011010",
24258 => "010100100110111101000100",
24259 => "001101110100001101010110",
24260 => "000100000010101101010010",
24261 => "111011101011001111101101",
24262 => "110110010101110010010101",
24263 => "110010001011101101001110",
24264 => "101110010010001110011010",
24265 => "101100011010001101111000",
24266 => "101101011001100010000100",
24267 => "101111011100000101010010",
24268 => "110000110000101111111010",
24269 => "110000110001101011100010",
24270 => "110000101001101011010010",
24271 => "110011001000001100100110",
24272 => "111000001010111011111111",
24273 => "111100111111110010011000",
24274 => "000001010010011111010000",
24275 => "000110000000100011001101",
24276 => "001001100101111101000100",
24277 => "001001010110001010010100",
24278 => "000100011000100001010100",
24279 => "111100111000010011001110",
24280 => "110101101111111000111000",
24281 => "101111101110100110000110",
24282 => "101011000010111010100010",
24283 => "101000010101110100010000",
24284 => "100111011010101111000100",
24285 => "101000010111000001110000",
24286 => "101011001101010011001110",
24287 => "101110111010010010110010",
24288 => "110011001000110111011100",
24289 => "111000001001110110001101",
24290 => "111101010111111110110000",
24291 => "000001110000110100001010",
24292 => "000011101100110110100100",
24293 => "000001111110110100011110",
24294 => "111101101101010010011110",
24295 => "111001000101100011101000",
24296 => "110101001100000001101001",
24297 => "110010001110011101010100",
24298 => "110001010110011101111100",
24299 => "110011100011001100001110",
24300 => "110110101111001110011100",
24301 => "111000101000010011111011",
24302 => "111010011100101010100111",
24303 => "111101001100111010100001",
24304 => "111111010100111011100111",
24305 => "111111110101110111001010",
24306 => "111111001110100100101111",
24307 => "111110000001111000000000",
24308 => "111100101001100001010011",
24309 => "111100000000010111000111",
24310 => "111101000010111100001011",
24311 => "111110111100000011110001",
24312 => "000000100111110110111101",
24313 => "000010101101110110011110",
24314 => "000100110001101110101001",
24315 => "000110001001010100001010",
24316 => "001000111011001011110001",
24317 => "001101011010101001101000",
24318 => "010000001001100001010010",
24319 => "010000001000110100101100",
24320 => "001111100101001100001000",
24321 => "001110100011101110101100",
24322 => "001011110011000011110111",
24323 => "001000101101000101001101",
24324 => "000111011000010001011101",
24325 => "000111101010101001101001",
24326 => "001001011000010000110011",
24327 => "001100110010101111000100",
24328 => "010001000001110100111100",
24329 => "010101011000001011010110",
24330 => "011000101110010101011100",
24331 => "011001100001011110011011",
24332 => "011001001110000101001111",
24333 => "011001011101000000111000",
24334 => "011000110111010100100101",
24335 => "010111001111001110111110",
24336 => "010101011001100010000010",
24337 => "010010011011101101001000",
24338 => "001101111011011010110100",
24339 => "001000110000001100111110",
24340 => "000100010000100010011100",
24341 => "000001010101100000110110",
24342 => "111111000000001111101011",
24343 => "111101101000110100000010",
24344 => "111111101110111000100111",
24345 => "000100100010101000100011",
24346 => "001000100111001011011010",
24347 => "001010001001001101110000",
24348 => "001001011000010000101111",
24349 => "000111001001111010100111",
24350 => "000011000110010110000011",
24351 => "111101001011100110101110",
24352 => "110110111011111001111110",
24353 => "101111101011000000011100",
24354 => "100111010011011011001010",
24355 => "100010011000100100011001",
24356 => "100010000000110101101011",
24357 => "100010000010111100111011",
24358 => "100001110101100110000001",
24359 => "100010101001110001111010",
24360 => "100011010010100010100101",
24361 => "100011111001000011101011",
24362 => "100101011111001100111111",
24363 => "100110100100110011000100",
24364 => "100110011000110100010111",
24365 => "100111000111010100100111",
24366 => "101001111111101110111110",
24367 => "101110000100100010110000",
24368 => "110011000011011011101010",
24369 => "111000101001111000101000",
24370 => "111101011010010111100111",
24371 => "000001110001001110110100",
24372 => "000111000010010001101010",
24373 => "001011100000001011101010",
24374 => "001110001110000001110100",
24375 => "010001010111000101001110",
24376 => "010011110101100010000000",
24377 => "010001111000011100111010",
24378 => "001101101011001110100100",
24379 => "001100000101110101100110",
24380 => "001011010101011010100000",
24381 => "001000001001000000001010",
24382 => "000101010111111000101010",
24383 => "000101010000000100000110",
24384 => "000101010000101100000111",
24385 => "000100101111100001001101",
24386 => "000101001110001001100000",
24387 => "000101101001111010011000",
24388 => "000100001001010100110100",
24389 => "000001110101001001111000",
24390 => "000010100101000110111100",
24391 => "001000000010101000110111",
24392 => "001110011110011001001110",
24393 => "010010100101111100001010",
24394 => "010110000001101110100100",
24395 => "011001011010101100010011",
24396 => "011001100010000101000100",
24397 => "010101100001100101100010",
24398 => "010000101001001101100010",
24399 => "001100001001011010010100",
24400 => "000110000011101110100100",
24401 => "111110011110010001011110",
24402 => "110111110100110011010011",
24403 => "110010111110011101000100",
24404 => "101111100101011001001100",
24405 => "101101001001100001001010",
24406 => "101011000110010001011010",
24407 => "101010110011011011011110",
24408 => "101101111010000110000000",
24409 => "110010101000000000001000",
24410 => "110101111111001110010101",
24411 => "110111011001011010110100",
24412 => "111000100111100000011110",
24413 => "111011110010100101010110",
24414 => "000000010101011100011100",
24415 => "000011101100111111101001",
24416 => "000101111001000010001011",
24417 => "001000111011000110111100",
24418 => "001100101110000110100100",
24419 => "001111010000010111000010",
24420 => "001111010010001101011010",
24421 => "001100100101010010100010",
24422 => "000111010100011100001010",
24423 => "000001011000000111000011",
24424 => "111101010110111111010101",
24425 => "111010100100011011110010",
24426 => "110111001010110011111111",
24427 => "110101001111110110011110",
24428 => "110110111101100111100100",
24429 => "111010010001011011100100",
24430 => "111101011001000010010100",
24431 => "000000101100010100011100",
24432 => "000011010101101111011110",
24433 => "000100000010001000010101",
24434 => "000010111100010100100111",
24435 => "000000001100111100111101",
24436 => "111011110011010111001010",
24437 => "110111001000010111010010",
24438 => "110100000010010011111111",
24439 => "110010110000100001110010",
24440 => "110001111111010101001000",
24441 => "110000101011111100001100",
24442 => "101110111101001110111110",
24443 => "101101011001010101100110",
24444 => "101100100111111000000100",
24445 => "101101000101101000010100",
24446 => "101110110000011011101110",
24447 => "110001010010000101011100",
24448 => "110011110101111001010110",
24449 => "110101001001000100001010",
24450 => "110101000011000110111001",
24451 => "110101000010011110010110",
24452 => "110110000111011011101001",
24453 => "110111111001011100000100",
24454 => "111001111011100010111100",
24455 => "111100010000111010001001",
24456 => "111110010111101010110110",
24457 => "111111011011010011100100",
24458 => "000000000101101001111000",
24459 => "000001010001110001110101",
24460 => "000010100100010110100011",
24461 => "000100010110101101010111",
24462 => "000111100100101011011011",
24463 => "001011000000100011111101",
24464 => "001101011001010110101110",
24465 => "001110110110111111110010",
24466 => "001110111010000101001100",
24467 => "001101110111011110101110",
24468 => "001110000000000111010000",
24469 => "010000000000001001000100",
24470 => "010001101100100100011110",
24471 => "010001111110001101010110",
24472 => "010011010100010001111000",
24473 => "010111000100011110110100",
24474 => "011001110111001001011011",
24475 => "011001111111011100111111",
24476 => "011001110100111111111001",
24477 => "011001101001100001111010",
24478 => "011000110100010111100100",
24479 => "011000101010111010011110",
24480 => "011000101111110111000111",
24481 => "011000001010010110100101",
24482 => "010111010100110000110010",
24483 => "010100010001110000100110",
24484 => "001110001110000111111010",
24485 => "001000111001010011101110",
24486 => "000101110001000101000000",
24487 => "000010011111011011101101",
24488 => "111111000111101100000111",
24489 => "111101111011110110011000",
24490 => "111110101001101111010100",
24491 => "111110100011101011001001",
24492 => "111100110010111000100101",
24493 => "111011000100101110011010",
24494 => "111010010101100100101101",
24495 => "111001100001011001101000",
24496 => "110101111001010100111000",
24497 => "101101101011000111111000",
24498 => "100100110101101100101000",
24499 => "100000111101001010010001",
24500 => "100000111111011110111101",
24501 => "100001010001100110100101",
24502 => "100001011000100000010001",
24503 => "100001110110101101001011",
24504 => "100010111011001101000001",
24505 => "100100010000111000000011",
24506 => "100100101010101111111111",
24507 => "100100101000000100001001",
24508 => "100101000000111010111000",
24509 => "100101110110111001100001",
24510 => "101010000011100001100010",
24511 => "110011001101001011100110",
24512 => "111100011110111110011000",
24513 => "000011000000101000001001",
24514 => "001001001000001001011100",
24515 => "001110001111101010110010",
24516 => "010000000011011010000110",
24517 => "010000010001100000110000",
24518 => "010000100010111011011100",
24519 => "001111001000101111101000",
24520 => "001011010101100000001101",
24521 => "000111101100101110111011",
24522 => "000110011000111110101010",
24523 => "000110110010110100100110",
24524 => "000111110101100010001011",
24525 => "001001001011011010010000",
24526 => "001010011010101110011000",
24527 => "001100000000010011101110",
24528 => "001101110001011100010110",
24529 => "001101010010110001111110",
24530 => "001010000011011000000110",
24531 => "000110100000101000110110",
24532 => "000100010010001100111011",
24533 => "000100010001011110100110",
24534 => "000110010010011100001001",
24535 => "001000100011011101100000",
24536 => "001011101001011111111110",
24537 => "010000010000111001001010",
24538 => "010010101011010001110000",
24539 => "010001010001001011111000",
24540 => "001111110000000111000110",
24541 => "001111001111011110010110",
24542 => "001101000011111011111110",
24543 => "001000011110001111100110",
24544 => "000010100000010001010010",
24545 => "111011110001100111011110",
24546 => "110101000110001000011100",
24547 => "101110111111011101000010",
24548 => "101001011101100011100000",
24549 => "100101011100111100000011",
24550 => "100100000101110011100010",
24551 => "100101000001111000101110",
24552 => "100110111100010110011011",
24553 => "100111111101000000110111",
24554 => "100111011110111110110001",
24555 => "101000001010000100110100",
24556 => "101011010011101101010100",
24557 => "101110110011110101110100",
24558 => "110010110001111000111000",
24559 => "111000110010111001000000",
24560 => "111111001001011011101000",
24561 => "000100011001110000100101",
24562 => "001000110000100101101111",
24563 => "001010011111111000101000",
24564 => "001000101010000100100001",
24565 => "000101011101100000101000",
24566 => "000010110001001101100101",
24567 => "000000010111111011100000",
24568 => "111101101011010111111110",
24569 => "111011000110100111000101",
24570 => "111001011110011001101011",
24571 => "111000110100001110000001",
24572 => "111001100110011111001101",
24573 => "111100100110101100100001",
24574 => "000000011100011010001111",
24575 => "000011011010001111010000",
24576 => "000101111110001001000001",
24577 => "001000010000100101011110",
24578 => "001000100011000100110000",
24579 => "000110010001011100000001",
24580 => "000100000001101111000000",
24581 => "000100100001001100001101",
24582 => "000111000100011101100111",
24583 => "001001100001000100100001",
24584 => "001011000010001000101001",
24585 => "001011110001101010100000",
24586 => "001100101011000001111010",
24587 => "001110000010110110111010",
24588 => "001101110110011101100010",
24589 => "001011001111111100110111",
24590 => "001000100111100101101110",
24591 => "000110100001100001101010",
24592 => "000010111001011111011111",
24593 => "111110011000010011001101",
24594 => "111011101111011001111110",
24595 => "111011001000010001101001",
24596 => "111011000001011110011011",
24597 => "111011010011000100101100",
24598 => "111100011011010100010110",
24599 => "111110100000101101000000",
24600 => "000001100100110010001111",
24601 => "000101000000001011011110",
24602 => "001000000000000001011010",
24603 => "001010011010110111010110",
24604 => "001011100000010111010010",
24605 => "001001111000101111101111",
24606 => "000101111110110110000110",
24607 => "000001111101100101011011",
24608 => "111110101100010101110111",
24609 => "111011001010110110000010",
24610 => "110111101101011101100100",
24611 => "110110101001001101111000",
24612 => "111000111111100101100101",
24613 => "111101100000010100000011",
24614 => "000010101000001111011110",
24615 => "000111011010001001100111",
24616 => "001011100011101001001100",
24617 => "001111000111110101000000",
24618 => "010001111111000101011000",
24619 => "010100010001100011111100",
24620 => "010110010100010110001110",
24621 => "010111110100010000001110",
24622 => "010111101010001000101000",
24623 => "010101000100111101110010",
24624 => "010001010110110011010110",
24625 => "001110010011111000100000",
24626 => "001011011010010011101001",
24627 => "000111111110111110101000",
24628 => "000101100100101000110000",
24629 => "000101000010010010110110",
24630 => "000100111111101100001111",
24631 => "000011111110110101001011",
24632 => "000001110000000011010010",
24633 => "111110101110011001001111",
24634 => "111011010111100000110011",
24635 => "111001000011010110111010",
24636 => "111001010011110000111110",
24637 => "111010100010100111111100",
24638 => "111001001101101011111100",
24639 => "110100010100010001000110",
24640 => "101101111010110111110110",
24641 => "101000111001000100100110",
24642 => "100110001111110011000001",
24643 => "100101000101011111111101",
24644 => "100101000110110001101110",
24645 => "100101001111100010011000",
24646 => "100011100110011100000111",
24647 => "100001111000000111100001",
24648 => "100010010110010000000101",
24649 => "100011011000010000101101",
24650 => "100011110000111101000011",
24651 => "100011111100100110110110",
24652 => "100100011010011111000001",
24653 => "101000001010111011000110",
24654 => "110001001011011010010110",
24655 => "111100001000011010001011",
24656 => "000101110100000011010011",
24657 => "001101100111001100000110",
24658 => "010011010011010101101110",
24659 => "010111111001110001100100",
24660 => "011011101001011101011111",
24661 => "011011101110011010000101",
24662 => "010110111101111001101110",
24663 => "001111111111110011010000",
24664 => "001001000011100010010111",
24665 => "000010101010011000011000",
24666 => "111101010000110100101110",
24667 => "111000110101001110110000",
24668 => "110101010001110000011100",
24669 => "110100100000010010111100",
24670 => "110111111111011011000011",
24671 => "111100111111111001001010",
24672 => "000000001111110000011000",
24673 => "000010001100111000101101",
24674 => "000100100011011000110011",
24675 => "001000000001100010101110",
24676 => "001100000110101000110000",
24677 => "001110110111110010100110",
24678 => "010000001101011111111110",
24679 => "010001110101011010110010",
24680 => "010010001111000010010000",
24681 => "001110110111101111011110",
24682 => "001001100010001001110110",
24683 => "000101100010111001111001",
24684 => "000011110010011111011011",
24685 => "000010111000010100100010",
24686 => "000000101010100110101011",
24687 => "111101000110001000010101",
24688 => "111010000011001001010110",
24689 => "110111100010110110010010",
24690 => "110100011110101010111010",
24691 => "110001100001110100101100",
24692 => "101111101110001110111110",
24693 => "101110110000101110100100",
24694 => "101101101010110001111110",
24695 => "101011100111100000001000",
24696 => "101001000010010111111110",
24697 => "100111100100101001011000",
24698 => "100111110111011001011101",
24699 => "101001010111000001000000",
24700 => "101100101010110100000000",
24701 => "110010101000011110000000",
24702 => "111001101010001101000100",
24703 => "000000001000110001101101",
24704 => "000110011001101001011000",
24705 => "001011010101101101100100",
24706 => "001100100101011010101010",
24707 => "001010010011111100110010",
24708 => "000110000111011100001110",
24709 => "000001000110100000110011",
24710 => "111100001001011111000001",
24711 => "110111001110001101110010",
24712 => "110010101010110101011100",
24713 => "101111111000110100011010",
24714 => "101110101100000001011110",
24715 => "101110010110101110001000",
24716 => "101111010101011100110100",
24717 => "110000111000001111101010",
24718 => "110010001000101110110100",
24719 => "110011111001101010101000",
24720 => "110101101101001110010110",
24721 => "110110010011000011101001",
24722 => "110110011110111011001110",
24723 => "110111101011111100000010",
24724 => "111010010100110011111100",
24725 => "111101110000011100110100",
24726 => "000000100001000000011101",
24727 => "000010001110010100110010",
24728 => "000011111001100010100000",
24729 => "000101110101011110010000",
24730 => "000111010110001111010010",
24731 => "000111110000110010000010",
24732 => "000110111000001000101110",
24733 => "000101000111011011011000",
24734 => "000010101011001011001100",
24735 => "111111001011000011011000",
24736 => "111011001110011100000010",
24737 => "111000110111111111000100",
24738 => "111001001110100010101001",
24739 => "111011001111010101110000",
24740 => "111101110001100101111000",
24741 => "000000110000000010010100",
24742 => "000100001001110000000001",
24743 => "000111111110101000110100",
24744 => "001100001001101110010010",
24745 => "010000100000010110101110",
24746 => "010101101110011110100010",
24747 => "011011010101011101000010",
24748 => "011110100001010010001111",
24749 => "011110110010000100011111",
24750 => "011110011100101100011010",
24751 => "011101100110000000111011",
24752 => "011011001001001001001001",
24753 => "011000011001001110000001",
24754 => "010111000010001001001110",
24755 => "010111000010010111100000",
24756 => "010111011011000011100000",
24757 => "010111100000101110011000",
24758 => "010111011110110111101010",
24759 => "010111011000100100110110",
24760 => "010111000011110011101010",
24761 => "010110111110011011010010",
24762 => "010111000010111101011110",
24763 => "010110101100111111111010",
24764 => "010110011010111111111000",
24765 => "010110001100110001010010",
24766 => "010100010011111011111010",
24767 => "001111010001010010111100",
24768 => "000111100000101001110011",
24769 => "111111100100001100110110",
24770 => "111010000110101000101010",
24771 => "110111010001000101000101",
24772 => "110101111101100001010101",
24773 => "110110001000111001101111",
24774 => "110111100001001011001011",
24775 => "111000110110110010011001",
24776 => "111001001110111010101000",
24777 => "111000100100111000010100",
24778 => "111000001001001110010010",
24779 => "111001010111111101010101",
24780 => "111010011110000110010010",
24781 => "110111101110011010001111",
24782 => "110000111010101011100010",
24783 => "101001010011111011110000",
24784 => "100011110110010001101101",
24785 => "100001101011100010110011",
24786 => "100001101100011111011100",
24787 => "100001110110010110000111",
24788 => "100010000010110011001111",
24789 => "100010111001010000101101",
24790 => "100011110110000110010001",
24791 => "100100101101000000100010",
24792 => "100101010010110011011101",
24793 => "100101100011110101011001",
24794 => "101000010010011011000100",
24795 => "101111110010111111101100",
24796 => "111001011011110000111110",
24797 => "000010010110010110111011",
24798 => "001011011011010111101111",
24799 => "010100111101010010010000",
24800 => "011100010000001011101001",
24801 => "011110111111111111011100",
24802 => "011110001001101111101001",
24803 => "011100101011010100010011",
24804 => "011011110001101110000011",
24805 => "011010101000100110010011",
24806 => "011001100010010000101001",
24807 => "011000111001010110110011",
24808 => "010110101111100110101000",
24809 => "010001100101101010101010",
24810 => "001011010001110011111000",
24811 => "000110100001001010000000",
24812 => "000100001111100001001101",
24813 => "000011100110100010001010",
24814 => "000011000000110010011010",
24815 => "000010000111110101100100",
24816 => "000010011001100001101100",
24817 => "000101010001010101100100",
24818 => "001010011100011010010110",
24819 => "001111011011000110001110",
24820 => "010010000101001100100110",
24821 => "010100000001000100110100",
24822 => "010110100011000011000010",
24823 => "010110000001001001011000",
24824 => "001111111101101011011110",
24825 => "001000000011111110011001",
24826 => "000001111011011011110001",
24827 => "111100101011001100000010",
24828 => "110101111001100011000100",
24829 => "101101010101011110111000",
24830 => "100101111010111110110111",
24831 => "100010010100110001111101",
24832 => "100001011101100011110010",
24833 => "100001100110101101011101",
24834 => "100011000111111000101101",
24835 => "100110001101101101110011",
24836 => "101010010101000111011000",
24837 => "101110100001101111111100",
24838 => "110000011010110001010010",
24839 => "101110111110110000111010",
24840 => "101101001001000010100000",
24841 => "101101001010011101001100",
24842 => "101101100000111001111010",
24843 => "101101000101000000111110",
24844 => "101101010110111100011000",
24845 => "101111110011101101001110",
24846 => "110100101000001100011000",
24847 => "111010110011101011101010",
24848 => "000000001001001100111010",
24849 => "000011001110100100100111",
24850 => "000101000001101111101000",
24851 => "000111001000101010010000",
24852 => "001000111001101110110000",
24853 => "001000001000101110010000",
24854 => "000101001011000010100000",
24855 => "000010010010010100100011",
24856 => "111111001010011111011110",
24857 => "111010111010000100000100",
24858 => "110111011101100110110010",
24859 => "110101100010001001100101",
24860 => "110011001111111110100010",
24861 => "110000111100110000010000",
24862 => "110000011010000000011000",
24863 => "110000111111100011001110",
24864 => "110001011011100011101110",
24865 => "110010001000010000111000",
24866 => "110011111100111010010000",
24867 => "110111010001010110110110",
24868 => "111011110010010100101010",
24869 => "111111110100000010000001",
24870 => "000001100101010011101101",
24871 => "000001111000101001000100",
24872 => "000010101001011101000100",
24873 => "000011000001101110010100",
24874 => "000000100110111110101010",
24875 => "111100000010100011001011",
24876 => "110111110110110101100110",
24877 => "110011101101100100100000",
24878 => "101110010110000001111000",
24879 => "101001110111011101011000",
24880 => "101000010011000111101110",
24881 => "101000100100001101101100",
24882 => "101010001100100000110100",
24883 => "101101101100111001000000",
24884 => "110010001110011011101010",
24885 => "110111001110001000111111",
24886 => "111100101101011110001110",
24887 => "000010000011010011001010",
24888 => "000111001111010000010010",
24889 => "001100010100011001101010",
24890 => "010000001000111110111110",
24891 => "010010000110111010001010",
24892 => "010010110001001000111000",
24893 => "010010100100100100001010",
24894 => "010001101111011111011100",
24895 => "010000110100001011101100",
24896 => "010000101011000101011100",
24897 => "010001101100011100001110",
24898 => "010011010100111111110100",
24899 => "010100101110010010110010",
24900 => "010101110011111000010110",
24901 => "010111100101010100001000",
24902 => "011001011111110100001001",
24903 => "011001101101110110001010",
24904 => "011001101011000111110101",
24905 => "011011000001110001000111",
24906 => "011011100011001011100111",
24907 => "011010110110101100101001",
24908 => "011010101011101111100011",
24909 => "011010010100111000010111",
24910 => "011001111101001101111011",
24911 => "011001110100110110010101",
24912 => "010111101110011000011100",
24913 => "010100101111001011111110",
24914 => "010011010011111010010000",
24915 => "010001100110011111111100",
24916 => "001110101010100011100000",
24917 => "001100001010001100001010",
24918 => "001001111010100001000110",
24919 => "000110101111101001011101",
24920 => "000010100001000000101111",
24921 => "111110110001111010001000",
24922 => "111100101111110001000111",
24923 => "111001011110101011111101",
24924 => "110001101101000111111110",
24925 => "101000000100100010001100",
24926 => "100010001110001100100001",
24927 => "100001011111000110110001",
24928 => "100001111011111000011111",
24929 => "100001011111010111101001",
24930 => "100001111101010111001000",
24931 => "100010111111100010111101",
24932 => "100011011001111101010111",
24933 => "100100001011101110010111",
24934 => "100100101101101001101001",
24935 => "100100101111110001000101",
24936 => "100101100001101100001111",
24937 => "100101101010011000110011",
24938 => "100110100101011000010001",
24939 => "101101100011000011011000",
24940 => "111001000001001110101011",
24941 => "000011100001011101010110",
24942 => "001100110100001100000010",
24943 => "010101101001000110101000",
24944 => "011011100100111000100000",
24945 => "011101011001111000111011",
24946 => "011101001101111001100010",
24947 => "011011101101101010110011",
24948 => "010110001100001011110110",
24949 => "001101010001011101111110",
24950 => "000110010001110101101111",
24951 => "000011000011111110010111",
24952 => "000001010001011001000010",
24953 => "111111100111100000101101",
24954 => "111110101110011001111101",
24955 => "111111110110000010001000",
24956 => "000010001110110000011111",
24957 => "000011010110010011001111",
24958 => "000011010111001100000100",
24959 => "000100010111001001000111",
24960 => "000111001100011110001101",
24961 => "001100001000010000111010",
24962 => "010010100001000000110100",
24963 => "011000010110110101010111",
24964 => "011011101110000111111101",
24965 => "011100000110111110011101",
24966 => "011011001000011111111011",
24967 => "011001111000101111000101",
24968 => "010111101000001000101010",
24969 => "010100110101111001001100",
24970 => "010001111000010101000010",
24971 => "001100011100001110101000",
24972 => "000011010000100010110000",
24973 => "111000010100111101010000",
24974 => "101110110110110101000010",
24975 => "101000100001001110010100",
24976 => "100100010111100011100001",
24977 => "100001111001011100011001",
24978 => "100001111010000010001011",
24979 => "100011111010000000111111",
24980 => "100111001001011111100111",
24981 => "101010110110001111110110",
24982 => "101101101000010100101110",
24983 => "110000101100011000111010",
24984 => "110101101101011011110101",
24985 => "111010111000111101111010",
24986 => "111111001110011010110011",
24987 => "000011110100010101010111",
24988 => "000111011101111010111000",
24989 => "001000001001000100111110",
24990 => "000110010101011110000100",
24991 => "000011010011110111110000",
24992 => "111111001000100101010111",
24993 => "111001111110011110111100",
24994 => "110101001011111100000111",
24995 => "110001110010111110100100",
24996 => "101111111010101010110010",
24997 => "101111110111001001001000",
24998 => "110001011111100010010010",
24999 => "110011110001100011100110",
25000 => "110110001010100001001100",
25001 => "111000110110011111011111",
25002 => "111011110111001001001000",
25003 => "111110001010001000111011",
25004 => "111110011111101111100011",
25005 => "111101011010001001101001",
25006 => "111011100111011101101000",
25007 => "111000111101110100110001",
25008 => "110110111101110010000001",
25009 => "110111000101000001010110",
25010 => "111000100000001111010100",
25011 => "111011001001110010110001",
25012 => "111111000110111101001010",
25013 => "000010101110000001011100",
25014 => "000101110001001010011010",
25015 => "001001000110000001100010",
25016 => "001011001000011001010100",
25017 => "001010000101100110001000",
25018 => "000110101000010110100101",
25019 => "000010000001001001100101",
25020 => "111100001110110011100011",
25021 => "110101001111100001111100",
25022 => "101110111000011011100110",
25023 => "101011000101011001000000",
25024 => "101001110001001010010010",
25025 => "101010111100001110001110",
25026 => "101111001011010111001000",
25027 => "110101001000011010100000",
25028 => "111011001010001010100001",
25029 => "000001011011010100101010",
25030 => "000111101000011110111100",
25031 => "001100100101111101001100",
25032 => "001111111001110101100000",
25033 => "010000101101111111101100",
25034 => "001110001100111100001000",
25035 => "001010011000110001110111",
25036 => "000111110101110101111000",
25037 => "000101110011100000010000",
25038 => "000010101010110000011000",
25039 => "111111011001100101111000",
25040 => "111110001001001111001111",
25041 => "111111011111111011000110",
25042 => "000010000001110010011011",
25043 => "000100100101111111101010",
25044 => "000111110011101110010010",
25045 => "001011011011101100010000",
25046 => "001101110101011110010000",
25047 => "001111100010111000001110",
25048 => "010010010011000000110010",
25049 => "010100110100101010111110",
25050 => "010100110100110011111100",
25051 => "010011010001010010011100",
25052 => "010010000001101001011010",
25053 => "001111111100000010001010",
25054 => "001011100111100001001001",
25055 => "000110110010100001110001",
25056 => "000011101111011000000001",
25057 => "000011000111110000110011",
25058 => "000100001110101101010110",
25059 => "000100111000110100111111",
25060 => "000100001010101101111001",
25061 => "000011111110110011011010",
25062 => "000100101100010111100000",
25063 => "000100101110101101110101",
25064 => "000100011110111110101101",
25065 => "000011110100000111110100",
25066 => "111111010110111100000000",
25067 => "110101101110100110100010",
25068 => "101011101001110101101100",
25069 => "100110110101000001011111",
25070 => "100110011110100010011111",
25071 => "100110001111101101001111",
25072 => "100110001001000101011111",
25073 => "101000010011110111110010",
25074 => "101011011101001101010000",
25075 => "101101000001010011000000",
25076 => "101100000111111000101010",
25077 => "101010010100110100001000",
25078 => "101011000000111001001110",
25079 => "101111010000101110010000",
25080 => "110101000001110111001110",
25081 => "111010110101000011010000",
25082 => "000000100000110001011110",
25083 => "000110100110100000001110",
25084 => "001101000101010001100100",
25085 => "010010101111101110100110",
25086 => "010111100001001001001000",
25087 => "011011010101011000110011",
25088 => "011100101000001010110001",
25089 => "011011110000111011011101",
25090 => "011001000111101111110001",
25091 => "010011000000101101101110",
25092 => "001011001110010000100100",
25093 => "000100110100100111001010",
25094 => "111110111000101100011111",
25095 => "111001001110001000011010",
25096 => "110101000110011001101111",
25097 => "110010010000000101010110",
25098 => "110001111000101010011010",
25099 => "110100001101111110110001",
25100 => "110100111110101110111101",
25101 => "110010111010001110010100",
25102 => "110010111000001000100100",
25103 => "111000001101001100111010",
25104 => "000000101110110111101010",
25105 => "001000100001001101010110",
25106 => "001110011011101000111100",
25107 => "010011101001011001110110",
25108 => "010111100000010011001110",
25109 => "010111110001110001011100",
25110 => "010100101100111100111000",
25111 => "010000101010000110110110",
25112 => "001100001111100111011000",
25113 => "000110011011001000100100",
25114 => "111111100110100110000100",
25115 => "111000010101011011010111",
25116 => "110000010011101111101000",
25117 => "101001110100001001100110",
25118 => "100111010011010011001000",
25119 => "100110101001010010111011",
25120 => "100110010101101100000101",
25121 => "101000011000011011100000",
25122 => "101100011100001100011010",
25123 => "110000000011001100011100",
25124 => "110010111011001100101110",
25125 => "110101111111101101101111",
25126 => "111010001001000011011010",
25127 => "111111100110111111110011",
25128 => "000101000001001111100101",
25129 => "001001101000100100000110",
25130 => "001110011000001111110010",
25131 => "010011000101101000011110",
25132 => "010110011111000100101000",
25133 => "010111110101101001110110",
25134 => "010110000111100110110100",
25135 => "010000100100010000100110",
25136 => "001000110111011100010100",
25137 => "000001100110010101010010",
25138 => "111011001100001010001110",
25139 => "110100111101110110111100",
25140 => "110000000011010000111100",
25141 => "101110011010100000110110",
25142 => "101111011101100100010100",
25143 => "110001000111110100011100",
25144 => "110100000010010000010110",
25145 => "111001101010001001010101",
25146 => "111111111100000010000100",
25147 => "000011111111001010101111",
25148 => "000101010111101000110001",
25149 => "000100100001111101111111",
25150 => "000010010101010100010101",
25151 => "111111110011111101100101",
25152 => "111100101111111100101111",
25153 => "111001010110111000000010",
25154 => "110110111100000000010010",
25155 => "110101000011110011110010",
25156 => "110010010001000101010110",
25157 => "101111011010100011100000",
25158 => "101110101111111100010000",
25159 => "110000011100100001011000",
25160 => "110010110010101101110110",
25161 => "110101000101001101101001",
25162 => "110111001000100011010000",
25163 => "110111100010011011110000",
25164 => "110101101101100101100010",
25165 => "110011001101000110001110",
25166 => "110001101010001101010110",
25167 => "110001100011010111001000",
25168 => "110010001111110000010100",
25169 => "110011010001101001111110",
25170 => "110101011111101001110001",
25171 => "111001001011110000101100",
25172 => "111101011010101001100101",
25173 => "000010010000000101110111",
25174 => "001000001100001100101111",
25175 => "001110011010110001100100",
25176 => "010011101110100011010010",
25177 => "010111110111111100011100",
25178 => "011011000101110010100110",
25179 => "011100101101101111100001",
25180 => "011011111110010000110100",
25181 => "011001101100100000110111",
25182 => "010110110101100111111110",
25183 => "010011011101001011011110",
25184 => "010000011011110000101000",
25185 => "001110101010100110010100",
25186 => "001101010100111010001000",
25187 => "001011010111110111100111",
25188 => "001001010011100111000100",
25189 => "001000111001010011001100",
25190 => "001010110110011101111000",
25191 => "001101011001000001001100",
25192 => "001111011010010001011100",
25193 => "010001111110101010110100",
25194 => "010100010000000000010100",
25195 => "010011100010110011110110",
25196 => "010000100010110110001110",
25197 => "001110001101001111001110",
25198 => "001100011111001101000100",
25199 => "001001100100011010000011",
25200 => "000101110001010100010001",
25201 => "000010010100100101101010",
25202 => "111111010000010100000100",
25203 => "111100001100010101000101",
25204 => "111001001000011000001110",
25205 => "110110111000100010100010",
25206 => "110101111111001100110111",
25207 => "110011110111010101101110",
25208 => "101101100011100111011100",
25209 => "100101110000011110110001",
25210 => "100001110000010111000001",
25211 => "100010000001100001010111",
25212 => "100011011000010101011011",
25213 => "100100000101001100011101",
25214 => "100100110001100101100001",
25215 => "100111001001000101010011",
25216 => "101011000101111010110100",
25217 => "101101110001101111100010",
25218 => "101110011101000101111010",
25219 => "101111011101100011110110",
25220 => "110000101010101001011010",
25221 => "110001100011011100100000",
25222 => "110100111110110000000100",
25223 => "111010110001111100001100",
25224 => "111111010101110100011001",
25225 => "000011001010110010010110",
25226 => "001000011001111001111101",
25227 => "001110110110010110011110",
25228 => "010110001111110001111100",
25229 => "011100011001010000110011",
25230 => "011110001101111000001011",
25231 => "011101100001000011110011",
25232 => "011101001111011100111101",
25233 => "011100111110110100000011",
25234 => "011100011001111110101111",
25235 => "011011110001010100001001",
25236 => "011010111000100110111011",
25237 => "011010010110000111110011",
25238 => "011010000111001010101001",
25239 => "011001101101110100011000",
25240 => "011001110000101001010001",
25241 => "011000101010000011001101",
25242 => "010011001010000101110100",
25243 => "001010100011101111001011",
25244 => "000011011011001110100001",
25245 => "111111001100001011011001",
25246 => "111101000000110010000010",
25247 => "111101100011100010001111",
25248 => "000000110111011111001011",
25249 => "000100010101100101001110",
25250 => "000110001110000111111010",
25251 => "000111010010110010101000",
25252 => "001000010100011110010011",
25253 => "001001100111001011001111",
25254 => "001011000100100011010101",
25255 => "001010110000000000001111",
25256 => "000110100011100111011110",
25257 => "111110001111111111111110",
25258 => "110010110100011001011000",
25259 => "100111110110101111100100",
25260 => "100010001010010110000001",
25261 => "100001010110001001001001",
25262 => "100001100000011110011001",
25263 => "100001110111001011110111",
25264 => "100010011001011101111110",
25265 => "100001110110111000010111",
25266 => "100001011101001101000101",
25267 => "100010110000001000011111",
25268 => "100101011000001100100111",
25269 => "101010101000001000101100",
25270 => "110011000111010000011100",
25271 => "111011010110100100111101",
25272 => "000001011111000101011110",
25273 => "000111010101000101010100",
25274 => "001100100011110100101000",
25275 => "001110101001111100000100",
25276 => "001101100111111001001110",
25277 => "001011011100010000001111",
25278 => "001000101111010111111100",
25279 => "000101001101111010000110",
25280 => "000001011101000001000000",
25281 => "111101111111110111011011",
25282 => "111010011000111010000100",
25283 => "110110111011111111000110",
25284 => "110101011001000110101101",
25285 => "110110001110010100100100",
25286 => "111000000101111100100111",
25287 => "111011010101001111111111",
25288 => "000001001111111101001001",
25289 => "000111100101010100010011",
25290 => "001010110111100110110001",
25291 => "001011001100100001100000",
25292 => "001001110001110001010110",
25293 => "000111010011000101100001",
25294 => "000101110100011000010010",
25295 => "000110011110100001010110",
25296 => "000111011001011001010111",
25297 => "000110010101100100101001",
25298 => "000010111011110001101001",
25299 => "111110100000100100000010",
25300 => "111010010011101111110011",
25301 => "110110101101010001110000",
25302 => "110011111111111010111100",
25303 => "110001110101111011101100",
25304 => "110000000101111011010000",
25305 => "101111110100101101110110",
25306 => "110000010100010100001110",
25307 => "110000001010111101001000",
25308 => "110001001010110000011100",
25309 => "110100010000110100111100",
25310 => "110111001101001011010010",
25311 => "111001001011001100100010",
25312 => "111010101111100110101011",
25313 => "111011011000011001000000",
25314 => "111010111011110101000010",
25315 => "111010001110100010101001",
25316 => "111010000010001001111000",
25317 => "111010101001100100110100",
25318 => "111011111001010011011010",
25319 => "111101100010111110101000",
25320 => "111111001011010001000100",
25321 => "000000101011011011001011",
25322 => "000010111011111000000110",
25323 => "000110001111000011100000",
25324 => "001001110000111110011011",
25325 => "001101000000000110010000",
25326 => "001111111111101111010100",
25327 => "010010101111001011110110",
25328 => "010100010010011100011100",
25329 => "010011101010010101011010",
25330 => "010001101001100101000010",
25331 => "001111100011110011100000",
25332 => "001101101100101001000010",
25333 => "001100001011111000111110",
25334 => "001011010110000110001000",
25335 => "001011011011101101000010",
25336 => "001011110010000000111100",
25337 => "001011010011000111111100",
25338 => "001011000010100111010101",
25339 => "001100001100101011101110",
25340 => "001101011101101011011010",
25341 => "001110011011001101000000",
25342 => "001111110000110110110000",
25343 => "010000101100010111101100",
25344 => "010000011100001011100000",
25345 => "001101110110110001100100",
25346 => "000111111001010000100000",
25347 => "000000111101110111111100",
25348 => "111011110100001111000101",
25349 => "110111101010000111010100",
25350 => "110010010010100000100000",
25351 => "101010101101111101011000",
25352 => "100011101110011001110010",
25353 => "100001011100010010011001",
25354 => "100010011100111110111010",
25355 => "100010111101010000111001",
25356 => "100011000100010100111010",
25357 => "100011111101100100111111",
25358 => "100110000101011010111101",
25359 => "101001011101100001001110",
25360 => "101100001000111110101000",
25361 => "101100110001110000010100",
25362 => "101100001001111000001110",
25363 => "101010100000000100000100",
25364 => "101000100001100001110000",
25365 => "101000011000111011001010",
25366 => "101010100000011011011010",
25367 => "101101100111110111111110",
25368 => "110001111110111111110010",
25369 => "111000010011000110111101",
25370 => "111111001000011101000111",
25371 => "000100110111100110000111",
25372 => "001010010110101101100110",
25373 => "010000000110110110111110",
25374 => "010011111111010000001010",
25375 => "010100111000011000110110",
25376 => "010100000000010110110110",
25377 => "010001101111101111101110",
25378 => "001110011010111101001000",
25379 => "001100001011010000100010",
25380 => "001100000010011010010110",
25381 => "001100101010000000000100",
25382 => "001101010000111111000100",
25383 => "001101100110101100001010",
25384 => "001100111001010100110010",
25385 => "001011101101000011100000",
25386 => "001010101100101101100011",
25387 => "001000110000110110100011",
25388 => "000110001100111111100001",
25389 => "000101110111001001011110",
25390 => "001001010001011011010000",
25391 => "001110110110011110000110",
25392 => "010011011101001011100000",
25393 => "010101001101001001110000",
25394 => "010101110100011000111100",
25395 => "010111011110011101110010",
25396 => "011000110101000111000101",
25397 => "011000110010101111001111",
25398 => "011000110110100111100001",
25399 => "011000010110100100110100",
25400 => "010100010010001101100110",
25401 => "001100100100111111101010",
25402 => "000100010111001001101110",
25403 => "111101101100011101001000",
25404 => "111000011101011001101011",
25405 => "110011101001111001111110",
25406 => "101111000011001011101110",
25407 => "101100011011010111001110",
25408 => "101100011010100011011100",
25409 => "101101001110101001111000",
25410 => "101110001101011000011010",
25411 => "101111011010110010010000",
25412 => "110001000001101010111100",
25413 => "110101001010111100001011",
25414 => "111100101111111010101111",
25415 => "000100001000110111011100",
25416 => "001000110011110001100101",
25417 => "001100110010010010010000",
25418 => "001111011110100100001110",
25419 => "001101001010000000111010",
25420 => "000110011111111000010000",
25421 => "111110101110101010111000",
25422 => "110111011001010101011010",
25423 => "110001101001100101100100",
25424 => "101110010001111001010000",
25425 => "101100101011001101111000",
25426 => "101011101100011111100000",
25427 => "101100000100001001110010",
25428 => "101111011101110000100010",
25429 => "110100101100100001100111",
25430 => "111001011100111010101100",
25431 => "111110010100001000000110",
25432 => "000100010100101001001001",
25433 => "001001001100111010101100",
25434 => "001010001111100000101001",
25435 => "001000011100011011010011",
25436 => "000101111101011011000100",
25437 => "000010111001101010000111",
25438 => "111111011010101001010001",
25439 => "111100101000111100100101",
25440 => "111010111100010110110111",
25441 => "111010001001110100010101",
25442 => "111010000001010010010010",
25443 => "111001111011010000101000",
25444 => "111001100001011111100111",
25445 => "111001010110001110110100",
25446 => "111010010111000011000100",
25447 => "111100010001111010111010",
25448 => "111101101111101001111111",
25449 => "111110011001110010100011",
25450 => "111111000111101100010010",
25451 => "000000101110111010010001",
25452 => "000010010100000100110110",
25453 => "000010101100001110100110",
25454 => "000010110100111101101101",
25455 => "000010110100111110010110",
25456 => "000001101010000001110011",
25457 => "000000000100110011001001",
25458 => "000000001100111001101111",
25459 => "000011001011010001100010",
25460 => "000110010011010100010001",
25461 => "000110101011110111101111",
25462 => "000110001110010001001001",
25463 => "000110110010111011010000",
25464 => "000111000110110110110110",
25465 => "000110010100001111011010",
25466 => "000101110000100111101000",
25467 => "000111001011110000001011",
25468 => "001010001100100011111010",
25469 => "001101000000111101111010",
25470 => "001111100001011101001110",
25471 => "010010100011101001101110",
25472 => "010101000110000111100100",
25473 => "010101101111100000010110",
25474 => "010101000101000011110110",
25475 => "010100000100010110110110",
25476 => "010010010110100101100110",
25477 => "001110010010001001101110",
25478 => "000110111001110110111111",
25479 => "111110010010010000101001",
25480 => "111000000101110101010100",
25481 => "110101010011101001011010",
25482 => "110011001110010100001110",
25483 => "110001100000000000011100",
25484 => "110011011011101001011100",
25485 => "111000110001101110010011",
25486 => "111110101111010111001010",
25487 => "000100101011111101101111",
25488 => "001001111110100011110110",
25489 => "001100110101000000000100",
25490 => "001011100111111110101111",
25491 => "000110110000101101110001",
25492 => "000001101011110111010111",
25493 => "111100010010100001100011",
25494 => "110001100011101110110000",
25495 => "100101011000100111100000",
25496 => "100001000011000011010111",
25497 => "100001100101100001111001",
25498 => "100001010101001010010110",
25499 => "100001011111001001100000",
25500 => "100001111110101111011010",
25501 => "100100110001100111111000",
25502 => "101011100011111000010000",
25503 => "110001001010001011100110",
25504 => "110100001111100100101110",
25505 => "110111111001111011011100",
25506 => "111010011111001001010011",
25507 => "111001101100101100001010",
25508 => "110111001001010000111001",
25509 => "110101010011111010000111",
25510 => "110100110110110100010000",
25511 => "110101000101010101111100",
25512 => "110110001000100000011101",
25513 => "111000111000100010000010",
25514 => "111101001000011011111101",
25515 => "000010011011001100100111",
25516 => "001000011010111111010000",
25517 => "001101000101011011000000",
25518 => "001110111100001010010110",
25519 => "001111100010110100010110",
25520 => "001111101110010100001100",
25521 => "001110000011010100000010",
25522 => "001011000011011000111011",
25523 => "001001001101000000100111",
25524 => "001000010111010100100001",
25525 => "000110010101100110110001",
25526 => "000011000111101100110110",
25527 => "000000001111010010000110",
25528 => "111101010001001100100010",
25529 => "111001101001010111000010",
25530 => "110111000011100100110111",
25531 => "110110010000011100111110",
25532 => "110110011101110011101110",
25533 => "110111011001011010001110",
25534 => "111001100011000101101101",
25535 => "111101010101111000101000",
25536 => "000000000100101001110101",
25537 => "111111111011110001100010",
25538 => "000000100101110101000110",
25539 => "000011101111100000011111",
25540 => "000110101101100100110110",
25541 => "000111110111101111000010",
25542 => "001000001011100111000100",
25543 => "001000100011010100001010",
25544 => "000110111010111100010010",
25545 => "000010000100001110100001",
25546 => "111100001010011001011110",
25547 => "110111101010001100111011",
25548 => "110101000000100010011010",
25549 => "110010000110000000111010",
25550 => "101111010011111010000100",
25551 => "101111100010010011100000",
25552 => "110001101100010101111110",
25553 => "110100000001001001000010",
25554 => "110110110001111000011001",
25555 => "111010000001110000000000",
25556 => "111110101100101001011011",
25557 => "000101010110000110100100",
25558 => "001100001101100101110010",
25559 => "010001011010001000001100",
25560 => "010100110101101000101000",
25561 => "010111011001111111000010",
25562 => "011000111101001110111001",
25563 => "010111111011001111010110",
25564 => "010100110110101001000110",
25565 => "010010110111001111101010",
25566 => "010001110011010000110000",
25567 => "001110111100010000100100",
25568 => "001010011110000010111100",
25569 => "000110011101001101111011",
25570 => "000011111001001100100101",
25571 => "000001111110000011111110",
25572 => "000000010110000000111110",
25573 => "111111100101100010100001",
25574 => "111110110101101010101101",
25575 => "111110011001001001010011",
25576 => "111111001001100001000110",
25577 => "111111010000101010111111",
25578 => "111101111111101010001101",
25579 => "111100110010001100110000",
25580 => "111011100111000101000010",
25581 => "111001011010010001101100",
25582 => "110101110010100111110001",
25583 => "110001011010000110101110",
25584 => "101101011010101000001000",
25585 => "101010100101000001001100",
25586 => "101001011111100110001100",
25587 => "101010001001110110000100",
25588 => "101011100101111110000100",
25589 => "101100111011101111000100",
25590 => "101101011000010010110110",
25591 => "101101111011101101010100",
25592 => "110000101001110111101010",
25593 => "110011111101010011111110",
25594 => "110110010100000001101001",
25595 => "111000111001000111110000",
25596 => "111011000001010110100110",
25597 => "111011111110001011101011",
25598 => "111100011111010011010110",
25599 => "111100110111010000110101",
25600 => "111100111101110100111010",
25601 => "111100110101101101000110",
25602 => "111110010011111000110100",
25603 => "000001111100001110101000",
25604 => "000101100100100001101111",
25605 => "001001000101011100000101",
25606 => "001100111011111111100110",
25607 => "001111101100010011010010",
25608 => "010000100011110010100010",
25609 => "010000011101100110100110",
25610 => "010001001001110011111000",
25611 => "010011001101101000000000",
25612 => "010101111100000101000100",
25613 => "011001001011111011000001",
25614 => "011100000001001110111110",
25615 => "011100100100011111101101",
25616 => "011011110010111000001101",
25617 => "011011010110000100100000",
25618 => "011010100110011001000111",
25619 => "011010000000011011001011",
25620 => "011001110100000111101010",
25621 => "011001101001001011001111",
25622 => "011001010101111000010011",
25623 => "010101010010010111100110",
25624 => "001101011011000110011100",
25625 => "000111100100001011001001",
25626 => "000100001111001111100100",
25627 => "000000111110000100111000",
25628 => "111110001010111010111010",
25629 => "111101001110100011001000",
25630 => "111111011010100101001101",
25631 => "000010111100111100111000",
25632 => "000100101100111111001000",
25633 => "000100101111011001000010",
25634 => "000100010111000011110110",
25635 => "000100001000101010000101",
25636 => "000011011000000111111100",
25637 => "111111111101010000011000",
25638 => "111000110111111000001101",
25639 => "101111010011011011111010",
25640 => "100110011000101101001100",
25641 => "100001110000001111100001",
25642 => "100001000001000010111011",
25643 => "100001010000110010100111",
25644 => "100001101011110000001111",
25645 => "100010011001111100001111",
25646 => "100100011000110101000101",
25647 => "100111111111011111101011",
25648 => "101011001010110010100010",
25649 => "101101111110001000111010",
25650 => "110010001001111011000000",
25651 => "110110100100011111000010",
25652 => "111000001111100100000111",
25653 => "110111010100000001001100",
25654 => "111000010100001110111100",
25655 => "111100011111101001010101",
25656 => "111111111110010111110100",
25657 => "000010011010100010010111",
25658 => "000110100100010110010011",
25659 => "001100000100000110111100",
25660 => "010001000000111110001100",
25661 => "010100011100111111000000",
25662 => "010101101000111100110110",
25663 => "010101011000100000011100",
25664 => "010101000011011000000010",
25665 => "010100001010010110111110",
25666 => "010010001000101000011110",
25667 => "001111000111010001010000",
25668 => "001011110101000001110110",
25669 => "001000110100010101010111",
25670 => "000101101111111011011101",
25671 => "000010111111010011011100",
25672 => "111111011110110101111000",
25673 => "111010011001010011011101",
25674 => "110110010110000100000011",
25675 => "110100101011111010000001",
25676 => "110101001101100111110101",
25677 => "110111011001101000011100",
25678 => "111010000010001001010110",
25679 => "111101011101110000101010",
25680 => "000001000100111010101010",
25681 => "000010101000101101000001",
25682 => "000010001101011010000100",
25683 => "000010111110101011110100",
25684 => "000110001111101000111000",
25685 => "000111011111011110101110",
25686 => "000100010100111011101100",
25687 => "111111110010000100101111",
25688 => "111011100001111110100000",
25689 => "110110011000101101101100",
25690 => "101110000011011101101010",
25691 => "100101000010100111101001",
25692 => "100001010100111100100101",
25693 => "100001100000101000000111",
25694 => "100001111010011110101001",
25695 => "100011000101110111011001",
25696 => "100011111110110000100101",
25697 => "100100110010111101101101",
25698 => "101001010000101111101010",
25699 => "110000110100000011000110",
25700 => "110111110100111100111011",
25701 => "111110010010011001110011",
25702 => "000101011101010011100000",
25703 => "001011101011010011101100",
25704 => "001110001110001111101000",
25705 => "001101011010010000001110",
25706 => "001100001110111010111100",
25707 => "001011111000010100110110",
25708 => "001011000011100000100010",
25709 => "001001100100001010010100",
25710 => "001000010111000011001010",
25711 => "000111011001001110001101",
25712 => "000111000111000111011100",
25713 => "000111100010010110111111",
25714 => "000110110000110101110101",
25715 => "000101100001101100101011",
25716 => "000110000011000101111101",
25717 => "000111110100101011101010",
25718 => "001001100100010110000111",
25719 => "001010000011110001101110",
25720 => "001001100101100010111110",
25721 => "001000110001000100000000",
25722 => "000110110010111001010110",
25723 => "000100111110111111111001",
25724 => "000100000101000100010001",
25725 => "000011011100100010000010",
25726 => "000011100010100011011011",
25727 => "000011001101000011010010",
25728 => "000010010010110011110101",
25729 => "000001110110010011010001",
25730 => "000001010100100110000110",
25731 => "000000110011011001101110",
25732 => "000000000000011110000110",
25733 => "111110111111011110001000",
25734 => "111110100110000010001010",
25735 => "111101110010011111001111",
25736 => "111100000001000101110101",
25737 => "111001101011011001100001",
25738 => "110110100000001011100110",
25739 => "110011010001111110111000",
25740 => "110001100010010001101010",
25741 => "110001001111111011010010",
25742 => "110001101010111011010100",
25743 => "110010011101001111111010",
25744 => "110010101101111101100110",
25745 => "110001111101000100010100",
25746 => "110001000111110101111100",
25747 => "110001110000011010111010",
25748 => "110100001011010010001110",
25749 => "110110111110101010001000",
25750 => "111010001101110011010100",
25751 => "111110010111011100110011",
25752 => "000001100101000110100101",
25753 => "000011100000000101010000",
25754 => "000110010110111010011100",
25755 => "001010110010111001000111",
25756 => "001110110101111101011010",
25757 => "010001100010101111001000",
25758 => "010100010001100001101010",
25759 => "010111011111011100001010",
25760 => "011001100110001011111101",
25761 => "011001011000000000001101",
25762 => "010111110011001010011100",
25763 => "010100101110011011101010",
25764 => "001111011000000011001110",
25765 => "001010111001000100110110",
25766 => "001000001100001000011000",
25767 => "000100111111010101011001",
25768 => "000001111100110111000110",
25769 => "111111110111010100110110",
25770 => "111111100001101111010000",
25771 => "000001001101101101111111",
25772 => "000011101100111011000010",
25773 => "000111011001110010001101",
25774 => "001011001010000101100010",
25775 => "001101110010001101101110",
25776 => "010000100011000101110000",
25777 => "010010010011111011101110",
25778 => "010001100010101110101000",
25779 => "001111000010010111101100",
25780 => "001100011111001001110110",
25781 => "001001011100100011010100",
25782 => "000001111111101010110101",
25783 => "110111001011000110101100",
25784 => "101111101010001100011010",
25785 => "101100001000001010010010",
25786 => "101000001110011010110010",
25787 => "100100010110011011111000",
25788 => "100100101011110100111111",
25789 => "101001000001001010000000",
25790 => "101100011100100110110000",
25791 => "101101000110111101011100",
25792 => "101101010001011101110000",
25793 => "101111000001011101110110",
25794 => "110010111111011011001100",
25795 => "110111000110110100101101",
25796 => "111001011100111111010000",
25797 => "111011011110000100011011",
25798 => "111101111101001101000111",
25799 => "000000100100001100100111",
25800 => "000011000100100011001001",
25801 => "000100101001001101100101",
25802 => "000110000000011001010010",
25803 => "001000010011011011111100",
25804 => "001010010000011100111111",
25805 => "001001011010101001010110",
25806 => "000110001001001011110010",
25807 => "000010100101010010011011",
25808 => "111110001111001100110011",
25809 => "111010011001010100000001",
25810 => "111001100100000100011001",
25811 => "111010000001010100001001",
25812 => "111011011110011100001000",
25813 => "111111110110101001010111",
25814 => "000110010000101010100100",
25815 => "001010111000011011000100",
25816 => "001010100010111110000010",
25817 => "000111010001111100010100",
25818 => "000100110011010110010100",
25819 => "000011111110100101001110",
25820 => "000011000110110101111100",
25821 => "000000100011000101010001",
25822 => "111110100111111010100000",
25823 => "111110101111101101000111",
25824 => "111110011000110100000010",
25825 => "111100101100011001010010",
25826 => "111011011101110010011000",
25827 => "111101001010111100100000",
25828 => "000010010100001001001000",
25829 => "000111111011100011110110",
25830 => "001010100001000101100111",
25831 => "001001101001110111010011",
25832 => "000111000110011101001101",
25833 => "000011001101110111100111",
25834 => "111110001100011001100000",
25835 => "111000010011011101000100",
25836 => "110001111000100011011110",
25837 => "101101101110011011101010",
25838 => "101100100011100010100010",
25839 => "101011110110001101000000",
25840 => "101010111010010000011010",
25841 => "101011001001010010110110",
25842 => "101101111001101010001010",
25843 => "110010101100100101010110",
25844 => "111000011000101101010011",
25845 => "111110010001000001011101",
25846 => "000011111000101101101011",
25847 => "001001101111110100110000",
25848 => "001110001000110011111110",
25849 => "001110001110000110111000",
25850 => "001011100100000011101100",
25851 => "001001011101111110011100",
25852 => "001000001101001101011110",
25853 => "000110001010110100100000",
25854 => "000011010100111010110100",
25855 => "000001011101011010000101",
25856 => "000000110000000110101101",
25857 => "111111011001001001110000",
25858 => "111101010010100100000010",
25859 => "111011111101111101100110",
25860 => "111011101111001101100011",
25861 => "111100110100110001110011",
25862 => "111110111010111001010001",
25863 => "000000000101100100101000",
25864 => "111111110111111111000010",
25865 => "111111010101100110010011",
25866 => "111110111010010101101100",
25867 => "111110011000001101110110",
25868 => "111101110100001111001111",
25869 => "111110000100001001011101",
25870 => "111110111010011001100100",
25871 => "111111011100010110000110",
25872 => "111111101001000111100110",
25873 => "111111110001010001100000",
25874 => "000000001100011001000100",
25875 => "000001000101011000111001",
25876 => "000001111011101110101000",
25877 => "000010010001110110110000",
25878 => "000010010011001010010100",
25879 => "000001100001111100010100",
25880 => "111110111010010011000011",
25881 => "111011001001011010010001",
25882 => "111000001111010000111010",
25883 => "110111101101101110000001",
25884 => "111000111010100111011000",
25885 => "111001110010111100000111",
25886 => "111010101111101000010101",
25887 => "111101000110100001000011",
25888 => "000000100111100110000101",
25889 => "000100010101010111110101",
25890 => "000111111011101001100010",
25891 => "001100010001100101000110",
25892 => "010000111101001011111000",
25893 => "010100011110111000101100",
25894 => "010110001101101011111000",
25895 => "010110101001001101010000",
25896 => "010111000100000110000000",
25897 => "010110100111011010011100",
25898 => "010100000101100001110100",
25899 => "010001000011111111111010",
25900 => "001110111010010011000000",
25901 => "001100111110001011110000",
25902 => "001001111111001011110000",
25903 => "000110110101000010001101",
25904 => "000101101100001100111011",
25905 => "000110101011000001100110",
25906 => "000111011101110100001010",
25907 => "000101100110000100101011",
25908 => "000010001000001001010001",
25909 => "111111001101011111001000",
25910 => "111100101010110111111000",
25911 => "111010110001000100010101",
25912 => "111001110000010000000100",
25913 => "111001010111100111101010",
25914 => "111001101011110000100011",
25915 => "111011000010011111101010",
25916 => "111101111111001111000011",
25917 => "000001011001000011101111",
25918 => "000100000001010000110010",
25919 => "000101101011110011100100",
25920 => "000110100110110010110100",
25921 => "000111001011000110010010",
25922 => "000110000001010000000000",
25923 => "000011010111101101100011",
25924 => "000000001101011110011110",
25925 => "111010000101110000110100",
25926 => "110000011010111111010010",
25927 => "100110110001111100000101",
25928 => "100001110000011110000100",
25929 => "100001101110101001010001",
25930 => "100001111100000101011001",
25931 => "100010011110010001011000",
25932 => "100111001000010110101001",
25933 => "101110010011111101101110",
25934 => "110100111101011110110101",
25935 => "111010010100111111011110",
25936 => "111101110101111101000101",
25937 => "000000010011010101101101",
25938 => "000011011110010000011101",
25939 => "000110111100110000011100",
25940 => "001001011011000100011100",
25941 => "001010110100100100000110",
25942 => "001010110011110111001000",
25943 => "001000111011100000011010",
25944 => "000110111111100110101010",
25945 => "000111011110111010100110",
25946 => "001001111110111001000101",
25947 => "001100111100101111100010",
25948 => "001111001011101011000100",
25949 => "001110101010111010110000",
25950 => "001011010010100001101010",
25951 => "000110111000010000000010",
25952 => "000010010111000100111110",
25953 => "111101111100011010110000",
25954 => "111010011010110101000001",
25955 => "111001110010100111111111",
25956 => "111011111001001010010010",
25957 => "111111000001111011110111",
25958 => "000100000100011110111110",
25959 => "001001010010111000111110",
25960 => "001010101001100100110000",
25961 => "001000111101100101111100",
25962 => "000111000001110000011001",
25963 => "000101111101000100101010",
25964 => "000101101110111000100100",
25965 => "000011111110111100001101",
25966 => "111110110011110001111001",
25967 => "111000010001110101100110",
25968 => "110010010110010000100000",
25969 => "101100101010101000010000",
25970 => "100111110110101000100100",
25971 => "100101101111100010101000",
25972 => "100111100011000000010001",
25973 => "101100101000001101000000",
25974 => "110010100110101000010110",
25975 => "110111000001011100110100",
25976 => "111001011101111101011001",
25977 => "111011101111111010011010",
25978 => "111101111101111101001011",
25979 => "111110111100000111010101",
25980 => "111110010010001011001010",
25981 => "111011000101010111111110",
25982 => "110111001000011001010111",
25983 => "110100011101000100111010",
25984 => "110000101101100110000110",
25985 => "101100000111011110101010",
25986 => "101010111101001101011000",
25987 => "101110110010000110101010",
25988 => "110101100010001011111000",
25989 => "111101010000010110000000",
25990 => "000100010100001011100110",
25991 => "001001111010000001100000",
25992 => "001111100100010010001000",
25993 => "010011010011110101000100",
25994 => "010001101111011011111110",
25995 => "001101110011011001010100",
25996 => "001011001001000100000011",
25997 => "001010000000010010100001",
25998 => "001000000101100110011101",
25999 => "000011111001010000101000",
26000 => "000000100110000101001010",
26001 => "111111101101000011001101",
26002 => "111111110001110100110100",
26003 => "000000001111001011110111",
26004 => "000000011101011010111101",
26005 => "000000101111010001000010",
26006 => "000001100101100011010111",
26007 => "000010011100110111110000",
26008 => "000001101010000000101110",
26009 => "111110111110111010111110",
26010 => "111101001011010001100111",
26011 => "111100011011111010000010",
26012 => "111011000110000000110100",
26013 => "111000110010111000010010",
26014 => "110101101000101110110101",
26015 => "110010011110110110101100",
26016 => "101111100000011101011000",
26017 => "101110000000011011010010",
26018 => "101110101100111101101100",
26019 => "101111001000001010011000",
26020 => "110000000111001110000110",
26021 => "110010101001001001001100",
26022 => "110011111010010010100110",
26023 => "110011110011101000001110",
26024 => "110011110010110000110110",
26025 => "110100000101010011110110",
26026 => "110100111011101010101011",
26027 => "110110010111010001101101",
26028 => "111000000100000101011111",
26029 => "111001011000001010000101",
26030 => "111010100100111110110111",
26031 => "111100100001111101110001",
26032 => "111111000000000110010000",
26033 => "000001100100110011000111",
26034 => "000100001000110011101000",
26035 => "000111010100101111000010",
26036 => "001011010010000110010101",
26037 => "001110100110110111010100",
26038 => "010001001101011100100000",
26039 => "010011010000000110111010",
26040 => "010100011001111100011010",
26041 => "010101110111010110101010",
26042 => "010111101011010000011010",
26043 => "011000111110010001010011",
26044 => "011001011100011001110001",
26045 => "011001010100100111100001",
26046 => "011010010000000010011111",
26047 => "011011011011001000001101",
26048 => "011011011010001011000101",
26049 => "011011100000001100100001",
26050 => "011011100101011110011110",
26051 => "011011010110111011011111",
26052 => "011011001110001110010100",
26053 => "011010111000010001011100",
26054 => "011001101010011000110011",
26055 => "010110010101111100000100",
26056 => "010001111111011101110000",
26057 => "001101101100010111000010",
26058 => "001001101001110000100100",
26059 => "000111101000001110110110",
26060 => "000111110011111110011001",
26061 => "001001100101111110001010",
26062 => "001011000000110011100010",
26063 => "001010101000110110011011",
26064 => "001010001000110011101100",
26065 => "001001010100000011110010",
26066 => "001000100101001110100010",
26067 => "000110110101110011111111",
26068 => "000001100010101001110001",
26069 => "111001100100001101111100",
26070 => "101101010001101000000000",
26071 => "100010011100111010000101",
26072 => "100001011100011100001001",
26073 => "100010101010101111010110",
26074 => "100001111011011010111111",
26075 => "100010000010110010010011",
26076 => "100010001010110011100100",
26077 => "100110101000110111101111",
26078 => "101111110010101111110100",
26079 => "110111110111110001101001",
26080 => "111111000010101011001011",
26081 => "000110001110101110110010",
26082 => "001011111010000010011100",
26083 => "001111001001111000010110",
26084 => "010000110100100001000000",
26085 => "010001101101110000110100",
26086 => "001111110101001100011110",
26087 => "001001011100000010111010",
26088 => "000000001110110111000011",
26089 => "111001001010110010010001",
26090 => "110110111000010110101001",
26091 => "110110111100101011010100",
26092 => "110111111100010011001110",
26093 => "111000110111000010111000",
26094 => "111000001011011010110001",
26095 => "110111001101101000010000",
26096 => "110111110110110000111000",
26097 => "111010110101110111010100",
26098 => "111110010100000010010111",
26099 => "000000011001101101101110",
26100 => "000100000111101111101010",
26101 => "001010011111110000100010",
26102 => "010000000001011111001110",
26103 => "010011010101110110011100",
26104 => "010100111001001001110100",
26105 => "010100110001000111000010",
26106 => "010011011101011011001000",
26107 => "010011000110001101010110",
26108 => "010011110011100110000010",
26109 => "010010001111010000010010",
26110 => "001110011011001111101100",
26111 => "001000000011111101011110",
26112 => "111101010001010011111011",
26113 => "110001101011011101011000",
26114 => "101000000010001100011000",
26115 => "100001111101110111010101",
26116 => "100001000101000110111000",
26117 => "100001101011001001111001",
26118 => "100100000001011110011111",
26119 => "101010100110000000001000",
26120 => "110001011010100100001010",
26121 => "110110101100100001000111",
26122 => "111100111101001001010000",
26123 => "000101000011001011100000",
26124 => "001011110001100111111000",
26125 => "001101011010110010011110",
26126 => "001010100000100010010110",
26127 => "000011111111110001000110",
26128 => "111010100001100111010101",
26129 => "110000100001001111111000",
26130 => "101000001010100110010100",
26131 => "100011010111011100001011",
26132 => "100011000101100100000001",
26133 => "100110101011101101100011",
26134 => "101100110100110110000110",
26135 => "110100000011011001110000",
26136 => "111010011101111100011001",
26137 => "111110101011001011011110",
26138 => "000001111100000010111000",
26139 => "000100100101010100000100",
26140 => "000100101100001010111100",
26141 => "000011001011011011110100",
26142 => "000010110111011110100011",
26143 => "000011111111101110111011",
26144 => "000100011000011111111100",
26145 => "000011100110100010110000",
26146 => "000011010111011010100011",
26147 => "000011101101010000111010",
26148 => "000011101011001100010111",
26149 => "000011000101011100001101",
26150 => "000010001101010111000101",
26151 => "000001100011101100111001",
26152 => "000001001011010111010110",
26153 => "000000101100000111110010",
26154 => "000000001001011110100110",
26155 => "000000010001000011011011",
26156 => "000000101111001001001010",
26157 => "000000010100001010101001",
26158 => "111110010101101010000001",
26159 => "111010100101111000110100",
26160 => "110110010100100110101110",
26161 => "110010100010110100001110",
26162 => "101110111110100100101110",
26163 => "101100100010001100111100",
26164 => "101011100011010110001000",
26165 => "101011011110111111101000",
26166 => "101100001111001011101110",
26167 => "101101000000110101110110",
26168 => "101110000101011111101000",
26169 => "110000110010110111011000",
26170 => "110100101111010000000111",
26171 => "111000000110010110011110",
26172 => "111001011111000110001010",
26173 => "111001001101011010101110",
26174 => "111000111100111111001111",
26175 => "111001010111011000101010",
26176 => "111001100100111001000000",
26177 => "111010000000010011111001",
26178 => "111011011100001100001101",
26179 => "111100110000111100011101",
26180 => "111101101000111010100101",
26181 => "111110100010010111001010",
26182 => "111110111001111010010110",
26183 => "111110110110110111110110",
26184 => "111111011100101001010101",
26185 => "000001010010111111000100",
26186 => "000011110110100101100101",
26187 => "000101111010111001000110",
26188 => "000111010111001101000001",
26189 => "001000110000010001000110",
26190 => "001001111111100101100000",
26191 => "001011001110001100000010",
26192 => "001101011111111010100110",
26193 => "010001011110010000110010",
26194 => "010110010100110000110100",
26195 => "011001011110101001110111",
26196 => "011001100011101010111000",
26197 => "011000101000000111010001",
26198 => "010111100000101111000100",
26199 => "010100101101101000110110",
26200 => "010000101001101101000110",
26201 => "001101001100110010101000",
26202 => "001011001100111111010110",
26203 => "001010000001110111000010",
26204 => "001001010111000010000101",
26205 => "001001101111111110110100",
26206 => "001011000110111100110010",
26207 => "001100111011001011111110",
26208 => "001110010101110110011000",
26209 => "001111001000010001100110",
26210 => "001111111111111010001000",
26211 => "010000011101100101110110",
26212 => "001111100101011101010000",
26213 => "001100100010110011010010",
26214 => "000110000010011101111110",
26215 => "111101000001011100100111",
26216 => "110101101011111011010100",
26217 => "110010001001000001001110",
26218 => "110000101011000111111110",
26219 => "110001100111111001001110",
26220 => "110110001101101110010111",
26221 => "111100000111111110100110",
26222 => "000000101001101110100010",
26223 => "000010011101111001110101",
26224 => "000010011001100101111101",
26225 => "000011011110110101010110",
26226 => "000110011001000011011011",
26227 => "001000111010111100101000",
26228 => "001001101001001001101111",
26229 => "001000111110111110001010",
26230 => "000110110110111100001110",
26231 => "000001110010001100111000",
26232 => "111001111111111011010100",
26233 => "110001111100101110100100",
26234 => "101011100001111011010110",
26235 => "100111110100100110010101",
26236 => "101000000101110010011110",
26237 => "101011100110011000110110",
26238 => "101111011100011111001010",
26239 => "110010110110001011101000",
26240 => "110110011101010111000100",
26241 => "111010011011101000010000",
26242 => "111111010110111011111101",
26243 => "000100100010001110110101",
26244 => "001000100110111101100010",
26245 => "001100011011100010111100",
26246 => "010000101110000000011000",
26247 => "010010100000110100000010",
26248 => "001111010110001100101010",
26249 => "001001110011000111101000",
26250 => "000100101010001000011111",
26251 => "000001010011001001001110",
26252 => "000000001110001111011110",
26253 => "111110101100110011100011",
26254 => "111100000111110101101100",
26255 => "111010100011111010000010",
26256 => "111000101001110110010101",
26257 => "110100010000010111111001",
26258 => "101111000001010010010000",
26259 => "101101100101100010110010",
26260 => "110001001000000010010110",
26261 => "110101111100010011001001",
26262 => "111010010001011100101011",
26263 => "111110010101110010110111",
26264 => "000011001011000100001100",
26265 => "001001011001000011010000",
26266 => "001110000110111010111000",
26267 => "010000110101011111101010",
26268 => "010011101000100011111000",
26269 => "010100111011011111010110",
26270 => "010011100010001101100100",
26271 => "001111111001110000111010",
26272 => "001001011100011011001111",
26273 => "000001010010101101111001",
26274 => "111010100101011110010000",
26275 => "110110110000110011100010",
26276 => "110100110010010001000000",
26277 => "110100110011101100010000",
26278 => "110111110111110010000100",
26279 => "111100100110111000001011",
26280 => "000001110100111001010011",
26281 => "000110101100110000111000",
26282 => "001001101100011110001010",
26283 => "001011111010010011100100",
26284 => "001110011010111100110110",
26285 => "001111011000011011100010",
26286 => "001110010010111000100100",
26287 => "001101110101010100001010",
26288 => "001110111111110111001110",
26289 => "001110100011010100011000",
26290 => "001011001011111000001100",
26291 => "000110111110110110101111",
26292 => "000011010011110010110000",
26293 => "000000110101111111100010",
26294 => "111101110101000110111001",
26295 => "111000111110011001111100",
26296 => "110100101011101000000001",
26297 => "110010010011111011011010",
26298 => "110010011110010010001000",
26299 => "110100101000010110100100",
26300 => "110110111010010000000010",
26301 => "111001100011000001100011",
26302 => "111011100011110010011000",
26303 => "111011001100110100100000",
26304 => "111000010001101110001100",
26305 => "110011011000010100111000",
26306 => "101110001011110111001000",
26307 => "101000100001110100101100",
26308 => "100100000010000111011111",
26309 => "100011110001111000100011",
26310 => "100101001101111101111001",
26311 => "100110110001000000011101",
26312 => "101001001001100110101110",
26313 => "101011100100010011110010",
26314 => "101111110010010101000100",
26315 => "110110001010110001001100",
26316 => "111011100111010100001011",
26317 => "111110111111010100010100",
26318 => "000001010000000011001100",
26319 => "000011001110111011011101",
26320 => "000100001000101000100110",
26321 => "000011001001001000111011",
26322 => "000001000001011110101100",
26323 => "111110101011101100011110",
26324 => "111100101011010011000101",
26325 => "111010110011010111001001",
26326 => "111001001010001001110111",
26327 => "111000010101100010010000",
26328 => "111000000010110010011001",
26329 => "111000100010010100111010",
26330 => "111011001000111101011000",
26331 => "000000100101010011111011",
26332 => "000110110000010110000100",
26333 => "001010011111111001100101",
26334 => "001100111100001011100010",
26335 => "010000001001110110100110",
26336 => "010010110001101111011000",
26337 => "010100010101111011010000",
26338 => "010110000100100100111100",
26339 => "010111010010100001011010",
26340 => "010101111110100010100100",
26341 => "010010000000000010000000",
26342 => "001101011010101000001010",
26343 => "001001010101011101010101",
26344 => "000101010111100000000110",
26345 => "000000111010010001110001",
26346 => "111100001101010101011010",
26347 => "111001010101110100100101",
26348 => "111001001001111011001000",
26349 => "111001110111011010011011",
26350 => "111010110101000011100110",
26351 => "111101001110110001100111",
26352 => "000001011110001010110100",
26353 => "000101010010100101001001",
26354 => "000110001111110111111101",
26355 => "000101111100110001000110",
26356 => "000110111100000001011110",
26357 => "000111011110101101110111",
26358 => "000011100000010101101100",
26359 => "111011000001101100000010",
26360 => "110011000110100110101000",
26361 => "101110111000110110110110",
26362 => "101101011111111101111000",
26363 => "101101111011110111100010",
26364 => "110000100010111000010100",
26365 => "110101111110100011001010",
26366 => "111100001110010011100100",
26367 => "000000010000000011100111",
26368 => "000010110100110001111000",
26369 => "000110010000111000101001",
26370 => "001010111000110100010110",
26371 => "001111110110110100111010",
26372 => "010100010100010110010010",
26373 => "010110111100001010110010",
26374 => "010110100011111101001000",
26375 => "010011111110110111001000",
26376 => "010000010100101101011000",
26377 => "001011110111111000010000",
26378 => "000110110111001010011111",
26379 => "000001010100010000011010",
26380 => "111100110111111000100000",
26381 => "111011010100101011111000",
26382 => "111011000101011011001100",
26383 => "111010010000110111111011",
26384 => "111010000100111000001101",
26385 => "111100101011000101011010",
26386 => "000001001011100011010010",
26387 => "000100100110110110111011",
26388 => "000110101110010110101101",
26389 => "001001110001100100110101",
26390 => "001101111110001110010010",
26391 => "010000100001001101010100",
26392 => "001110101111101100110110",
26393 => "001000100101001001101100",
26394 => "000000101001011111101000",
26395 => "111010010100111110101010",
26396 => "110101101110000011010100",
26397 => "110000111100011011111010",
26398 => "101101000101010001010010",
26399 => "101011100010011011100010",
26400 => "101011000001101101010100",
26401 => "101010010000001101101100",
26402 => "101001000010100101010010",
26403 => "101000110011111110101100",
26404 => "101100001011000110001110",
26405 => "110010100110000011010010",
26406 => "111000100111000110001000",
26407 => "111100111110111111101111",
26408 => "000000000000101100101010",
26409 => "000001101101111010111101",
26410 => "000011110101011001010000",
26411 => "000110101100111001010011",
26412 => "000110110110000000010111",
26413 => "000011011011100000001001",
26414 => "000000010001000000001101",
26415 => "111110110100101100010100",
26416 => "111100010101101110111101",
26417 => "110111000000000011011000",
26418 => "110001000101010110110010",
26419 => "101110101111010011010000",
26420 => "110000101111100101011100",
26421 => "110100010001101100000001",
26422 => "111000101010110011000110",
26423 => "111111011011111110011101",
26424 => "000111100011010100000100",
26425 => "001110010100101010011100",
26426 => "010010101101000010001100",
26427 => "010100101111111101001110",
26428 => "010101000111111111101010",
26429 => "010101101100011010110000",
26430 => "010110000101110100011110",
26431 => "010011100111010001001100",
26432 => "001111111110011110111010",
26433 => "001111010111110010001010",
26434 => "010000101010101001001000",
26435 => "001111110111100010101110",
26436 => "001100001111011100011110",
26437 => "001000011100000100001010",
26438 => "000110101100100000010101",
26439 => "000101011010011110010100",
26440 => "000001110010100010010000",
26441 => "111100100101000010000110",
26442 => "111000100010111110101110",
26443 => "110111100011001001001101",
26444 => "111001100011010101111010",
26445 => "111011110011000011110011",
26446 => "111100101101000111011111",
26447 => "111110000110011000100111",
26448 => "111111101011110010011000",
26449 => "111110110111111100111000",
26450 => "111100000011001101100101",
26451 => "111001000011001011011011",
26452 => "110101111000001110101110",
26453 => "110001111111011111101100",
26454 => "101101101010101100111010",
26455 => "101001101000010111010110",
26456 => "100110101110001101011101",
26457 => "100101100011110001010001",
26458 => "100110001101011000010101",
26459 => "101000010111010100010000",
26460 => "101011110011000010010010",
26461 => "110000001101000011110010",
26462 => "110100100001000101001010",
26463 => "110111111011011010111000",
26464 => "111010110111111111111001",
26465 => "111101001100010011100011",
26466 => "111101110000010100010011",
26467 => "111100100111011100101011",
26468 => "111011010010001010100110",
26469 => "111010101000101110100101",
26470 => "111001110001000011100010",
26471 => "111000100110000110001110",
26472 => "111001000011001010111000",
26473 => "111011011010111101101010",
26474 => "111110100010011001100010",
26475 => "000010110010000110000101",
26476 => "000111110100011010000011",
26477 => "001100000011011001001110",
26478 => "010000001010010010111000",
26479 => "010100101110101010001100",
26480 => "010111101000011101110010",
26481 => "011000001000110010101101",
26482 => "010111110000111110100100",
26483 => "010111010000001001001010",
26484 => "010110100011100001110010",
26485 => "010100111110110100100100",
26486 => "010001110111011110101100",
26487 => "001110011110010111000100",
26488 => "001011111111010011111000",
26489 => "001001110111011001110111",
26490 => "001000010111111100001110",
26491 => "001000000000000000100111",
26492 => "000111011001001000101101",
26493 => "000110010011010011000000",
26494 => "000110011101101011110011",
26495 => "001000000100111011001001",
26496 => "001001100111101110011111",
26497 => "001010000011001100110010",
26498 => "001001011110011000001011",
26499 => "001000100100101011100111",
26500 => "000111001011111100010100",
26501 => "000100110010111110010000",
26502 => "000001101000110010100101",
26503 => "111100111100000101101100",
26504 => "110101101110100110001101",
26505 => "101110110100111110111110",
26506 => "101100001110101001011100",
26507 => "101101001010001111111000",
26508 => "101110101011001111111010",
26509 => "110001000000001110000100",
26510 => "110101001110111011011100",
26511 => "111001101011100001101101",
26512 => "111100001111010001110110",
26513 => "111101001101101001000001",
26514 => "111110010111001010010101",
26515 => "000000110101001001000101",
26516 => "000011111010001110110000",
26517 => "000110001110000111101110",
26518 => "000111100110111001010111",
26519 => "000111101010001011010001",
26520 => "000101010011010100010001",
26521 => "000001100000101011001001",
26522 => "111110001000100111000111",
26523 => "111011100100010101100110",
26524 => "111001111111011110110000",
26525 => "111000111101111001110010",
26526 => "110111001110011111000110",
26527 => "110101100110000111001101",
26528 => "110110000011111100000010",
26529 => "111001000000011000011100",
26530 => "111110000100101101000001",
26531 => "000011111100000111000111",
26532 => "001000100101000101011010",
26533 => "001100110100010101011100",
26534 => "010010100101111110101000",
26535 => "010111110001000100101000",
26536 => "011000101110111111000011",
26537 => "010101100010010111001010",
26538 => "010000000100110110001100",
26539 => "001010000001000000101001",
26540 => "000101101010000100100101",
26541 => "000011001011001011101111",
26542 => "000000000100000100001101",
26543 => "111101001001000101100110",
26544 => "111101001001111101110000",
26545 => "111101110110100101010010",
26546 => "111011111000111001110010",
26547 => "111000111101010101011000",
26548 => "111000011011111010000010",
26549 => "111011011001111010011110",
26550 => "111111110100011111101001",
26551 => "000010001100010101111010",
26552 => "000010100010001000110110",
26553 => "000011010010011100000111",
26554 => "000011111000111111110000",
26555 => "000010111101010100111110",
26556 => "000000110010100100110101",
26557 => "111100110000001100111111",
26558 => "110111000011111001001010",
26559 => "110010010000111100100100",
26560 => "101111000000100100001100",
26561 => "101100000100000100001110",
26562 => "101001010100000111010010",
26563 => "100110111010001010011111",
26564 => "100110001000011001100011",
26565 => "101001100000010011110110",
26566 => "110000000011100010111110",
26567 => "110110110111101000001101",
26568 => "111110011011010011100011",
26569 => "000110111011110001000000",
26570 => "001101100010111011010010",
26571 => "010001000010011001011010",
26572 => "010001110010000100001010",
26573 => "001111100010010111111100",
26574 => "001011011111110101111010",
26575 => "000110111000011001111100",
26576 => "000001000011101001000001",
26577 => "111011010000001010011000",
26578 => "111000100000110101001011",
26579 => "111001010100011010011111",
26580 => "111011110001001110011010",
26581 => "111110000011001101010111",
26582 => "111111101011100111000111",
26583 => "000001110111111010000011",
26584 => "000100111101111101010000",
26585 => "000110101011010010000110",
26586 => "000101100010110000001111",
26587 => "000011010010010100010110",
26588 => "000010001100000100100010",
26589 => "000010101111010101110110",
26590 => "000011011010110000101001",
26591 => "000010100001001001100001",
26592 => "000001001000000010000100",
26593 => "000000110101000100001111",
26594 => "111111101101001011101101",
26595 => "111100101011111011100011",
26596 => "111010011110010110111110",
26597 => "111001011001011111000100",
26598 => "110111000101111011000100",
26599 => "110100000010001011000110",
26600 => "110001101000110110101000",
26601 => "101111111000001100000100",
26602 => "101111011000010101111010",
26603 => "110000010010001100100010",
26604 => "110001010111001011010100",
26605 => "110010011011110111110110",
26606 => "110100010000111100111010",
26607 => "110111010010011100011100",
26608 => "111011011010011011101000",
26609 => "111111010110010011110010",
26610 => "000001100011011000111110",
26611 => "000001111111101110110011",
26612 => "000001100100101100101100",
26613 => "000001000000010111110000",
26614 => "000000011011000101010000",
26615 => "111110111100000010110001",
26616 => "111011111110101101101100",
26617 => "111001001010111101111111",
26618 => "111000001111101000011000",
26619 => "111000001101110010101100",
26620 => "110111110111100001100110",
26621 => "111000010101001100111110",
26622 => "111010110110101111100010",
26623 => "111111010000101101011101",
26624 => "000100011000111110110111",
26625 => "001000100100000110111010",
26626 => "001011110001011110100000",
26627 => "001111010011111111001000",
26628 => "010010000110100100101110",
26629 => "010010011110101011001110",
26630 => "010001101011011100100100",
26631 => "010000101110011110110110",
26632 => "001110011111101110011010",
26633 => "001011000111000101010111",
26634 => "001000010110101001110100",
26635 => "000110110001011010011100",
26636 => "000101100011111101110010",
26637 => "000100001101101000011110",
26638 => "000011001111111111001100",
26639 => "000100000101000011011011",
26640 => "000110110001101110101110",
26641 => "001000110010001000011101",
26642 => "001000110010110010111110",
26643 => "001000101010000100100010",
26644 => "001000110011011110010010",
26645 => "000111011000011100001000",
26646 => "000100001000001001101110",
26647 => "111111111101101110010101",
26648 => "111010111111000001001000",
26649 => "110101001011110011100011",
26650 => "101111010101011110011100",
26651 => "101011010001011000001100",
26652 => "101010111010010111000000",
26653 => "101110011000110110100110",
26654 => "110011110111110101011000",
26655 => "111000111011001001010100",
26656 => "111100100000111011010011",
26657 => "111111000000101110000101",
26658 => "111111111010101110001011",
26659 => "111111011110101011100000",
26660 => "000000000110100101010111",
26661 => "000010000011110100100100",
26662 => "000011100010010111001010",
26663 => "000100110011111111100111",
26664 => "000110010100010011011110",
26665 => "000110100101101011101101",
26666 => "000100100110010000000000",
26667 => "000000111001001011010101",
26668 => "111101101110101001110110",
26669 => "111100111111110011000110",
26670 => "111100101111100001011101",
26671 => "111001110010111100011010",
26672 => "110100110101011100100100",
26673 => "110001001100100111011110",
26674 => "110000100000011010111010",
26675 => "110001101001110101011000",
26676 => "110011110010010000000010",
26677 => "110111101001010010000111",
26678 => "111100111010010111100111",
26679 => "000010000011110100110010",
26680 => "000110011010100011000100",
26681 => "001001001000010111101001",
26682 => "001001001111011000000100",
26683 => "000111100000011110011010",
26684 => "000101001110110001010010",
26685 => "000011100010001111110000",
26686 => "000100000100110100110010",
26687 => "000110101010110110111000",
26688 => "001000101001101100111101",
26689 => "001000110011001110011110",
26690 => "000111101100100101111101",
26691 => "000100111011100100111101",
26692 => "000001000111111010001011",
26693 => "111111100111011101100111",
26694 => "000001101001101111001111",
26695 => "000100001001110001000101",
26696 => "000100011110111000000010",
26697 => "000011100111000110101010",
26698 => "000100001011111011001111",
26699 => "000110101001111010101010",
26700 => "001000010110111000101110",
26701 => "001000101010111011101011",
26702 => "001010110000010111010111",
26703 => "001110101111101010010110",
26704 => "010000101000110010100100",
26705 => "001111010100010110010010",
26706 => "001100110001100010001110",
26707 => "001001100111111111000111",
26708 => "000110000100011000011001",
26709 => "000011010011100000001000",
26710 => "000010010001011001110101",
26711 => "000011110000100110111111",
26712 => "000111100100110100000001",
26713 => "001011010000110100011010",
26714 => "001101010111111101001110",
26715 => "001111000111110000111000",
26716 => "010000011100100111101000",
26717 => "010000000100110110011000",
26718 => "001110010111111010011010",
26719 => "001011000101000000011110",
26720 => "000101010011001011011000",
26721 => "111110110001101000010110",
26722 => "111001001011100010010110",
26723 => "110100011101000010010011",
26724 => "110001111011110011011100",
26725 => "110010101001010000001100",
26726 => "110101001100000110001111",
26727 => "111000101101111100001000",
26728 => "111101001101101100010011",
26729 => "000001110101011010010111",
26730 => "000101001111000001001110",
26731 => "000101111010010001010110",
26732 => "000011110100111111110100",
26733 => "000000110101111011001101",
26734 => "111101111011000000101100",
26735 => "111011000101110110001110",
26736 => "111000100101100100011100",
26737 => "110101110111100111011110",
26738 => "110010011010011101001010",
26739 => "101110101100011110110100",
26740 => "101011010010100001011110",
26741 => "101000110010011100111010",
26742 => "100111100100111000000111",
26743 => "100111100011111000011100",
26744 => "101000100010110001111110",
26745 => "101001110100101010100000",
26746 => "101011001111110000011110",
26747 => "101101111111011100001000",
26748 => "110010000000100101111100",
26749 => "110101110101010010011010",
26750 => "111001001000100100010011",
26751 => "111100010001101010100100",
26752 => "111110111111001010111011",
26753 => "000000101110001111111000",
26754 => "000001010000000000011000",
26755 => "000000110000000101000110",
26756 => "111111010011011000010101",
26757 => "111101101001001010111100",
26758 => "111101110111101101111001",
26759 => "000000011011101100100001",
26760 => "000010100100001001010111",
26761 => "000010000110011100010010",
26762 => "000000011110000001010101",
26763 => "000000101001010011101011",
26764 => "000010111001101001001001",
26765 => "000100101011110011100100",
26766 => "000101011011010011001111",
26767 => "000111010101101111000111",
26768 => "001011000101111001110100",
26769 => "001111001000010011010100",
26770 => "010010001111101000000000",
26771 => "010100001100110111000110",
26772 => "010101010110011010010000",
26773 => "010110010000110110111000",
26774 => "010110110011011001000000",
26775 => "010110000110010110101100",
26776 => "010100000011001011001010",
26777 => "010001001001101101101010",
26778 => "001100111100110001011100",
26779 => "000111100111010001011111",
26780 => "000010110110111000000010",
26781 => "111110111001000000001100",
26782 => "111010111010100110110110",
26783 => "110111110110000001011000",
26784 => "110110101100011100000100",
26785 => "110111101001111111110011",
26786 => "111010010110001001010101",
26787 => "111100111000100011011010",
26788 => "111110011011010110110000",
26789 => "000000010111100011000110",
26790 => "000010011001010110010010",
26791 => "000010100110101010011100",
26792 => "000001000011001000011000",
26793 => "111111001011100010000110",
26794 => "111100111011011000101111",
26795 => "111000011010011011101011",
26796 => "110001101001001011011000",
26797 => "101100001011001100110000",
26798 => "101010101110110111011100",
26799 => "101100100001001100101000",
26800 => "101111010111001011000110",
26801 => "110010000111001110011010",
26802 => "110101010010001111111001",
26803 => "111000100010001111101001",
26804 => "111001110110111011111100",
26805 => "111001100100011111010101",
26806 => "111001111110111000011001",
26807 => "111011101011100010111000",
26808 => "111110001011101000100101",
26809 => "000000101111000001111001",
26810 => "000010010110011111010111",
26811 => "000011000000111001111010",
26812 => "000010010110010110100100",
26813 => "111111100100110000001100",
26814 => "111100011000001111010100",
26815 => "111011000110100010000100",
26816 => "111010100111010010000011",
26817 => "111000011010010100011001",
26818 => "110101100101011100100110",
26819 => "110101001010001110110010",
26820 => "110110101011110001000110",
26821 => "111000000000000001100000",
26822 => "111001010111111000010010",
26823 => "111011011011101011110010",
26824 => "111110010010000001101001",
26825 => "000010011000101110101110",
26826 => "000110000101101111101100",
26827 => "000110111100000111101000",
26828 => "000101011100101011111001",
26829 => "000010110011000011111001",
26830 => "111110111111100010101100",
26831 => "111011101011101001111011",
26832 => "111011101010010000110101",
26833 => "111110010111001110010011",
26834 => "000000001100100011110101",
26835 => "111111111001110010010101",
26836 => "111110101001111011111000",
26837 => "111100100010000011010010",
26838 => "111010000010000100100111",
26839 => "111000101001100001011000",
26840 => "111000011100000001111100",
26841 => "111001000101001110111100",
26842 => "111001111001101100010011",
26843 => "111001101000100010100111",
26844 => "111001101010101000010111",
26845 => "111011100000010011100111",
26846 => "111101010111100010101100",
26847 => "111111000110101101101110",
26848 => "000010100100110111000000",
26849 => "000110011100101110011110",
26850 => "001000011010100110101010",
26851 => "001000110000000010111100",
26852 => "001000010011100001100110",
26853 => "000111001000111110101011",
26854 => "000101001001001100001110",
26855 => "000010100101000001101110",
26856 => "000000111101111000110001",
26857 => "000010010110011010000011",
26858 => "000110011001010110001110",
26859 => "001010101000111100000101",
26860 => "001110010001111001010100",
26861 => "010001110111000110001100",
26862 => "010100011100111001111110",
26863 => "010101000001101010100110",
26864 => "010011011101111110111000",
26865 => "010000001011000101000110",
26866 => "001101011000011111000110",
26867 => "001100011111010101011100",
26868 => "001011100001111011010010",
26869 => "001001111111001011000011",
26870 => "001001110001111111101110",
26871 => "001010111000000100111010",
26872 => "001100011001111111000110",
26873 => "001110100011110100110000",
26874 => "010000011011100110000000",
26875 => "010000001110001101111100",
26876 => "001101110000011010111010",
26877 => "001010011000000001011000",
26878 => "000110100011010111011101",
26879 => "000010001000001111101111",
26880 => "111110100110111111010110",
26881 => "111100101000010000011011",
26882 => "111001100111101001010100",
26883 => "110100110100110100011111",
26884 => "110000101001100100110100",
26885 => "101101001110001000100100",
26886 => "101001000100011100001010",
26887 => "100101010110101001101101",
26888 => "100011110011110010010101",
26889 => "100011110011101011101000",
26890 => "100100010010010100001001",
26891 => "100101111000011010010011",
26892 => "101001010111100100000000",
26893 => "101101110100110000111010",
26894 => "110010010001000100101010",
26895 => "110110110110111001110000",
26896 => "111010110101000110110101",
26897 => "111100110100010011111101",
26898 => "111101101111011101000000",
26899 => "111110110110101000100010",
26900 => "111110010110101111001111",
26901 => "111010110010010101100111",
26902 => "110110110101010111101111",
26903 => "110101010100000111010111",
26904 => "110101001000011001100011",
26905 => "110100101110010010110101",
26906 => "110101000110110100111110",
26907 => "110110111011101110000011",
26908 => "111001001011101000100100",
26909 => "111011111010011000101100",
26910 => "111111111101111000110100",
26911 => "000100100111001011100110",
26912 => "001000110110011100010011",
26913 => "001101011110100000101000",
26914 => "010011101101001100111010",
26915 => "011010010101000100101100",
26916 => "011110001101101100110101",
26917 => "011110110101100010000101",
26918 => "011110100111111100001011",
26919 => "011110001100010110010100",
26920 => "011100111100100010010011",
26921 => "011011110100001011110111",
26922 => "011011001000010010010101",
26923 => "011010100110101111001001",
26924 => "011010010011011001010011",
26925 => "011000011100010001100001",
26926 => "010011101010000111101100",
26927 => "001101110101010111100110",
26928 => "001000110100100110111011",
26929 => "000101011010001011001000",
26930 => "000100110111111101100011",
26931 => "000111010101110001010110",
26932 => "001010101110000100110000",
26933 => "001100101101011010100100",
26934 => "001101011101100000110100",
26935 => "001110101011100011001010",
26936 => "001111111001100001010010",
26937 => "010000000111011110111100",
26938 => "010000001011101001000100",
26939 => "001110111111110100000010",
26940 => "001001101111011000001011",
26941 => "000000001101100101100110",
26942 => "110100011111100010011101",
26943 => "101010001110011001111010",
26944 => "100100111011110001110101",
26945 => "100011110101101001001011",
26946 => "100100000011110111000001",
26947 => "100100111101001010111111",
26948 => "100110001000101001100011",
26949 => "100110010011001100010001",
26950 => "100101111000110001011000",
26951 => "100111001110110110010001",
26952 => "101011100100000111101110",
26953 => "110001101000111000100010",
26954 => "110111101001010110100010",
26955 => "111100011110101001111011",
26956 => "111111011101011101001000",
26957 => "000000101000001101100101",
26958 => "111111111110111111000101",
26959 => "111101011100010101000010",
26960 => "111010100101001010011100",
26961 => "111000111000110100000010",
26962 => "110111101010001011111000",
26963 => "110110100010101000000011",
26964 => "110110001110000000110001",
26965 => "110101111110001111100111",
26966 => "110100110010011111000110",
26967 => "110100000111001011101111",
26968 => "110110000001001010011011",
26969 => "111001011100111100001000",
26970 => "111011111000011000010000",
26971 => "111101100100001101011101",
26972 => "000000000110000000100011",
26973 => "000010100000011011110111",
26974 => "000010001101010101100100",
26975 => "111110011101100110110010",
26976 => "111010001000100000100110",
26977 => "111001101010001001001100",
26978 => "111110010111011010010010",
26979 => "000100110110001001101011",
26980 => "001001000000101001011010",
26981 => "001010001100010100100100",
26982 => "001001100001101001111101",
26983 => "000110111101000000010010",
26984 => "000010110000111100101001",
26985 => "111110010101111100110010",
26986 => "111010011010110010000101",
26987 => "111000000010011100001100",
26988 => "110111110110000010010100",
26989 => "110111101111110111110110",
26990 => "110110000000110101011000",
26991 => "110011101100100101111100",
26992 => "110011000001000001011000",
26993 => "110101111110000111000100",
26994 => "111011000101101100010100",
26995 => "111110000100010100011110",
26996 => "111110110010010110010110",
26997 => "000000000011000000101000",
26998 => "000000110100110111011101",
26999 => "111110100001010000011000",
27000 => "111001100111111000000001",
27001 => "110101010110010111000010",
27002 => "110100111111011110110000",
27003 => "111000010011101111011101",
27004 => "111011110111010010001000",
27005 => "111110010000001000100001",
27006 => "000001001110011001000000",
27007 => "000101011100100011100011",
27008 => "001000110000010000011100",
27009 => "001001010110010010001010",
27010 => "001000011000011001011011",
27011 => "000111111111101110001001",
27012 => "001000100001111100100110",
27013 => "001000100110111001110100",
27014 => "000111000111100001000000",
27015 => "000101001111000111101111",
27016 => "000101011000001111001001",
27017 => "000111101000001010000010",
27018 => "001001110011111100110111",
27019 => "001010111010001001010101",
27020 => "001011110010111010101000",
27021 => "001101001000111100010010",
27022 => "001101111010100001101000",
27023 => "001100100000011010011010",
27024 => "001001011110100000001010",
27025 => "000111011000011101010001",
27026 => "000111000000101010110111",
27027 => "000110101001101101010001",
27028 => "000101011101101001111001",
27029 => "000100010000001100110000",
27030 => "000011100011101100000101",
27031 => "000010110111111100101101",
27032 => "000000110011000111000101",
27033 => "111101000100100111000011",
27034 => "111010000100101010111110",
27035 => "111000111101100111110010",
27036 => "110111111011010010101110",
27037 => "110110011101010011111111",
27038 => "110101110010000010101110",
27039 => "110110001001011111101010",
27040 => "110111001101011110000111",
27041 => "111000000110000110010000",
27042 => "111000001000111000011110",
27043 => "111000011011011111100101",
27044 => "111000111011001010010110",
27045 => "110111010111001000111011",
27046 => "110011101010011011010100",
27047 => "101111111101101000011110",
27048 => "101100110010011010011000",
27049 => "101001110110001000011010",
27050 => "101000010000011111100000",
27051 => "101000111111010001100000",
27052 => "101011001110011110000000",
27053 => "101110000111011011100110",
27054 => "110010010111010101010110",
27055 => "111000110011101110000001",
27056 => "000000011111001100010100",
27057 => "000111010001100001111100",
27058 => "001100100001111000010100",
27059 => "010001010111010110110010",
27060 => "010101101000101001000010",
27061 => "011000001011110000101100",
27062 => "011001001011101011100001",
27063 => "011000010101110110000101",
27064 => "010100110111110000110110",
27065 => "010000110001010110111100",
27066 => "001110010000011100110000",
27067 => "001100000100001101111100",
27068 => "001001001100010100111011",
27069 => "000111100100011011001011",
27070 => "000111110010001001110001",
27071 => "000111010010010101001111",
27072 => "000101100001110011100000",
27073 => "000101011110001110001000",
27074 => "000111101110111110011001",
27075 => "001001110100110000101100",
27076 => "001011101011100000111011",
27077 => "001111000001001000001110",
27078 => "010011001110010011110100",
27079 => "010110011011001100000100",
27080 => "010111101001001110011000",
27081 => "010111000010001010100100",
27082 => "010101011100000001000000",
27083 => "010011000111100010010100",
27084 => "010000010001011001011010",
27085 => "001101110101000010100000",
27086 => "001010100000110100111000",
27087 => "000011000010100000101111",
27088 => "111000010101001111000100",
27089 => "101111100010010001110010",
27090 => "101010111000001111110010",
27091 => "101000110111011111101010",
27092 => "101000101110010001000010",
27093 => "101010110101010000100100",
27094 => "101111001001001010000100",
27095 => "110100000110100011011001",
27096 => "110111010000110100110000",
27097 => "111001001101001011111000",
27098 => "111101001000101011100100",
27099 => "000011010010001000000000",
27100 => "001001010100101101111011",
27101 => "001101111010111010000000",
27102 => "001111111001111110001110",
27103 => "001101111100110110011000",
27104 => "000111101100110010110100",
27105 => "111110011000111010010110",
27106 => "110101011000101111111110",
27107 => "101111010011101001011110",
27108 => "101011000111010110000000",
27109 => "100111010001001110001101",
27110 => "100100110110010001001101",
27111 => "100101100101101011111111",
27112 => "101000111101100011010000",
27113 => "101100110111011111011010",
27114 => "110001001101101101000000",
27115 => "110111100011111100101110",
27116 => "111111010001110001110101",
27117 => "000110000110010101100011",
27118 => "001010011100101110110000",
27119 => "001011010010101010101010",
27120 => "001000101111010110000010",
27121 => "000100000101110100110000",
27122 => "111110110110011010010011",
27123 => "111011100000100000101011",
27124 => "111100001000100110110110",
27125 => "111111000110100000001101",
27126 => "000001010001000111001110",
27127 => "000010010111100010010100",
27128 => "000011100000010100111100",
27129 => "000011110110110011101111",
27130 => "000010100111111011101100",
27131 => "000001011101010010101001",
27132 => "000001110100000100101101",
27133 => "000010100001000011001111",
27134 => "000001101011011010000111",
27135 => "111111001110010110111011",
27136 => "111100110000100100101110",
27137 => "111011001011010111111001",
27138 => "111010001000100100010111",
27139 => "111010100001011110101100",
27140 => "111101100100001001011001",
27141 => "000001100011100010001000",
27142 => "000100001100011010100010",
27143 => "000101101101000010110011",
27144 => "000110011110001111110110",
27145 => "000101100110111101010000",
27146 => "000011000011011000000100",
27147 => "000000010111110100010110",
27148 => "111111101010010101110010",
27149 => "000001100110111111100000",
27150 => "000100010000010010000110",
27151 => "000101101100111110011010",
27152 => "000110110001100111001011",
27153 => "001000001011010111110101",
27154 => "001000011101100100010100",
27155 => "000110111000010110101101",
27156 => "000100011011100101011001",
27157 => "000010010010011000101000",
27158 => "000001001100101100001000",
27159 => "000000011100001111101111",
27160 => "111110100100110111100001",
27161 => "111100011110000000000010",
27162 => "111011111101100101101000",
27163 => "111100011101011001010010",
27164 => "111100010001110001001000",
27165 => "111011100011010100101101",
27166 => "111011111110100010001101",
27167 => "111110000110011110100110",
27168 => "111111110000101010011100",
27169 => "111110110111011010100011",
27170 => "111100010101110001000110",
27171 => "111010010111000110000101",
27172 => "111001111011001111111001",
27173 => "111010110001101101100000",
27174 => "111011110111101001001010",
27175 => "111100101000001010001001",
27176 => "111101101010001100111001",
27177 => "111110100111100000100111",
27178 => "111101101010001100100011",
27179 => "111010110110110010011111",
27180 => "111000010001001111001100",
27181 => "110110010001111100110111",
27182 => "110100010111110010001001",
27183 => "110011011010000100011100",
27184 => "110011110001010110110110",
27185 => "110100100101001101101100",
27186 => "110101010010100100100000",
27187 => "110110000011001111101011",
27188 => "110111100010100100010111",
27189 => "111001101010100011101011",
27190 => "111011001010001000100110",
27191 => "111100010010111100110011",
27192 => "111110011100110101101100",
27193 => "000001000101111111010100",
27194 => "000011000111101100111100",
27195 => "000100011111100101100100",
27196 => "000101001100100111010100",
27197 => "000101001110110111111011",
27198 => "000101001001010100000111",
27199 => "000101110100110011110001",
27200 => "000111100001011010111000",
27201 => "001001000110011001110111",
27202 => "001010000001001111001011",
27203 => "001011011010001100000001",
27204 => "001101100000100001010000",
27205 => "001111001101110100100000",
27206 => "010000100011010011111100",
27207 => "010010010110001100011110",
27208 => "010011011100110000001000",
27209 => "010001001010100010111100",
27210 => "001011100001000110111110",
27211 => "000101110001011001111011",
27212 => "000010000101110101001000",
27213 => "000000001110010011110010",
27214 => "111111010111111110101101",
27215 => "111110111111010000001111",
27216 => "111110111110111110111101",
27217 => "111111101100100010000011",
27218 => "000001110010111101011000",
27219 => "000101010100101110011000",
27220 => "000111111110101010101010",
27221 => "001000011111010101100101",
27222 => "001010000011111010111100",
27223 => "001110011001100110101100",
27224 => "010001110001001101001110",
27225 => "010001100111110110010000",
27226 => "001111101101100010011100",
27227 => "001101000100001101101000",
27228 => "001000100100110000111100",
27229 => "000010110000110111001000",
27230 => "111110010101101111010111",
27231 => "111100000101001100111001",
27232 => "111000111111110111111010",
27233 => "110010001110000010101000",
27234 => "101001010011001010101000",
27235 => "100010110000111001100011",
27236 => "100000111111000001110101",
27237 => "100010110111010001010111",
27238 => "100110101111011100110001",
27239 => "101011111010100100100010",
27240 => "110010001010010001001110",
27241 => "111000100101111100101000",
27242 => "111101001101001110111111",
27243 => "111111110101010010010010",
27244 => "000011001101011100111001",
27245 => "001000010111110111001100",
27246 => "001101010100111111100100",
27247 => "010000110100001101111110",
27248 => "010010110111001110111010",
27249 => "010010100110101010100000",
27250 => "001110101000101011011000",
27251 => "000111100001101101001101",
27252 => "000000001001001001111000",
27253 => "111010011011100011101001",
27254 => "110101111010100001011110",
27255 => "110010000010000101000000",
27256 => "101111101111011100100110",
27257 => "110000000111010000111010",
27258 => "110010010101001011010100",
27259 => "110101000001110001001011",
27260 => "111000110110110111101111",
27261 => "111110101000111100000101",
27262 => "000101011100001101111010",
27263 => "001100000010101110010110",
27264 => "010000111110100011111000",
27265 => "010010110100111110110110",
27266 => "010001001101001111011010",
27267 => "001011010000000001111100",
27268 => "000001101110010100010110",
27269 => "111001111110100001100000",
27270 => "110111100110010001100110",
27271 => "110111100000100001110101",
27272 => "110110100001111000100011",
27273 => "110101110111101100111010",
27274 => "110110011101001110001101",
27275 => "110110111011011111111000",
27276 => "110111001110101000101100",
27277 => "111000010101000111011001",
27278 => "111001111110011111000011",
27279 => "111011110111011010001000",
27280 => "111100111101100010001000",
27281 => "111011011010100000000001",
27282 => "111000011111111010001111",
27283 => "110110010001001000001110",
27284 => "110100000001010001011001",
27285 => "110011000001010111111010",
27286 => "110101100000001010101010",
27287 => "111001000010100001011101",
27288 => "111011010001111011000100",
27289 => "111101010110101101000011",
27290 => "111111001000011101000010",
27291 => "111111011001010110110000",
27292 => "111110100011000110000100",
27293 => "111101100011100111001101",
27294 => "111101111101001100000101",
27295 => "000000111010100110101110",
27296 => "000100100001011010110110",
27297 => "000110011010101101011111",
27298 => "000111100011011000010010",
27299 => "001000110101001100110111",
27300 => "001000100011011000000000",
27301 => "000110001101101000100100",
27302 => "000011001110010110100011",
27303 => "000000100001111101000101",
27304 => "111111010101111101000110",
27305 => "111111110000010100001000",
27306 => "111111100001011111011111",
27307 => "111110110100010011000000",
27308 => "000000011000100111010011",
27309 => "000011111101001101010001",
27310 => "000111000111000110101111",
27311 => "001001001110010100010100",
27312 => "001010111101101000010010",
27313 => "001100100010010110100010",
27314 => "001100111111101001001100",
27315 => "001010110001110101000010",
27316 => "000101101100110111111000",
27317 => "111111111111000001011111",
27318 => "111100000110110100111001",
27319 => "111001110100101100011100",
27320 => "110111100101010011101000",
27321 => "110101101000001011111100",
27322 => "110100100100010111011000",
27323 => "110011010110110100001110",
27324 => "110000111111101100101000",
27325 => "101110010110111100101000",
27326 => "101100110111011011110010",
27327 => "101100000100000110110100",
27328 => "101011000110001001010000",
27329 => "101010111101110101110010",
27330 => "101100000011000111110100",
27331 => "101101110010011100110100",
27332 => "110000111011001110010100",
27333 => "110100101111000111100101",
27334 => "110110111000101001000000",
27335 => "110111101001110000010011",
27336 => "111000100011100000000111",
27337 => "111001100010100101100001",
27338 => "111010000110111010100010",
27339 => "111010101000010011101000",
27340 => "111011111100000111000010",
27341 => "111101011000111110100000",
27342 => "111110001001000110000110",
27343 => "111111101001111000101100",
27344 => "000010010101111011010001",
27345 => "000101001000100011101110",
27346 => "001001000000111111101110",
27347 => "001110010101000110101100",
27348 => "010011111011011110100000",
27349 => "011001100111011111000011",
27350 => "011101101110010101011001",
27351 => "011110101011010010101111",
27352 => "011110011001001010100000",
27353 => "011110010001010110110110",
27354 => "011101110011010001101010",
27355 => "011101001001011001001101",
27356 => "011100100011101010100011",
27357 => "011100000001000100011101",
27358 => "011011011101110100101101",
27359 => "011010110100011111010001",
27360 => "011010010010110101001100",
27361 => "011001101000100110101110",
27362 => "011000110111110110011001",
27363 => "011000100100110101000001",
27364 => "011000011111100000000101",
27365 => "011000101001000111001001",
27366 => "011000010100001110000101",
27367 => "010101110101001110001110",
27368 => "010011000110100000000000",
27369 => "010010101001111000000010",
27370 => "010010011101111001001010",
27371 => "010000100001100011110110",
27372 => "001100101110111011100100",
27373 => "000110101111010011011100",
27374 => "111111001011000101011111",
27375 => "110111001111100110010110",
27376 => "110000100110001110010000",
27377 => "101100101000101101010010",
27378 => "101001001010111010011100",
27379 => "100100100010010010111000",
27380 => "100001011101100100110100",
27381 => "100001000111011110000110",
27382 => "100001011011010111111000",
27383 => "100001000101011111011001",
27384 => "100001000011011001011101",
27385 => "100100010100100001011011",
27386 => "101011001110000001010110",
27387 => "110001101111101111111100",
27388 => "110110001011010100000110",
27389 => "111001001101111000101110",
27390 => "111010000100110010011010",
27391 => "111001100011011010110011",
27392 => "111010011001111011000000",
27393 => "111101000110111110011001",
27394 => "111111100011100011110001",
27395 => "111111001111110010011011",
27396 => "111011111100101010000010",
27397 => "110111110111110010101001",
27398 => "110100100111100000000000",
27399 => "110010100111001001100100",
27400 => "110001010101001100100010",
27401 => "101111100101000101010010",
27402 => "101111000111001100011010",
27403 => "110011000011010010110000",
27404 => "111001100000111110111010",
27405 => "111110100110110111111001",
27406 => "000010110001101101000100",
27407 => "001000001111110110010101",
27408 => "001110111011000110110110",
27409 => "010101000111101101111010",
27410 => "011001100101010101110101",
27411 => "011100011100000100100101",
27412 => "011101001011111000110101",
27413 => "011001000111001011011011",
27414 => "001111110000010101110110",
27415 => "000110001000110010111110",
27416 => "000001001001100110001100",
27417 => "111111111000000101010011",
27418 => "111110110011000101010001",
27419 => "111101101001011010000001",
27420 => "111110000011100110101101",
27421 => "111110111111010101000000",
27422 => "111110111101000011100011",
27423 => "111111010111110110000011",
27424 => "000000111110011011011011",
27425 => "000001111101010101101011",
27426 => "000001100111101000001101",
27427 => "000000110110011111010010",
27428 => "111111111011100011100011",
27429 => "111110000010010010101010",
27430 => "111010011111111001011101",
27431 => "110110110101101001000110",
27432 => "110101000100111110011100",
27433 => "110100011101101101100100",
27434 => "110011101110001110010110",
27435 => "110010111011011111100000",
27436 => "110001101011101010101110",
27437 => "110000001010010100000100",
27438 => "101111011011101011111110",
27439 => "101111001010111101001100",
27440 => "101111101110110011000110",
27441 => "110011001000000010100110",
27442 => "111000101100100010011111",
27443 => "111101100100101101001000",
27444 => "000001010000110000101110",
27445 => "000100011001001110100100",
27446 => "000101101100010111111011",
27447 => "000100000000100011010001",
27448 => "000000010100111110110101",
27449 => "111100001111110100011001",
27450 => "111000111010010100000011",
27451 => "110110101111010110100010",
27452 => "110101001100010011101111",
27453 => "110100101110000000011100",
27454 => "110111001111111110011101",
27455 => "111100101011100010100001",
27456 => "000010010110110110111100",
27457 => "000110110111101011010010",
27458 => "001010101101001111101100",
27459 => "001101110000100111100000",
27460 => "001110111110011111001100",
27461 => "001101101101100111101100",
27462 => "001010000101001100010111",
27463 => "000100111101111110001000",
27464 => "000000000110000011011011",
27465 => "111100101111101000010001",
27466 => "111010100100111001101101",
27467 => "111000101010110000101001",
27468 => "110110111101001110010010",
27469 => "110101110111010001010010",
27470 => "110101000011111100010000",
27471 => "110011111000011100001100",
27472 => "110010110010010010111100",
27473 => "110010010010000010111110",
27474 => "110001100111011001100110",
27475 => "110000110101110101100100",
27476 => "110001000011000110111100",
27477 => "110010001010111010101100",
27478 => "110011111000111101101010",
27479 => "110110000001101010100001",
27480 => "110111000100110100011100",
27481 => "110110011100001010101110",
27482 => "110101111111110001000101",
27483 => "110110110001000100011010",
27484 => "110111010101001001010101",
27485 => "110110011111111000000010",
27486 => "110101010000011011111010",
27487 => "110100111110101000110101",
27488 => "110101000111011101010001",
27489 => "110101000010000110100100",
27490 => "110101111011000010111001",
27491 => "111000010001110100000110",
27492 => "111011000000111010100111",
27493 => "111110000010100000111010",
27494 => "000001111000101010110100",
27495 => "000101111101100000111000",
27496 => "001001100100011000001010",
27497 => "001100100011111110000000",
27498 => "001110110111100011001000",
27499 => "010000111001001100000100",
27500 => "010010111100110100100110",
27501 => "010100010011110010111110",
27502 => "010100101011101100010010",
27503 => "010101001000011111111110",
27504 => "010110011001001000111100",
27505 => "010111111110000101101110",
27506 => "011001000100110011111011",
27507 => "011001111001001101000111",
27508 => "011011001110101000010101",
27509 => "011100001011010110011110",
27510 => "011011000110011000110011",
27511 => "011001010000000010000001",
27512 => "011000100010011001101100",
27513 => "010111101010100001110000",
27514 => "010101100110011100000110",
27515 => "010100011110111100010110",
27516 => "010101010000100000011010",
27517 => "010101011110111001101010",
27518 => "010011101000101111000000",
27519 => "010001000011101110011100",
27520 => "001110110100011101010110",
27521 => "001100011110111101110010",
27522 => "001001110001100101110100",
27523 => "000111011001110010000100",
27524 => "000110010000010001011101",
27525 => "000100101110101001011001",
27526 => "111111010101010011001111",
27527 => "110111001101111100010000",
27528 => "110001101101100111100110",
27529 => "101111111010100101010010",
27530 => "101111100101100010000010",
27531 => "110000111110011111101100",
27532 => "110100010100111111100100",
27533 => "110111100100100001110011",
27534 => "111001000111111111010010",
27535 => "111000100010101001101001",
27536 => "110101110101001110000111",
27537 => "110010001101011101101000",
27538 => "101111110011100010111010",
27539 => "101111101001010011111110",
27540 => "110000101101001111100010",
27541 => "110001110101100111111010",
27542 => "110010110011010000111000",
27543 => "110010110110011101111110",
27544 => "110001110001010000110110",
27545 => "110001111000100110100110",
27546 => "110101010010110010101101",
27547 => "111001101111000100101110",
27548 => "111011010100000111000000",
27549 => "111011011101001000011010",
27550 => "111110011011000011011111",
27551 => "000010001111011101001011",
27552 => "000010011010010001101011",
27553 => "000001000110010001000010",
27554 => "000001111010101111100011",
27555 => "000011001010111100111010",
27556 => "000011001010111100011111",
27557 => "000011011100101111001100",
27558 => "000100010110000010110101",
27559 => "000011110011010000100000",
27560 => "000000111100001100100101",
27561 => "111110000010101011111000",
27562 => "111110011011011010100100",
27563 => "000010101110110101011000",
27564 => "001000000100011001011001",
27565 => "001011110011010001111101",
27566 => "001110010101011010000000",
27567 => "010000001101000010110110",
27568 => "010000011110100010011100",
27569 => "001111111110110010001010",
27570 => "010000001111011010011010",
27571 => "010000001010011101010110",
27572 => "001110101001101011010110",
27573 => "001100010001001101000010",
27574 => "001001100001100110001010",
27575 => "000111011100110000010000",
27576 => "000110100000110101001000",
27577 => "000101001010011000001100",
27578 => "000011011000101000000011",
27579 => "000011001010001101000001",
27580 => "000100000011101001100110",
27581 => "000011111011001110000000",
27582 => "000010001101100010000110",
27583 => "111111100011110011010101",
27584 => "111100110000100000111011",
27585 => "111010011100010110101010",
27586 => "111001001110101011110001",
27587 => "111010100111001111110001",
27588 => "111111000001001101101000",
27589 => "000011101101100000010011",
27590 => "000110111100110001000011",
27591 => "001010001001001001101010",
27592 => "001100101010000010101110",
27593 => "001011010010111100000101",
27594 => "000101010101000100000111",
27595 => "111100100101001110110010",
27596 => "110011101100111101110010",
27597 => "101101011011101000110000",
27598 => "101001011011011010011110",
27599 => "100101001011101000101011",
27600 => "100010000000110111011110",
27601 => "100100000001110001010101",
27602 => "101011001011100111000110",
27603 => "110011011110101000001000",
27604 => "111010111110011000011011",
27605 => "000010010111110100000101",
27606 => "001001000011101010111010",
27607 => "001100111110000011011010",
27608 => "001101000011100110001000",
27609 => "001001101110011011110111",
27610 => "000100010101111010001110",
27611 => "111110001100101101101101",
27612 => "110111111000010101011111",
27613 => "110010010001111000011000",
27614 => "101110001010101101000010",
27615 => "101010110101111100000100",
27616 => "100111010111011000000101",
27617 => "100100010110111000100100",
27618 => "100011101010000100101101",
27619 => "100101110101001101010111",
27620 => "101001000000001011111110",
27621 => "101100001100000111001100",
27622 => "110000100101111111101100",
27623 => "110101111001101010111110",
27624 => "111010011110100011100111",
27625 => "111110010011100100010010",
27626 => "000001001001001001111001",
27627 => "000001010011000100100111",
27628 => "111110101001101100011110",
27629 => "111011001011001010100101",
27630 => "110111111000100011001110",
27631 => "110100011001111000010000",
27632 => "110001101101011110101010",
27633 => "110001101011100010001000",
27634 => "110011101101011000010010",
27635 => "110101110110000010000010",
27636 => "111000001101011100100101",
27637 => "111011101001101110011010",
27638 => "111111100011010111000110",
27639 => "000011010100110010100001",
27640 => "000111000100101111110010",
27641 => "001010001101000110011011",
27642 => "001100000010011011111110",
27643 => "001100110111011011110000",
27644 => "001100101100100000111010",
27645 => "001011100100110111110010",
27646 => "001010111111001100000000",
27647 => "001011001111011101101110",
27648 => "001010100000001111101010",
27649 => "001000111011101100011110",
27650 => "001000011100000100010010",
27651 => "001000101110000101011000",
27652 => "001000111110110000100010",
27653 => "001010001110111110010011",
27654 => "001100010000010100010100",
27655 => "001100110110010001101100",
27656 => "001011110110010011010110",
27657 => "001011100110011010111101",
27658 => "001101000010001101110110",
27659 => "001110010110001100011000",
27660 => "001101011100101000001000",
27661 => "001010110000101010001001",
27662 => "001001001001111111100100",
27663 => "001001010111110000010001",
27664 => "001000010101011101101000",
27665 => "000101001000000001000101",
27666 => "000010011100011110011000",
27667 => "000000111001010101010111",
27668 => "111110110111011101011001",
27669 => "111100010100110000001100",
27670 => "111010101111000110000101",
27671 => "111011000000111111011110",
27672 => "111010111010101010011010",
27673 => "110111000001100100101000",
27674 => "110001101001101001000010",
27675 => "110000011101001101000110",
27676 => "110011110100010010010010",
27677 => "111000100110010011010101",
27678 => "111101101101110111111101",
27679 => "000010101001001111110000",
27680 => "000110001000100000001111",
27681 => "000111101111010010111010",
27682 => "000111011010100011000011",
27683 => "000101111100101010100111",
27684 => "000110000111001110000101",
27685 => "001000111001001100010000",
27686 => "001011001100101101000100",
27687 => "001011100010010111111100",
27688 => "001011011001010110101110",
27689 => "001001101011001001100111",
27690 => "000101010001010010000001",
27691 => "000001111001101011001011",
27692 => "000010000011010010100011",
27693 => "000010111000000110110011",
27694 => "000010000000010011110001",
27695 => "000000111000010110101001",
27696 => "000001010101101011000000",
27697 => "000010010011110100100011",
27698 => "000001110011100110011100",
27699 => "000000100001010011101000",
27700 => "111111101000100111011001",
27701 => "111110010111011110101101",
27702 => "111100111000001011000110",
27703 => "111100000101001000100100",
27704 => "111010110011111000010000",
27705 => "111000000111011010000110",
27706 => "110101000001010010100010",
27707 => "110010011100111011001010",
27708 => "110001011010000011110000",
27709 => "110011101011001100001010",
27710 => "111001010100101111110100",
27711 => "111111110010100010011100",
27712 => "000100110100110010000000",
27713 => "000111110011101011010111",
27714 => "001000001101010100001011",
27715 => "000101111110100110100101",
27716 => "000010111000010100100010",
27717 => "000000101110101110001000",
27718 => "111111000110111011110110",
27719 => "111100001001111000001001",
27720 => "110111010101110011101101",
27721 => "110010110010101011000000",
27722 => "110000110011100000110100",
27723 => "110000111011010001100000",
27724 => "110001101100000000010000",
27725 => "110011111111101010110000",
27726 => "111001011111011011110010",
27727 => "000000001011110111001010",
27728 => "000011111001011010101101",
27729 => "000011111110100111100010",
27730 => "000011000010011111010100",
27731 => "000010000111110000011110",
27732 => "000000110110001010010110",
27733 => "000000010110101011000111",
27734 => "000010010110001110000000",
27735 => "000110100001110001011110",
27736 => "001010111101101101010111",
27737 => "001110001111101010110010",
27738 => "010000000000100000100000",
27739 => "010000100000000010111100",
27740 => "010000100000110111010000",
27741 => "001111110100001010101100",
27742 => "001100110110011111110000",
27743 => "001000010000001110100000",
27744 => "000100101011111010111011",
27745 => "000010010001000011101000",
27746 => "111111011001100001010010",
27747 => "111101000001110110100101",
27748 => "111101010001110110111100",
27749 => "111111110111011101111111",
27750 => "000011000011001001110110",
27751 => "000110001101010011110010",
27752 => "001001011011011000111010",
27753 => "001011111010101000101011",
27754 => "001100010101111101110000",
27755 => "001010001101000011011010",
27756 => "000110010101100001111111",
27757 => "000010010001110000000100",
27758 => "111110110110111110101110",
27759 => "111011001011111001110010",
27760 => "110101111100110110110100",
27761 => "110000000010011000111100",
27762 => "101011001001100110011010",
27763 => "100110110110111111011101",
27764 => "100011011001100011001011",
27765 => "100010101111001110101011",
27766 => "100011110010111011000010",
27767 => "100100110100010011100100",
27768 => "100111100111100111100001",
27769 => "101100001011010101000110",
27770 => "110000001100110101010010",
27771 => "110100011111110110111010",
27772 => "111001000011101011010000",
27773 => "111011001011101011110110",
27774 => "111011000111100011110101",
27775 => "111010100111001110010100",
27776 => "111001011101001111111100",
27777 => "110111101000011101100011",
27778 => "110101110100011100010000",
27779 => "110100101101100010010110",
27780 => "110101001011111111000011",
27781 => "110111010011101001000101",
27782 => "111010100011011110111110",
27783 => "111110101011001000001111",
27784 => "000011010000111100011111",
27785 => "000111101110010001110010",
27786 => "001011100101110100001011",
27787 => "001111001000001000011000",
27788 => "010010100010110110001100",
27789 => "010100110011100011101010",
27790 => "010101101010101000101100",
27791 => "010110001110010000100110",
27792 => "010110010110010010011100",
27793 => "010101101010111001110100",
27794 => "010100101011101010000100",
27795 => "010011011010110110111000",
27796 => "010010100100111101101010",
27797 => "010011000011001111101100",
27798 => "010011101100000011010010",
27799 => "010011101001101101111010",
27800 => "010011111111010111101100",
27801 => "010100111101011110110010",
27802 => "010101010010010010001000",
27803 => "010011111011000100011010",
27804 => "010001100010010111101110",
27805 => "001111101100101101010110",
27806 => "001101111110101010111010",
27807 => "001010110000000100101011",
27808 => "000110110000110100010110",
27809 => "000011010010110000010001",
27810 => "111110101001010000001010",
27811 => "110111011101101101101001",
27812 => "110000100110001110111110",
27813 => "101101001111011100001000",
27814 => "101100101110000100010110",
27815 => "101100110110111010011110",
27816 => "101100110111110010000100",
27817 => "101101001000010011111010",
27818 => "101101110001110010010110",
27819 => "101101001010000000100110",
27820 => "101010000101100111010110",
27821 => "100111101001001011010111",
27822 => "101001010110110010100100",
27823 => "101101111110000100111110",
27824 => "110010011000101101011000",
27825 => "110110000001110000011111",
27826 => "111001101000011110001000",
27827 => "111011111101000111001010",
27828 => "111010101110110010011000",
27829 => "110111101101100010101111",
27830 => "110111101100100100101111",
27831 => "111011001000000101101110",
27832 => "111110000010101001011001",
27833 => "111111000101111110100100",
27834 => "000000011111111101010010",
27835 => "000010111001000101010100",
27836 => "000100001111101011011011",
27837 => "000100011001111110011101",
27838 => "000110000111111011000101",
27839 => "001010001110000111001101",
27840 => "001101111101011101110100",
27841 => "001110111010111110011000",
27842 => "001101110101001010110010",
27843 => "001101000000110011010110",
27844 => "001100101010011110100000",
27845 => "001011010110111111100111",
27846 => "001001110110101100010010",
27847 => "001001110000111011100000",
27848 => "001010111101001010101101",
27849 => "001101000111011100111000",
27850 => "001111011111001101100000",
27851 => "010000000000011100010100",
27852 => "001101111011000010111000",
27853 => "001010001110111001010101",
27854 => "000110001000101101011010",
27855 => "000011110000101101001110",
27856 => "000101011000100000100010",
27857 => "001001110101010111001100",
27858 => "001100101110000011111000",
27859 => "001100001010110001010000",
27860 => "001010011101101111110010",
27861 => "001000100001001100101111",
27862 => "000100111101110110001111",
27863 => "000000100110111011001010",
27864 => "111101010010011010110111",
27865 => "111001111101001100110011",
27866 => "110011011010011010111110",
27867 => "101001100111101111010000",
27868 => "100010011111100000100111",
27869 => "100001011011101000010111",
27870 => "100001100110110111001111",
27871 => "100001001000010011000011",
27872 => "100100111110001001100001",
27873 => "101100111111011110110100",
27874 => "110100010110100100101000",
27875 => "111010101100000000100011",
27876 => "000000101011111110001110",
27877 => "000011110110010110110101",
27878 => "000011000110010111011001",
27879 => "000000111001100101011000",
27880 => "111111101100100000000001",
27881 => "111111010011001000011101",
27882 => "111110010101100011100101",
27883 => "111100100011001100011110",
27884 => "111010100111100010111001",
27885 => "111001010101001111100000",
27886 => "111000110011110000001110",
27887 => "111000010100001100100000",
27888 => "111000000001110011010010",
27889 => "111000110001001000001100",
27890 => "111010010101011001010000",
27891 => "111100101001000001111000",
27892 => "111111101110011000100010",
27893 => "000010111100000001011000",
27894 => "000110110000110010110111",
27895 => "001011110101010001111111",
27896 => "010000110000111000010000",
27897 => "010100110101010101110100",
27898 => "011000101100110111110101",
27899 => "011011001110101011110000",
27900 => "011010101001001000001110",
27901 => "010111010000010001011000",
27902 => "010001111000111101100000",
27903 => "001011000001011111110100",
27904 => "000100100000001101000110",
27905 => "000000010110011001001101",
27906 => "111110000000000110011100",
27907 => "111011100111011101111000",
27908 => "111000110101001000101001",
27909 => "110110001110110101110001",
27910 => "110011101011000001001000",
27911 => "110000101100010001001110",
27912 => "101101111101000100101110",
27913 => "101100110100010000111110",
27914 => "101101100010011011010110",
27915 => "101111100011101111110010",
27916 => "110010110110110100110100",
27917 => "110111001001111000011100",
27918 => "111011001010110110011011",
27919 => "111101110100101011000111",
27920 => "111110111011110101111100",
27921 => "111110110010100000001010",
27922 => "111101101111101011001100",
27923 => "111011101110000100101000",
27924 => "110111111100010010110011",
27925 => "110010010101010111000010",
27926 => "101100111001001111011110",
27927 => "101001101010001100101000",
27928 => "101000001100000100001000",
27929 => "100111101010111001010111",
27930 => "101001000010011001011010",
27931 => "101100110110111001000100",
27932 => "110010011001100101110110",
27933 => "111001010001001000111110",
27934 => "000001001000011001001111",
27935 => "001000100001111111010100",
27936 => "001101111010010101111000",
27937 => "010001001001000100010110",
27938 => "010010110011101100111110",
27939 => "010011010001010010111010",
27940 => "010011001010011101011110",
27941 => "010010100011110110010000",
27942 => "010000101001000001001110",
27943 => "001110010101100000110010",
27944 => "001101011000010001000110",
27945 => "001101000011101011111000",
27946 => "001101000001110110100000",
27947 => "001110111110111000101110",
27948 => "010001111101011000101110",
27949 => "010010110111000010001100",
27950 => "010001111110100110011100",
27951 => "010001100110001011110100",
27952 => "010001001111111001100010",
27953 => "001111000101111101011000",
27954 => "001011011000011001100100",
27955 => "000111110100001110001111",
27956 => "000101011010010101000010",
27957 => "000011011111011000001100",
27958 => "000000011111101100110100",
27959 => "111101001010000011001111",
27960 => "111100001011000001001010",
27961 => "111101001101010011010000",
27962 => "111101110100011110000001",
27963 => "111110000101011011001100",
27964 => "111110001100011111011011",
27965 => "111100001100111000110010",
27966 => "110111101110111111000100",
27967 => "110010111010101000001000",
27968 => "101111110001010010001100",
27969 => "101110111111110100110110",
27970 => "101111101100110010001000",
27971 => "110000101101001101011110",
27972 => "110001110100011011101100",
27973 => "110010011111101000110100",
27974 => "110001111000001001101100",
27975 => "110000100101111110110100",
27976 => "110000001001110011000110",
27977 => "110001100101110001011000",
27978 => "110101011110001001000110",
27979 => "111011010011110110010000",
27980 => "000001010011001011110100",
27981 => "000101110101101110101001",
27982 => "000111111100001010111010",
27983 => "000110111001111111011010",
27984 => "000100001101010010010000",
27985 => "000011000000100111000011",
27986 => "000011100101000000001010",
27987 => "000010101101001010000110",
27988 => "111110101100111110110001",
27989 => "111010000010011111010110",
27990 => "110111110001000110010001",
27991 => "110111010100110100011000",
27992 => "110111011101000000100000",
27993 => "111001111100111110010111",
27994 => "111111010110010010101001",
27995 => "000101000111111101000010",
27996 => "001010100000101000001001",
27997 => "001111000010111000010000",
27998 => "010000010101100011010110",
27999 => "001110111010001101111000",
28000 => "001101101100111010000010",
28001 => "001101001000000111101100",
28002 => "001101011100001101000110",
28003 => "010000011101000110100100",
28004 => "010101000111101110101100",
28005 => "011000000001010011101100",
28006 => "011000010101111011110011",
28007 => "010110111000111000101100",
28008 => "010011110001010010000110",
28009 => "010000110011110001110000",
28010 => "001111101110010110100110",
28011 => "001110001110101011110100",
28012 => "001010100011110100000010",
28013 => "000101111110011011111111",
28014 => "000000100011000010011001",
28015 => "111010111101000000001101",
28016 => "111000000011011110111001",
28017 => "111000000100000011001110",
28018 => "111001110100101110100001",
28019 => "111101110101011010010101",
28020 => "000010110011011101100110",
28021 => "000110001111011010010000",
28022 => "000111111101010101100011",
28023 => "001000001010010000010000",
28024 => "000110010011101100001010",
28025 => "000010110110101001101010",
28026 => "111110110011010110001110",
28027 => "111010111101011011100100",
28028 => "111000001100010110001111",
28029 => "110110011100010010010100",
28030 => "110100100100101100010111",
28031 => "110010001101100010001000",
28032 => "101111010101001101111100",
28033 => "101011011101101010011100",
28034 => "101000011011100101110110",
28035 => "101000111011101100011000",
28036 => "101011011110110011000100",
28037 => "101101111001110011111100",
28038 => "110001101011110000101000",
28039 => "110111100000100001000111",
28040 => "111101111101001110001010",
28041 => "000100100110001000000000",
28042 => "001010100111000111100100",
28043 => "001110100000100011101000",
28044 => "010000011001110001110000",
28045 => "010000110011111110010000",
28046 => "001111000010010010011110",
28047 => "001010010101100110000011",
28048 => "000010111110101111111001",
28049 => "111001110100110100100001",
28050 => "110000110101101101000100",
28051 => "101011110110001011000100",
28052 => "101100101111000001001010",
28053 => "110000000011000011101010",
28054 => "110010001000000001100100",
28055 => "110011110111110100011010",
28056 => "110110110010010010010010",
28057 => "111001010011111100100110",
28058 => "111001111111011111100111",
28059 => "111010011100000100010110",
28060 => "111100000110001001000101",
28061 => "111101100111110010000010",
28062 => "111110010001011001010010",
28063 => "111110101000000100111101",
28064 => "111110001010110101110101",
28065 => "111101001110011111011100",
28066 => "111100111100000000100110",
28067 => "111100110011101100111100",
28068 => "111101001000100000010100",
28069 => "111110111110001000101000",
28070 => "000000111110100101001110",
28071 => "000001100011010110100100",
28072 => "000000100011101111100000",
28073 => "111110000101110001011110",
28074 => "111011010000100011100110",
28075 => "111001100100111010000110",
28076 => "111000111110111001101000",
28077 => "111000110101111110001001",
28078 => "111001011001001011101111",
28079 => "111011010100111011110100",
28080 => "111110110101011111001000",
28081 => "000011010110011110011111",
28082 => "000111111001111001000000",
28083 => "001011110001000101011010",
28084 => "001111001100110001111000",
28085 => "010010010110000011111010",
28086 => "010100001110110010101100",
28087 => "010100100001110000010100",
28088 => "010011001010111000100100",
28089 => "001111100110101111011110",
28090 => "001011001111111000010100",
28091 => "000111101111000011001010",
28092 => "000100011010110111111110",
28093 => "000001100110011100000110",
28094 => "000000001000100000010101",
28095 => "111111000001011000101110",
28096 => "111110000001010011001100",
28097 => "111101110100000000001101",
28098 => "111110011101111111110110",
28099 => "000000001110111100111000",
28100 => "000010011011111010101100",
28101 => "000011111110010111001110",
28102 => "000101001111001010110001",
28103 => "000101110111011001010100",
28104 => "000100011001000101110110",
28105 => "000001001110011101101111",
28106 => "111101111101011100100110",
28107 => "111011001011000111011110",
28108 => "111001000100101101011110",
28109 => "111000010001111100001111",
28110 => "111000000110101111011100",
28111 => "110110011011001110001001",
28112 => "110011011100001011100100",
28113 => "110001101000010100101010",
28114 => "110010000010010111011000",
28115 => "110100011100110110111101",
28116 => "110111110101001001001111",
28117 => "111010010010010101110111",
28118 => "111011100111000101111011",
28119 => "111100000010100001100000",
28120 => "111010100010101110100100",
28121 => "110111111001010101111110",
28122 => "110110001101011010110000",
28123 => "110110010100111000001000",
28124 => "111000101001000111111111",
28125 => "111100101111101001001111",
28126 => "000001011001011000110000",
28127 => "000110000011110110100000",
28128 => "001001110110110000000101",
28129 => "001011101010000010010010",
28130 => "001011111000001100110000",
28131 => "001011011001100011111100",
28132 => "001010001000111110001110",
28133 => "000111101100011101111010",
28134 => "000011110101000011010000",
28135 => "111101111110001110111010",
28136 => "110110010000101100001011",
28137 => "101111011110111000111110",
28138 => "101100010111101001101010",
28139 => "101100010100001101100000",
28140 => "101110001001111000010100",
28141 => "110001110000111111010000",
28142 => "110110100110110101011110",
28143 => "111100000100110101010110",
28144 => "000000010001010110000011",
28145 => "000000110000000110111011",
28146 => "111111010100110111101100",
28147 => "111111011011100000111010",
28148 => "000000100010101001010011",
28149 => "000001011001111110011101",
28150 => "000011001000000001011011",
28151 => "000101110101000100001100",
28152 => "000111011110111100010100",
28153 => "000110111100001100010110",
28154 => "000100111010000110011110",
28155 => "000010010011000111000010",
28156 => "000000100100101100001100",
28157 => "000001001010100011100111",
28158 => "000001111011110100000010",
28159 => "111111010101111000001000",
28160 => "111010001100001010101110",
28161 => "110101111000111011110001",
28162 => "110100000101010101011011",
28163 => "110100100101111111010000",
28164 => "110110110100111011001010",
28165 => "111010110001111110010101",
28166 => "000000000010001000000111",
28167 => "000100101001001101010100",
28168 => "000111100000001011000001",
28169 => "001001001100111001110110",
28170 => "001010001110100100100011",
28171 => "001011001110000010100111",
28172 => "001100111010000010110010",
28173 => "001110110000100111110100",
28174 => "001111111111101010011000",
28175 => "010000111101100110110110",
28176 => "010010000000001110011110",
28177 => "010010010100101101110110",
28178 => "010001100000011100101010",
28179 => "010000011100010000001010",
28180 => "001111011001001010101010",
28181 => "001101110110111001001110",
28182 => "001011111100011010011110",
28183 => "001001010111000110000011",
28184 => "000110000111011101010000",
28185 => "000100010011101011010100",
28186 => "000100111100000001000011",
28187 => "000101111010101101111011",
28188 => "000110010001001100111001",
28189 => "000111101001110010000101",
28190 => "001010001001010010100000",
28191 => "001011011101100000001110",
28192 => "001011000011100000000010",
28193 => "001010000001101110011100",
28194 => "000111100111111110111011",
28195 => "000010100100101101000100",
28196 => "111011110111000010101101",
28197 => "110101100111110100011100",
28198 => "110001010010010100011110",
28199 => "101110101000101101010110",
28200 => "101100101001000100000000",
28201 => "101011100001001001011010",
28202 => "101011110000101011101000",
28203 => "101100110011010011010010",
28204 => "101110100100111100001010",
28205 => "110001011010001101001110",
28206 => "110100010111000111101100",
28207 => "110110001100000100111110",
28208 => "110111001000100000101100",
28209 => "111000010000011011001101",
28210 => "111001011011101101011011",
28211 => "111001111111111010100011",
28212 => "111010010101110100100011",
28213 => "111010010111010010110001",
28214 => "111001010100111011100011",
28215 => "110111111110111100000000",
28216 => "110111100110110100111111",
28217 => "111000010111111111001101",
28218 => "111001100110101100100110",
28219 => "111010011101010001000001",
28220 => "111011100101010111011111",
28221 => "111110010101100001100111",
28222 => "000010001000000000100000",
28223 => "000101101000011001111000",
28224 => "001000100101001000100011",
28225 => "001011001000100011011000",
28226 => "001101111101010011001010",
28227 => "010001110000100011000100",
28228 => "010101101110000111101110",
28229 => "011000000000011000011111",
28230 => "011000100110001010110011",
28231 => "011001011110111001101011",
28232 => "011010100011000000000100",
28233 => "011010000001011110111000",
28234 => "011000110110010011110101",
28235 => "011000000111010111111011",
28236 => "010110110000101111100110",
28237 => "010100110010000100010010",
28238 => "010010011010001110101110",
28239 => "001111010100101100111000",
28240 => "001100100011010100010010",
28241 => "001001111000011001111000",
28242 => "000101101010000000000011",
28243 => "000000100110011101101001",
28244 => "111100110111100000000110",
28245 => "111011101110100110001110",
28246 => "111100111111110000001100",
28247 => "111111001011101101001111",
28248 => "000001001101011111110110",
28249 => "000010100100010011110100",
28250 => "000010111001001001011010",
28251 => "000010001000100000110100",
28252 => "000000000000011000000110",
28253 => "111101010111010110111011",
28254 => "111010110010000010110011",
28255 => "110110110110111010010010",
28256 => "110011000000100011100000",
28257 => "110000011000100000101010",
28258 => "101011000011010110010010",
28259 => "100100001011000000101001",
28260 => "100001011010101110110011",
28261 => "100001010110101100111000",
28262 => "100010010111000000110111",
28263 => "100110110010011011010000",
28264 => "101100001001111010110010",
28265 => "101111100011110110101000",
28266 => "110010000010010100010100",
28267 => "110010111101100011101010",
28268 => "110010101110011101010010",
28269 => "110100000011111111000000",
28270 => "110110111011011110101000",
28271 => "111010100110101101110001",
28272 => "111111101110011000110100",
28273 => "000101011011100010011100",
28274 => "001001111011110000110110",
28275 => "001100110001110000110000",
28276 => "001110101011010011111100",
28277 => "001111011011011110110010",
28278 => "001110001010000000111110",
28279 => "001100000100111011010100",
28280 => "001010000001110110100010",
28281 => "000101110010111010111000",
28282 => "111110100111000111011100",
28283 => "110110101011011110110100",
28284 => "110000001000001010110110",
28285 => "101100110100001100010010",
28286 => "101101100010111111011010",
28287 => "110000111000100110000010",
28288 => "110101000100010101100000",
28289 => "111001001010110001011111",
28290 => "111100111011110000010011",
28291 => "000000100101101011010010",
28292 => "000011100001001100111011",
28293 => "000100101001000001100101",
28294 => "000101000001011111010110",
28295 => "000110111101001010010101",
28296 => "001001100110011010110100",
28297 => "001010000010011011100111",
28298 => "001000100001101000010010",
28299 => "000110101110110110101000",
28300 => "000011100100001101110100",
28301 => "111110101011101000010001",
28302 => "111010100101011111001100",
28303 => "111000011011000000010110",
28304 => "110111000000110110010011",
28305 => "110101000110100110000111",
28306 => "110010001001100011001100",
28307 => "101110101101000100000000",
28308 => "101011100101001001101000",
28309 => "101001010111010110001110",
28310 => "101001100110001001100010",
28311 => "101100111101011111001100",
28312 => "110000111101110101110100",
28313 => "110011010111000111010000",
28314 => "110101001111111100011000",
28315 => "110111110110000100100100",
28316 => "111010001010001111000001",
28317 => "111011101011001000000100",
28318 => "111101010000100010110100",
28319 => "111111100010001011111110",
28320 => "000010101101010101100110",
28321 => "000110000111110010100001",
28322 => "001000100000000001010000",
28323 => "001010001000110000111111",
28324 => "001011100101001111001001",
28325 => "001011111001101110010101",
28326 => "001011010011011111001100",
28327 => "001010111001000111000001",
28328 => "001010011000100001001000",
28329 => "001001111011110110100110",
28330 => "001001111101000011001100",
28331 => "001001011000000011100000",
28332 => "001000011010000101011101",
28333 => "001000100110110001100011",
28334 => "001001101110110000011100",
28335 => "001011010111010111001000",
28336 => "001110001001110010001100",
28337 => "010001010110101000101100",
28338 => "010011110110011000111000",
28339 => "010101111111010110011010",
28340 => "010111000110010110001000",
28341 => "010101010110001011011110",
28342 => "010001101101100001110000",
28343 => "001111000000011010101110",
28344 => "001101001110001001010000",
28345 => "001011000001111010110010",
28346 => "001001000010000001011100",
28347 => "000111000101000100110000",
28348 => "000011101101111011101111",
28349 => "111111110101001000000110",
28350 => "111101000001011110010100",
28351 => "111010101011110101100100",
28352 => "111000001001001100100010",
28353 => "110101110011101111101001",
28354 => "110100000111110010010001",
28355 => "110011000111101101000100",
28356 => "110001111100111010000000",
28357 => "110000011111110000100010",
28358 => "110000000100001111101110",
28359 => "110000001111100001111100",
28360 => "101111101000001000110010",
28361 => "101110101100100000100000",
28362 => "101101011101111101011010",
28363 => "101011000101100111010010",
28364 => "101000110101011101010000",
28365 => "101000110100100111001110",
28366 => "101011001110000011101000",
28367 => "101110100101100001110110",
28368 => "110001110110001111011000",
28369 => "110101011111010010101010",
28370 => "111001101110101001100011",
28371 => "111101100010100100011101",
28372 => "000000110010010010100100",
28373 => "000100000001011010100001",
28374 => "000111000011100011101000",
28375 => "001001011111010000011000",
28376 => "001010110111110010110000",
28377 => "001011011110110110000011",
28378 => "001100011111001110011000",
28379 => "001101001110110000010110",
28380 => "001100000001001110100110",
28381 => "001010000111001001001110",
28382 => "001010001010111110110011",
28383 => "001011111010010100101100",
28384 => "001101000110010110011000",
28385 => "001101011100000000010000",
28386 => "001101111011001011111110",
28387 => "001110001001000111000100",
28388 => "001101101100001101000010",
28389 => "001101010100111100000000",
28390 => "001101001100000111110100",
28391 => "001101100001000110001000",
28392 => "001111001010101110000100",
28393 => "010001111001001100100110",
28394 => "010100111111110011110000",
28395 => "010111011010011000101000",
28396 => "010111000011101100100010",
28397 => "010011101111110001001000",
28398 => "001111101001101111011100",
28399 => "001011111100001000000111",
28400 => "001000100001001101010110",
28401 => "000101010100011100000001",
28402 => "000010000001011110111010",
28403 => "111101110011111011011100",
28404 => "110111100000101110011101",
28405 => "101111000011011010100010",
28406 => "100111001101010001010010",
28407 => "100011100110100101001111",
28408 => "100100011000000110110111",
28409 => "100110110111101110001000",
28410 => "101010111000101000000100",
28411 => "110001010101011011100010",
28412 => "110111011011100011000010",
28413 => "111010111111001011101110",
28414 => "111101111010110011111000",
28415 => "000000111101110110110000",
28416 => "000011100000000011010000",
28417 => "000110011000001010011001",
28418 => "001000111000110000010110",
28419 => "001001001101110000010011",
28420 => "000111110000001000010101",
28421 => "000101010011011110001110",
28422 => "000010010110110011101101",
28423 => "000000000100111101110001",
28424 => "111110101110011111111010",
28425 => "111101101010001100000011",
28426 => "111100111011001101111111",
28427 => "111100011110011011111110",
28428 => "111011011101001001100100",
28429 => "111001100010100100011100",
28430 => "110111000110000110110110",
28431 => "110100010110100010111010",
28432 => "110010111100011111010010",
28433 => "110101001011110000100100",
28434 => "111001101111010010001001",
28435 => "111101101100110110011111",
28436 => "000000111100101101000011",
28437 => "000011001101011111101000",
28438 => "000011010101000110010110",
28439 => "000010100100001011110010",
28440 => "000010110111001011101001",
28441 => "000101001000010011101010",
28442 => "001001001111100101110000",
28443 => "001100111000100101000110",
28444 => "001110101101101110001010",
28445 => "010000001100100011111010",
28446 => "010000110111000010011110",
28447 => "001110101101010101011100",
28448 => "001010111011011010010110",
28449 => "000111101111100110010000",
28450 => "000100101000010111010010",
28451 => "000000100100001000100010",
28452 => "111100010010100011101011",
28453 => "110111110011110100100111",
28454 => "110010010000001100101010",
28455 => "101101011100111111010110",
28456 => "101011100011110001010010",
28457 => "101011010101110111001110",
28458 => "101011111011011010111110",
28459 => "101101111011101111110010",
28460 => "110000000111100000101010",
28461 => "110001010111001010101100",
28462 => "110010100110001010011110",
28463 => "110100011101001001001011",
28464 => "110110110011110011101011",
28465 => "111001011111111000000110",
28466 => "111100010101101100000101",
28467 => "111111000001010011010011",
28468 => "000000110100000111010000",
28469 => "000001111110100001101001",
28470 => "000011011001001101100100",
28471 => "000011011110000110000010",
28472 => "000000110010010111011010",
28473 => "111110010110111101000101",
28474 => "111110111011110101001011",
28475 => "000000001000000111100101",
28476 => "111110110100111110010111",
28477 => "111011111111010111111110",
28478 => "111010000110100111100100",
28479 => "111001010100101110000100",
28480 => "111000011001001000111010",
28481 => "110111001100011111000010",
28482 => "110110110110110011000010",
28483 => "111000110000001100001010",
28484 => "111101000110111111101001",
28485 => "000001111010010001000010",
28486 => "000101010111100010101001",
28487 => "001000011000100001010110",
28488 => "001011101011101011101000",
28489 => "001101111010110100100000",
28490 => "001110110111001110000000",
28491 => "001111111010011111001110",
28492 => "010000110110100100111100",
28493 => "001111111101000101001000",
28494 => "001100100011110001100000",
28495 => "000111011001011010100000",
28496 => "000001011001100010010100",
28497 => "111011100101110000111011",
28498 => "110111100011010010000100",
28499 => "110101110110001001100011",
28500 => "110101010101011101011001",
28501 => "110101111001101110011110",
28502 => "110111111111101110110000",
28503 => "111010000010011100100101",
28504 => "111011000011101000001101",
28505 => "111011111101010010110110",
28506 => "111100110110010011101011",
28507 => "111110000011000010000111",
28508 => "000000011001000110001000",
28509 => "000010111010100001110100",
28510 => "000100100111011111011011",
28511 => "000101110000110010011100",
28512 => "000110001101100000100011",
28513 => "000101111000010111010101",
28514 => "000101001101100111011001",
28515 => "000100101111101101001101",
28516 => "000100101110011111111011",
28517 => "000100000111110010100000",
28518 => "000010011110010001101000",
28519 => "000001011000010000001011",
28520 => "000001011101100101011000",
28521 => "000001110010011001111100",
28522 => "000010001100110010001000",
28523 => "000011010100101001111001",
28524 => "000101011101001100000000",
28525 => "000111010000001101001011",
28526 => "000110011111010100000111",
28527 => "000011000101110111001110",
28528 => "111110110010110100111001",
28529 => "111011010111100010111000",
28530 => "111001111010100101001010",
28531 => "111001100100011001010100",
28532 => "111001011011000110010010",
28533 => "111010100011011001000110",
28534 => "111101000110000000111101",
28535 => "000000000111011000110110",
28536 => "000011111111000011010111",
28537 => "001000100110111001010010",
28538 => "001100101100101011011110",
28539 => "001111110011011101101100",
28540 => "010010010100100001000010",
28541 => "010100010011000111001110",
28542 => "010100101011010101111010",
28543 => "010001110101101010101000",
28544 => "001011101001101000111001",
28545 => "000100001001111011010011",
28546 => "111101111100010001101000",
28547 => "111010000010011110101100",
28548 => "110111110000001100000010",
28549 => "110110001100101111101000",
28550 => "110100010010010000111111",
28551 => "110000101101111101101010",
28552 => "101100001110000100011100",
28553 => "101001110001110111001100",
28554 => "101011010111010011101110",
28555 => "101111101100100001011110",
28556 => "110100101001111011011000",
28557 => "111010100000001010011101",
28558 => "000001100011010000110111",
28559 => "000111011110010011001011",
28560 => "001010101011010100011000",
28561 => "001100011011100101000100",
28562 => "001110000100101110110100",
28563 => "001111010111001111010110",
28564 => "001111101011111000111010",
28565 => "001111101001001011000000",
28566 => "010000000000101110011000",
28567 => "001111011101010100001110",
28568 => "001100011010101111011010",
28569 => "000111111010000101011011",
28570 => "000100000100110111000010",
28571 => "000001110011000101110000",
28572 => "000000010001110011011101",
28573 => "111110010110101010001001",
28574 => "111011100001101101010100",
28575 => "110111111000010001111011",
28576 => "110100101001010100100101",
28577 => "110010101010101101000010",
28578 => "110000110110011110010110",
28579 => "110000010011000010111000",
28580 => "110100001000100101110000",
28581 => "111011001000011010011001",
28582 => "000001011011100100101010",
28583 => "000101001000001001101111",
28584 => "000101000101011010111101",
28585 => "000001110110001100011101",
28586 => "111110011000001111010010",
28587 => "111100011111010100100111",
28588 => "111011111010000011100101",
28589 => "111011110010011000111110",
28590 => "111011011101100101011000",
28591 => "111011000101011001110101",
28592 => "111011001110110111100100",
28593 => "111100000100111000010001",
28594 => "111100111101101111010000",
28595 => "111101100110111111010010",
28596 => "111111010100010011110101",
28597 => "000001011101101101011010",
28598 => "000000101101100000010011",
28599 => "111101000011110100011111",
28600 => "111001001100001110011000",
28601 => "110101001000101000111001",
28602 => "110000001111110111111010",
28603 => "101011100110011110100000",
28604 => "101000111000010101100010",
28605 => "101001110111111101111010",
28606 => "101110001110111110100110",
28607 => "110011000010111110101010",
28608 => "110111000001011011010110",
28609 => "111011100001100101010101",
28610 => "000001011100010010101010",
28611 => "000111110101010000010001",
28612 => "001101001110100111000100",
28613 => "010000111100001010001000",
28614 => "010010110101011000011000",
28615 => "010010101110110011000010",
28616 => "010000001101100010011010",
28617 => "001011010000011101010000",
28618 => "000101100000010001101101",
28619 => "000000101111111010000011",
28620 => "111101000110000111001010",
28621 => "111010111011101001111100",
28622 => "111010110100110111011001",
28623 => "111011010111010101110110",
28624 => "111011100101100011110010",
28625 => "111100001110010100100100",
28626 => "111100111000011110110110",
28627 => "111101000100011000111000",
28628 => "111110010010000101000111",
28629 => "000001001010111100011100",
28630 => "000100000011110111000000",
28631 => "000110010000001001011011",
28632 => "001000011111001001110110",
28633 => "001001111110100001100111",
28634 => "001001110001100111101111",
28635 => "001001000010111101110001",
28636 => "001000010001110011110000",
28637 => "000110110001011101010110",
28638 => "000101001011000101100100",
28639 => "000011101010111010110010",
28640 => "000001000001001110111100",
28641 => "111101010011000000001010",
28642 => "111001101011010001001010",
28643 => "110110101110111111101011",
28644 => "110100101011110111100000",
28645 => "110011011010110011011110",
28646 => "110010011100000110011100",
28647 => "110001001110101001010110",
28648 => "101111111111101011001000",
28649 => "101111110011110011011010",
28650 => "110000101001111001010110",
28651 => "110001100110000000011100",
28652 => "110011010101101011000100",
28653 => "110110101110111101011110",
28654 => "111010101000000001000010",
28655 => "111110010010000011001111",
28656 => "000010010101110010010011",
28657 => "000110011001100101110110",
28658 => "001001001100010110011111",
28659 => "001011000010100000011110",
28660 => "001101010111011010001110",
28661 => "001111110110001000100010",
28662 => "010000101000111101010000",
28663 => "001111011010101110000000",
28664 => "001101011011110100010100",
28665 => "001011011110110001000001",
28666 => "001010000001101110001011",
28667 => "001001101101010011000100",
28668 => "001010010100011100100111",
28669 => "001011001011000110000000",
28670 => "001100011011100000001110",
28671 => "001110011001010100101000",
28672 => "010000011110110101000100",
28673 => "010001111010111101010010",
28674 => "010010100110101101110010",
28675 => "010010110101101000000010",
28676 => "010010000111011111111110",
28677 => "001111100111010000111100",
28678 => "001101001000011011111110",
28679 => "001101000111001010110010",
28680 => "001101100111110000011110",
28681 => "001100000101001111001010",
28682 => "001010001011010001100101",
28683 => "001001110100000011000100",
28684 => "001010110000000101110100",
28685 => "001100100000111001010110",
28686 => "001110000010000011100110",
28687 => "001110101001110100001110",
28688 => "001110111011101101101010",
28689 => "001110001000010111111110",
28690 => "001010100011000010000010",
28691 => "000011101011010110010010",
28692 => "111010011101001100110001",
28693 => "110001000100101010001000",
28694 => "101001100000111101101010",
28695 => "100100100010111011011011",
28696 => "100010001011000111101111",
28697 => "100001011010010100001011",
28698 => "100001011000000101011001",
28699 => "100001101110000101001101",
28700 => "100001100100011001111011",
28701 => "100010011000000110010010",
28702 => "100111011111011111111110",
28703 => "110000001010110001011100",
28704 => "111001011011000100111101",
28705 => "000010000010110100110000",
28706 => "000111101111100010000111",
28707 => "001001000101000111001101",
28708 => "001000111001000011011011",
28709 => "001000100111110100110001",
28710 => "000110010010011101001000",
28711 => "000010010101000111000000",
28712 => "111111101010000100000101",
28713 => "111111000111110111010010",
28714 => "111111010111000010000010",
28715 => "111111010000100001100100",
28716 => "111111101000001111100100",
28717 => "000010010110101001011101",
28718 => "000110111100100110000111",
28719 => "001010011011010101000101",
28720 => "001011010110001010101100",
28721 => "001010001000100101101001",
28722 => "000111000110101001011100",
28723 => "000011011111111100000001",
28724 => "000000101000110001100111",
28725 => "111101111101001001110000",
28726 => "111011111010001101100000",
28727 => "111100100000111111110101",
28728 => "111111010100010001011100",
28729 => "000010010010111101011111",
28730 => "000100101010110100001000",
28731 => "000101011100101000010001",
28732 => "000011101111111110100111",
28733 => "000001010011101111000101",
28734 => "000000101000110011101010",
28735 => "000001010010101111001000",
28736 => "000000111110100111101100",
28737 => "111111010111100101011111",
28738 => "111101110000100000111110",
28739 => "111100100100010110010110",
28740 => "111100000001000011111001",
28741 => "111100101010101101000111",
28742 => "111110010000000011000111",
28743 => "000000000010101101000110",
28744 => "000001001000001100111000",
28745 => "000000011101110100010000",
28746 => "111110010111100101000100",
28747 => "111011100010101110110100",
28748 => "110111001100010001100000",
28749 => "110001000111110111101000",
28750 => "101011000011111111101010",
28751 => "100110010101001110101011",
28752 => "100011001111101000010011",
28753 => "100010000010101000111111",
28754 => "100010011100101101001000",
28755 => "100100001001110011111001",
28756 => "100111110101101100000111",
28757 => "101101111100110101111010",
28758 => "110101101100100011001111",
28759 => "111110001001000100110000",
28760 => "000110100000111110001000",
28761 => "001101101000011101101110",
28762 => "010010001011000011101110",
28763 => "010011000111101011000110",
28764 => "010000100101100100110100",
28765 => "001100001100110001000010",
28766 => "000111001011000101011000",
28767 => "000001011011111001001011",
28768 => "111011110100011000101000",
28769 => "111000010100010011011110",
28770 => "110111011001100000100010",
28771 => "110111111001110000010010",
28772 => "111001011001011010110010",
28773 => "111011111101000101110100",
28774 => "111111001000100001101011",
28775 => "000011001100010000010010",
28776 => "001000001010000001101100",
28777 => "001011111110101001111111",
28778 => "001101101100000010101100",
28779 => "001110111001010000101000",
28780 => "001111101111110001000110",
28781 => "001110110110011000111100",
28782 => "001100010010110111101110",
28783 => "001000111001011110100111",
28784 => "000101011101001111111000",
28785 => "000010110011101101110101",
28786 => "000000011100111001010100",
28787 => "111101001111100011010101",
28788 => "111001010101100000110110",
28789 => "110101111011010100100000",
28790 => "110011101001110101001010",
28791 => "110001101110110110100010",
28792 => "101111110001000011011110",
28793 => "101110111010011011110110",
28794 => "101111001101000111101010",
28795 => "101111001011100110011000",
28796 => "101110100101111100011110",
28797 => "101101111001011011100110",
28798 => "101101001010000000100110",
28799 => "101101000000100100110110",
28800 => "101110000100011010011100",
28801 => "101111101000001011000110",
28802 => "110000110010000010110000",
28803 => "110010010000111001010010",
28804 => "110101000101100100011110",
28805 => "111000000000001100100010",
28806 => "111001110101010010011100",
28807 => "111100000100101110001100",
28808 => "111111010110110011010101",
28809 => "000001100101101101111010",
28810 => "000001100010100010111000",
28811 => "000000001010000110011100",
28812 => "111110101111011110000111",
28813 => "111101110010010110001101",
28814 => "111101001010110101110110",
28815 => "111101000001011110111000",
28816 => "111101101010001100011010",
28817 => "111111010111010011011010",
28818 => "000010100101001101101011",
28819 => "000110110001101100110100",
28820 => "001010110010010101110101",
28821 => "001110110011001001011100",
28822 => "010011001001001100001110",
28823 => "010110101110110000100110",
28824 => "011000110100101111100100",
28825 => "011010000010000010100001",
28826 => "011010110100110010100101",
28827 => "011010110011100000100010",
28828 => "011010000101011101010001",
28829 => "011001101010100111000111",
28830 => "011001010110110011011001",
28831 => "011000011101110000011101",
28832 => "011000010100001001001001",
28833 => "011001101011010001100101",
28834 => "011010011100010000010001",
28835 => "011001010001001001010111",
28836 => "010111001011110010010000",
28837 => "010100100011110011111110",
28838 => "010000100001001010110000",
28839 => "001011001110000001010000",
28840 => "000110011000011101001110",
28841 => "000011001110101000010111",
28842 => "000000110101001111001000",
28843 => "111101010111110110110110",
28844 => "111000101101110010110000",
28845 => "110100100000010110100000",
28846 => "110001110111010001011100",
28847 => "110000111110000001100000",
28848 => "110010010100101010010000",
28849 => "110101110011000001000010",
28850 => "111010001001001101011100",
28851 => "111110100000011001000010",
28852 => "000001101110010100100000",
28853 => "000010101001010111101111",
28854 => "000010101111101010011010",
28855 => "000011011111011000001000",
28856 => "000011000011100010010101",
28857 => "000000000110101111011011",
28858 => "111100011001010111010110",
28859 => "111001101110001100000000",
28860 => "111000000110010000100101",
28861 => "110111000000101010100110",
28862 => "110110111100111101100011",
28863 => "111001000010100001111100",
28864 => "111101001000010000000000",
28865 => "000010010101000101110100",
28866 => "001000100010111010100000",
28867 => "001110011110101001101110",
28868 => "010000010100011101101110",
28869 => "001100100100110111101010",
28870 => "000111100000010010001111",
28871 => "000101000011000011010010",
28872 => "000011011111101100011011",
28873 => "000000011111000100111101",
28874 => "111101010100010000001101",
28875 => "111011100110100100011001",
28876 => "111010111011101001001010",
28877 => "111010001001100111000011",
28878 => "111001010000101011011101",
28879 => "111001110101110000001010",
28880 => "111100001100011110110001",
28881 => "111111000100110110101011",
28882 => "000010100101000100011110",
28883 => "000110010110000011101100",
28884 => "001000110001011111101100",
28885 => "001010011100101010111110",
28886 => "001011101100101101111101",
28887 => "001010100001110010100100",
28888 => "001000000101101001111110",
28889 => "001000010001000111101101",
28890 => "001010100010001100011111",
28891 => "001010011110111110100001",
28892 => "000110000100001111110100",
28893 => "111111000011111011010100",
28894 => "111000010111011000110010",
28895 => "110100000000101000001101",
28896 => "110001110000111110001110",
28897 => "101110111111010111011000",
28898 => "101010100011001111000000",
28899 => "100110100101010101101111",
28900 => "100100010111111000101011",
28901 => "100011110010011111100011",
28902 => "100101001110010000010011",
28903 => "100111110110010100101101",
28904 => "101011100100000011111010",
28905 => "110010110111100111000100",
28906 => "111101001011010011100000",
28907 => "000110101001111110111101",
28908 => "001110000110101110101110",
28909 => "010011100011001010011010",
28910 => "010110000101011010101110",
28911 => "010101011100110110101110",
28912 => "010001010101000110100010",
28913 => "001010001110110000010011",
28914 => "000010011101011111010010",
28915 => "111011000000010111101011",
28916 => "110100000110001011111100",
28917 => "101111011000111000000110",
28918 => "101101000111101101000000",
28919 => "101011111110000001010000",
28920 => "101100001101111010000000",
28921 => "101110100111100001110110",
28922 => "110010111100011001011010",
28923 => "111001001111001100101001",
28924 => "000000111110000000100110",
28925 => "000111100110001000000110",
28926 => "001010110111010001110100",
28927 => "001011100001000000100110",
28928 => "001011100110010111011001",
28929 => "001011100001011000101010",
28930 => "001010101111111111110010",
28931 => "001001010100100000111000",
28932 => "000111001000011101001110",
28933 => "000011111100101010110100",
28934 => "000000001010110011110010",
28935 => "111100001010001001101110",
28936 => "111000000111111000100110",
28937 => "110101000101110101111010",
28938 => "110011111110100010000000",
28939 => "110100000001000010011000",
28940 => "110100000101001010000011",
28941 => "110100010111011011010110",
28942 => "110101000101101000100100",
28943 => "110101011111101110110010",
28944 => "110101010100110000011100",
28945 => "110100110110010011110101",
28946 => "110011101001100100001110",
28947 => "110001101000101010111000",
28948 => "101111111010100111101010",
28949 => "101111000110011100010000",
28950 => "101110110111110010100100",
28951 => "101111101011111100000110",
28952 => "110010100010111101010000",
28953 => "110111010000001110101001",
28954 => "111100100001000001010100",
28955 => "000001001111000001110001",
28956 => "000100111011001011110111",
28957 => "000111000110110100011111",
28958 => "000111000010111011100101",
28959 => "000100111011011111010101",
28960 => "000001110111101010001101",
28961 => "111110000010011010110111",
28962 => "111001101001100110001011",
28963 => "110110011111010010111010",
28964 => "110101001100000011100100",
28965 => "110100100110000111010010",
28966 => "110100110110011101101001",
28967 => "110110111011010011110111",
28968 => "111010111011011000111101",
28969 => "000000011000101111001010",
28970 => "000101111010000010111011",
28971 => "001010010000000110110110",
28972 => "001101101100110011000000",
28973 => "010000001101001000000110",
28974 => "010001000111100011110010",
28975 => "010000101111000110111100",
28976 => "001111101101101000111000",
28977 => "001110110111111001100010",
28978 => "001111001001110111001000",
28979 => "010000010110000100011010",
28980 => "010001011111010110001100",
28981 => "010001101001011011111000",
28982 => "010000001110001101110010",
28983 => "001101111010001100101110",
28984 => "001011011010010110100000",
28985 => "001000000110010010110000",
28986 => "000100000110000111000010",
28987 => "000000111011100001110111",
28988 => "111111000010010010001010",
28989 => "111101000110010001111110",
28990 => "111010001001101101111010",
28991 => "110110101010100010101100",
28992 => "110011010100000010100110",
28993 => "110001000001000100101010",
28994 => "110001110001110110001100",
28995 => "110110010110111100010010",
28996 => "111100111100000101000000",
28997 => "000011101101000001100101",
28998 => "001001110111110001001010",
28999 => "001110100011101001110010",
29000 => "010000101010011111111010",
29001 => "010000001110001111010010",
29002 => "001111001101010000111010",
29003 => "001110111001101011100000",
29004 => "001110100001101110110110",
29005 => "001110010100010111100010",
29006 => "001110101111110101010010",
29007 => "001110001100111001010110",
29008 => "001100000100111111110100",
29009 => "001001100000110011101100",
29010 => "000111100101011011111110",
29011 => "001000001001110000101010",
29012 => "001011100010111111110101",
29013 => "001111001000101010110010",
29014 => "010001001100100001000110",
29015 => "010000111100111011001010",
29016 => "001101101000110111100000",
29017 => "001000111101010111111010",
29018 => "000100110000010001111010",
29019 => "000000011110000111101100",
29020 => "111100100011110001010100",
29021 => "111010001100011011110011",
29022 => "110111100110010110100000",
29023 => "110010011001001011000000",
29024 => "101011101001100000010100",
29025 => "100110000100111101010111",
29026 => "100011000100011101110010",
29027 => "100011100110110100000110",
29028 => "101000000001101100001010",
29029 => "101110001110010101010000",
29030 => "110100011011001100000111",
29031 => "111011000110110011010111",
29032 => "000001011101000011000100",
29033 => "000101010101110101110110",
29034 => "000110011110100000000100",
29035 => "000101100011101110101101",
29036 => "000011110000001000111001",
29037 => "000011010000001010001111",
29038 => "000100000101000100011111",
29039 => "000011001010011001101010",
29040 => "111111010000110100100111",
29041 => "111010001111000100100011",
29042 => "110101010011010001111011",
29043 => "110001010000001101001100",
29044 => "101111100010110101000000",
29045 => "101111011001110100110000",
29046 => "101110111101100010000100",
29047 => "101110010100011100011010",
29048 => "101101001100001111010110",
29049 => "101011110010000010110100",
29050 => "101101001001000011011110",
29051 => "110001111100011000000000",
29052 => "111000000000000001110101",
29053 => "111111101100111110110100",
29054 => "001001100000000100101000",
29055 => "010011010010100011110010",
29056 => "011010111100101101010010",
29057 => "011110101000001101000110",
29058 => "011110100011111011000111",
29059 => "011101001011001010110011",
29060 => "011001111011001110100101",
29061 => "010011110100100110000100",
29062 => "001101111110110111011110",
29063 => "001001101001101010011010",
29064 => "000100100000010110011000",
29065 => "111111010101100001100111",
29066 => "111100100110101111011010",
29067 => "111011010111100010011100",
29068 => "111010010111000110100100",
29069 => "111010011100111010100010",
29070 => "111011010111110111001111",
29071 => "111100011101100001101110",
29072 => "111111001111010110011000",
29073 => "000011101101001110000111",
29074 => "000111011101011001110110",
29075 => "001010110000000010101101",
29076 => "001111000001101110000010",
29077 => "010011010000110010011100",
29078 => "010110101000000010111000",
29079 => "011000100110010010100010",
29080 => "010110111000101000111010",
29081 => "010000011011011100101100",
29082 => "000110110111010101111011",
29083 => "111100010100011011101010",
29084 => "110010111110110011110010",
29085 => "101100100100010001000000",
29086 => "101001001110100101101000",
29087 => "101000010000001100101110",
29088 => "101000111001000110100010",
29089 => "101010110010010110100000",
29090 => "101101111110011110000100",
29091 => "110001110100101100001100",
29092 => "110101001011101100011001",
29093 => "110111110011011101101101",
29094 => "111001101001100001001101",
29095 => "111010000001011000001101",
29096 => "111001010111111000101000",
29097 => "111001001011010101101111",
29098 => "111000111011110100101001",
29099 => "110111101100100010000111",
29100 => "110111011110100001010100",
29101 => "111010001010101101000100",
29102 => "111110001110110100010011",
29103 => "000001110110001111011110",
29104 => "000101000011010001011110",
29105 => "000111011001010010111010",
29106 => "000111010110111001110000",
29107 => "000100101101100010100001",
29108 => "000000101111101110101000",
29109 => "111100010101100101111110",
29110 => "111000011001010001001110",
29111 => "110110010010100000011100",
29112 => "110101101000010111000100",
29113 => "110101010001111010110110",
29114 => "110110010101101110111101",
29115 => "111001110010001110001010",
29116 => "111101111111001010000100",
29117 => "000001101110111010001110",
29118 => "000110000001100111001000",
29119 => "001011001011100110110100",
29120 => "001111001110110011010010",
29121 => "010000110111011010001010",
29122 => "010001010011100010111100",
29123 => "010001100010001100001010",
29124 => "010000101100110010001110",
29125 => "001110001011101010011000",
29126 => "001011000011100100011101",
29127 => "001001001001011010101000",
29128 => "001000001111100100101110",
29129 => "000101100111011010000100",
29130 => "000000001010100011111100",
29131 => "111001111011011000100001",
29132 => "110101001000110110100010",
29133 => "110010100101011111011000",
29134 => "110001011000001000011000",
29135 => "110000100011010011110010",
29136 => "110000111001100101010110",
29137 => "110001111101111101110100",
29138 => "110000110100011100110000",
29139 => "101101000110010000000010",
29140 => "101010011100110010110000",
29141 => "101011010101101000011110",
29142 => "101110001000110100001100",
29143 => "110000111010000011111100",
29144 => "110100101001001001011010",
29145 => "111001100101110000000101",
29146 => "111101010001111111010100",
29147 => "111110111110111001110100",
29148 => "000000100110110110110101",
29149 => "000011100010101101100110",
29150 => "000111001110010101110000",
29151 => "001001110010110000001110",
29152 => "001011011001011110001011",
29153 => "001101101010001010001010",
29154 => "001110101110011000101000",
29155 => "001100100010101111110110",
29156 => "001001110010111110011010",
29157 => "001001010110000101101101",
29158 => "001011010110000000110110",
29159 => "001111000100100111110110",
29160 => "010010110010111101000100",
29161 => "010101000100001000101010",
29162 => "010110000101110000101010",
29163 => "010110000010110011011010",
29164 => "010100011001111101011010",
29165 => "010001001101001100000000",
29166 => "001110001100000101001100",
29167 => "001101000100101101011100",
29168 => "001100011110100101111100",
29169 => "001010011000000101011001",
29170 => "000111000110111100011100",
29171 => "000010111110101001001011",
29172 => "111110000000101010000101",
29173 => "111001111110000110111001",
29174 => "111000110000111101010101",
29175 => "111010010111111111001100",
29176 => "111101001011101100010100",
29177 => "111111110001111011111010",
29178 => "000001111001111111110011",
29179 => "000011011000110111000000",
29180 => "000011111001111110011100",
29181 => "000011000011110110100110",
29182 => "000000111011100001011010",
29183 => "111111010001011000100111",
29184 => "111110001000101101010001",
29185 => "111011010001110110101011",
29186 => "111000001101101111111110",
29187 => "110110101011010011011110",
29188 => "110011001110100111011110",
29189 => "101101001110100110011100",
29190 => "101000010000110011111000",
29191 => "100100110000011000010111",
29192 => "100010101100000011011111",
29193 => "100011000110110011010001",
29194 => "100100000000000101110101",
29195 => "100100000000101010011010",
29196 => "100100010110000011100000",
29197 => "100101011010001001100011",
29198 => "101000101100100100101100",
29199 => "101111101101001011011110",
29200 => "110111101101100010001000",
29201 => "111110111000011001010011",
29202 => "000111010100010001101110",
29203 => "010000000100101110011000",
29204 => "010101010010100010011010",
29205 => "010111000011100101111100",
29206 => "010110111111111111011110",
29207 => "010100010001011110001010",
29208 => "001111011000100000001100",
29209 => "001010010001101010111100",
29210 => "000101000101000101100001",
29211 => "000000110100011000101010",
29212 => "111111000101110111000110",
29213 => "111110001111010101100100",
29214 => "111101100000111011110010",
29215 => "111111010000001010111101",
29216 => "000010110100110010000110",
29217 => "000101010111011100110010",
29218 => "000111000001000010000000",
29219 => "001000110110101011110110",
29220 => "001010101111000110001000",
29221 => "001100101110110010000100",
29222 => "001110011000110110101110",
29223 => "001111001011010000011000",
29224 => "010000010111010000011010",
29225 => "010010011010110100110110",
29226 => "010011010111010000111000",
29227 => "010010001101001010010010",
29228 => "001111011110010111010010",
29229 => "001011000101001001011110",
29230 => "000101101001001001110110",
29231 => "000000100101011101110010",
29232 => "111011100000011000000111",
29233 => "110101011110111010110110",
29234 => "101111101101011111111010",
29235 => "101011111111001101001100",
29236 => "101010100100101010111100",
29237 => "101010101011110110101010",
29238 => "101011111100111110110100",
29239 => "101110011100001111100110",
29240 => "110001011000011010111010",
29241 => "110011101001101111101110",
29242 => "110101011000001111100010",
29243 => "110110111100111101000110",
29244 => "110111101010000100000001",
29245 => "110111001101110010010010",
29246 => "110110101110101101001000",
29247 => "110110101011100111001000",
29248 => "110110100101100010101101",
29249 => "110110110100010000000000",
29250 => "110111010010000110100010",
29251 => "110110100111000000010110",
29252 => "110101111000000111100110",
29253 => "110111110011010111010010",
29254 => "111011001001101100011100",
29255 => "111100110100100100010010",
29256 => "111101100000101010011011",
29257 => "111111100110000101110011",
29258 => "000010100101110000000011",
29259 => "000100010101100101001101",
29260 => "000100101010110001100000",
29261 => "000101000100010010110111",
29262 => "000101101010001110101000",
29263 => "000101110001001010110110",
29264 => "000101110111001101111000",
29265 => "000110010110001001000011",
29266 => "000110111110010000011111",
29267 => "000111110011101000110000",
29268 => "001001000011000000111100",
29269 => "001011000101001010100000",
29270 => "001101111110010111100110",
29271 => "010000100111000010100100",
29272 => "010010010100001110110100",
29273 => "010011101111101101011000",
29274 => "010100111111001010010100",
29275 => "010101000001111001111010",
29276 => "010011010110010101101100",
29277 => "010000101101010010110110",
29278 => "001101101010111100011110",
29279 => "001001010101011100110111",
29280 => "000011010110111011001111",
29281 => "111101101000001011010011",
29282 => "111010000100101110111100",
29283 => "111000000101101110011000",
29284 => "110101000111110110101010",
29285 => "101111111111100000111100",
29286 => "101010011001110001000010",
29287 => "100110100010010111001010",
29288 => "100101100110010101001011",
29289 => "100111111111110000000001",
29290 => "101100110111010001100010",
29291 => "110011001001100111111110",
29292 => "111010001001111010011011",
29293 => "000000000100100110000110",
29294 => "000011010110100101100001",
29295 => "000100011110110010110011",
29296 => "000100101001000111001010",
29297 => "000101000001011100101100",
29298 => "000110011000001110010101",
29299 => "000111111001010001011010",
29300 => "001000010110010000010110",
29301 => "000111110111100001100100",
29302 => "000111010100111101100100",
29303 => "000110111110011111100110",
29304 => "000110100111100110101101",
29305 => "000110100100000011010010",
29306 => "000111100010000001111100",
29307 => "001010001000110111100010",
29308 => "001101010110101111110110",
29309 => "001101111001000110100010",
29310 => "001011010101110111101000",
29311 => "001010000100101011100110",
29312 => "001011011010011011101011",
29313 => "001100000000010010010000",
29314 => "001010110010000111010100",
29315 => "001001100111101111000001",
29316 => "001001111011100001101101",
29317 => "001011000011101001100000",
29318 => "001001110101011010010010",
29319 => "000100100100010101101111",
29320 => "111101101001010110011110",
29321 => "111000010011001101111110",
29322 => "110110011100001000111010",
29323 => "110110111110000000101110",
29324 => "110110101100100111011100",
29325 => "110110101010001000010111",
29326 => "111001111111011110000001",
29327 => "111110000011011000001010",
29328 => "111111000000010101110011",
29329 => "111110100010100100101000",
29330 => "111111010011000111100011",
29331 => "000001001111101000101111",
29332 => "000011101010111100111100",
29333 => "000101000000000000100000",
29334 => "000011100100001001000001",
29335 => "000001001101110111110111",
29336 => "000000111111001001011000",
29337 => "000001111111101001111000",
29338 => "000010001001111001100101",
29339 => "000001001001110000100001",
29340 => "111110010010011010111011",
29341 => "111010010111100100000101",
29342 => "110111110010101000111010",
29343 => "110100111000110010010101",
29344 => "101111010101111000111100",
29345 => "101001101101111101100000",
29346 => "100110100111000101100111",
29347 => "100110111100111100010101",
29348 => "101011110010001010100100",
29349 => "110011010000110000110010",
29350 => "111011000011110010011010",
29351 => "000011111100011111010110",
29352 => "001100100110111010110110",
29353 => "010000110111001010011100",
29354 => "010000000001010101110100",
29355 => "001100111111001110000000",
29356 => "001001100010111101001000",
29357 => "000101000011110110100100",
29358 => "111110110000101101100011",
29359 => "111000010111110010111111",
29360 => "110101000101001110011000",
29361 => "110101010100001010110010",
29362 => "110110011111000100011101",
29363 => "111000010110111111111000",
29364 => "111101001101011010001011",
29365 => "000011011000100001010110",
29366 => "000111001000010000001011",
29367 => "001000111001001010100010",
29368 => "001001101111100001101000",
29369 => "001000110100101001011010",
29370 => "000111011101000011101011",
29371 => "000111000000101101101010",
29372 => "000110000100101101010000",
29373 => "000100001110001001011110",
29374 => "000010110100001101101101",
29375 => "000010010001000100101111",
29376 => "000001100011011010111010",
29377 => "111111011101101101111010",
29378 => "111100101111100101011000",
29379 => "111011001100010110000011",
29380 => "111010010001101101011000",
29381 => "111000101010111110101000",
29382 => "110110111001001111001101",
29383 => "110101100110010110100100",
29384 => "110100111000100111100110",
29385 => "110101000001011110110101",
29386 => "110101110100001100011000",
29387 => "110110111110111001011101",
29388 => "111000110110011000010110",
29389 => "111011010000110011010110",
29390 => "111100111101101111011011",
29391 => "111101000000111001100101",
29392 => "111011110100111001100010",
29393 => "111010001011001110001000",
29394 => "111000101111110101110011",
29395 => "111000001111011000110110",
29396 => "111000011011010110010000",
29397 => "111000110100000111001111",
29398 => "111001100011000011000010",
29399 => "111010001011010111010010",
29400 => "111010001110110011110011",
29401 => "111010101010100111100110",
29402 => "111100001110111000110000",
29403 => "111110011001000011100111",
29404 => "000000011100001110111101",
29405 => "000010001101100001110001",
29406 => "000100010001100101111100",
29407 => "000110100010011100111100",
29408 => "000111100001111100000100",
29409 => "000111010010101011000110",
29410 => "000111000011000110011101",
29411 => "000110001100110000010111",
29412 => "000100011010111100011111",
29413 => "000011000111110101111001",
29414 => "000010001010000011101110",
29415 => "000000000100111101101100",
29416 => "111101111101111000110100",
29417 => "111101101001110111001110",
29418 => "111110000011010011010110",
29419 => "111110111010100111111000",
29420 => "000010100000011110000111",
29421 => "001000010000101001000101",
29422 => "001101100100111101011010",
29423 => "010001100110111001011110",
29424 => "010011100111101101110000",
29425 => "010011001001101011010010",
29426 => "010000111110011011110000",
29427 => "001101001011101111001110",
29428 => "000111111001010101011000",
29429 => "000010000100100110010011",
29430 => "111011111111011011110001",
29431 => "110110001100010101110000",
29432 => "110001001110000000101100",
29433 => "101011111110011100011000",
29434 => "100110100100000111011001",
29435 => "100011010010011111000101",
29436 => "100011101101001110010101",
29437 => "101000000110110000000100",
29438 => "101111100011010100101100",
29439 => "111000000101111110111001",
29440 => "000000010000011000101100",
29441 => "000110011111110100011110",
29442 => "001000111011010011010001",
29443 => "001000000011010110100001",
29444 => "000110111111100110100111",
29445 => "000111010000011001111010",
29446 => "000111101000100111100100",
29447 => "000111010001110111111100",
29448 => "000110011110000011111010",
29449 => "000101010110101011010011",
29450 => "000011110110111110100110",
29451 => "000010101101101101101110",
29452 => "000010111010010000000000",
29453 => "000100000011110110100111",
29454 => "000101110100111000010101",
29455 => "001000011001100111000100",
29456 => "001010001001001111101100",
29457 => "001001000110000101110010",
29458 => "000110001101101011110010",
29459 => "000100000101000010001111",
29460 => "000011011111011110101110",
29461 => "000011110000100010000000",
29462 => "000100101001100110011010",
29463 => "000101011011100010000111",
29464 => "000100110000010010101101",
29465 => "000010001111100011110011",
29466 => "111101111110011011010111",
29467 => "111000100001110110010110",
29468 => "110011100001101001000100",
29469 => "101111111000101011000010",
29470 => "101101101010011001000010",
29471 => "101110000001000000001010",
29472 => "110000111100101111100110",
29473 => "110011100110100011101000",
29474 => "110101100010101100000100",
29475 => "111000111001001000000011",
29476 => "111100000010001110110111",
29477 => "111100110101110110101001",
29478 => "111110000111010011000000",
29479 => "000001011000000001100011",
29480 => "000011001010100101100011",
29481 => "000001111011110011111001",
29482 => "111111011000010101100000",
29483 => "111100011010001010110000",
29484 => "111010011100011101000101",
29485 => "111010011001100010000011",
29486 => "111010011000001011110100",
29487 => "111010000110111100001010",
29488 => "111011010110001011011001",
29489 => "111100110010010101110100",
29490 => "111100011011010100000000",
29491 => "111100000001100011000000",
29492 => "111100111100110010010001",
29493 => "111110000000100000101101",
29494 => "111111100100011010011111",
29495 => "000001111010101110011111",
29496 => "000100001110101001000111",
29497 => "001000010010001101100000",
29498 => "001110011011011110110110",
29499 => "010011100000101111110110",
29500 => "010111011100101010110010",
29501 => "011011101100011011110111",
29502 => "011110001010010110010011",
29503 => "011101111010100110101001",
29504 => "011100111011001001010001",
29505 => "011010100110011110100010",
29506 => "010110100100011001010110",
29507 => "010011010000011011001100",
29508 => "010000000100011101000100",
29509 => "001100011101000011001100",
29510 => "001011010100010101010111",
29511 => "001011011101111110111111",
29512 => "001010000111111000010000",
29513 => "001001100001001110110000",
29514 => "001010000111100011000010",
29515 => "001000110110011101011000",
29516 => "000110001000101100101100",
29517 => "000100000010000000100001",
29518 => "000010110111010010101101",
29519 => "000010111000101111111110",
29520 => "000010101111010110100001",
29521 => "000000001100000000011011",
29522 => "111100001000111100010110",
29523 => "111001000000110111000001",
29524 => "110111100100000010000110",
29525 => "110111001110010011101001",
29526 => "110111100001000000110100",
29527 => "111000001000000011000011",
29528 => "111000110100110110100111",
29529 => "111001111001111110001000",
29530 => "111010100111111111000111",
29531 => "111001101001110100110100",
29532 => "110111100111001000100010",
29533 => "110110000101010000000011",
29534 => "110101101011000000100001",
29535 => "110101010000110110001110",
29536 => "110100000110100100110101",
29537 => "110011101101100101001110",
29538 => "110011111111100001001000",
29539 => "110010011100111111000010",
29540 => "101111000010100101000000",
29541 => "101100011010111100111000",
29542 => "101100000000111001000110",
29543 => "101101000100111100101010",
29544 => "101111100000110000000110",
29545 => "110011011000010010001110",
29546 => "110110110110100111011110",
29547 => "111001010111101100111100",
29548 => "111100100110101111011001",
29549 => "000000011100100011101000",
29550 => "000011110100001111011101",
29551 => "000111100000100011011000",
29552 => "001011011010001100001111",
29553 => "001110001101010001101000",
29554 => "010000010010100110011000",
29555 => "010001011000110111100100",
29556 => "010000001100000101010100",
29557 => "001100110000011001011010",
29558 => "001000000000000110010000",
29559 => "000100100001001111111001",
29560 => "000011101110101011011110",
29561 => "000010100000101001001101",
29562 => "111111100100011001100100",
29563 => "111101010100101101100010",
29564 => "111011111011011100010011",
29565 => "111010111101111000000010",
29566 => "111100000111000001101110",
29567 => "111110101011011010011101",
29568 => "000001000010000110000011",
29569 => "000101001010010011110100",
29570 => "001011100010110011110011",
29571 => "010000111011010011100010",
29572 => "010100100011111100000110",
29573 => "010111010011011100100000",
29574 => "010111011011010010100100",
29575 => "010100000001100000111000",
29576 => "001110110010010111100100",
29577 => "001000011010011011011101",
29578 => "000000111011100110001010",
29579 => "110111110100111111001010",
29580 => "101100001110100111011010",
29581 => "100011000110000100101011",
29582 => "100001001010100000101011",
29583 => "100001100110101001111000",
29584 => "100000111011011001010001",
29585 => "100001000000011111101100",
29586 => "100010101011000011000111",
29587 => "101000100111011101000010",
29588 => "110010111001101011111010",
29589 => "111100000010111010101110",
29590 => "000010101011011110111101",
29591 => "000111111111010010000100",
29592 => "001011001111111000010011",
29593 => "001101100110100110110100",
29594 => "001110111011110010110010",
29595 => "001101001000010111001110",
29596 => "001010000110001010011000",
29597 => "000111100010110100110010",
29598 => "000011111011111010000000",
29599 => "000000001111100110100100",
29600 => "111110101101100101011101",
29601 => "111111110111100010100000",
29602 => "000011001100100001100101",
29603 => "000110010001101101010111",
29604 => "000111100001001000011111",
29605 => "001000011100001100000010",
29606 => "001010011000100110000000",
29607 => "001100000100011101100000",
29608 => "001011100101100100110011",
29609 => "001001111111111010111000",
29610 => "001001110000000100100001",
29611 => "001010010100001110111001",
29612 => "001000111010101001000100",
29613 => "000100000101001010010111",
29614 => "111101010010000010011111",
29615 => "110111010001010001001010",
29616 => "110010111101100000011010",
29617 => "101111000111101000110000",
29618 => "101011110101100010010000",
29619 => "101011000010110001110000",
29620 => "101100101101111110100000",
29621 => "101111011001100110111010",
29622 => "110001110100110010101110",
29623 => "110011001010100111101110",
29624 => "110100100101001101000100",
29625 => "110110101101100010010101",
29626 => "111000101101111111111101",
29627 => "111010011000111110110000",
29628 => "111010100110000010001110",
29629 => "111000100000101100000010",
29630 => "110101011000100101000000",
29631 => "110010000110100000010100",
29632 => "101110100001010101100100",
29633 => "101011010010011111011110",
29634 => "101010101110000100000010",
29635 => "101101011001011100111110",
29636 => "110000100001111011000010",
29637 => "110010010001010110111100",
29638 => "110010110000011010101110",
29639 => "110010101010000001111000",
29640 => "110011011101101011100010",
29641 => "110101000101101101000111",
29642 => "110101111000100000101011",
29643 => "110111011001010101100001",
29644 => "111011101010010011110110",
29645 => "000000010111010100011101",
29646 => "000100010010011101000010",
29647 => "001000110001101100000100",
29648 => "001100111111111111011010",
29649 => "010000011101001010110000",
29650 => "010011101110001111011010",
29651 => "010101101101011110011100",
29652 => "010110000100110011011110",
29653 => "010101111101101011111110",
29654 => "010101001111101010011110",
29655 => "010011011111010001111010",
29656 => "010001101110101100111100",
29657 => "001111110100011110101110",
29658 => "001101100100000000111100",
29659 => "001101101001101110011100",
29660 => "001111111110100001111010",
29661 => "010000111000110101100100",
29662 => "010000011010110100110110",
29663 => "010000100010010011001110",
29664 => "010000100000111110011010",
29665 => "001111100011010111000110",
29666 => "001110010110011000011100",
29667 => "001100100110011010000010",
29668 => "001010101001011000011011",
29669 => "001010011000100101001110",
29670 => "001010000011111101100011",
29671 => "000111000010000011001111",
29672 => "000011000110111011010100",
29673 => "000000010001110101111010",
29674 => "111110101001110010011000",
29675 => "111110000101011011101011",
29676 => "111110000111110111010110",
29677 => "111110011100001011101010",
29678 => "111110110000010100111111",
29679 => "111110011111110101001110",
29680 => "111100011000101111101001",
29681 => "111000000110110101100110",
29682 => "110100000110111000010110",
29683 => "110010011100100101001010",
29684 => "110010010101010111001000",
29685 => "110001011101011011000100",
29686 => "101110101110110101010110",
29687 => "101011101101000110010110",
29688 => "101001011110110111111000",
29689 => "100111001101011110011101",
29690 => "100101110101110000100001",
29691 => "100111110100111001000010",
29692 => "101100100010100011001000",
29693 => "110001110000010101100010",
29694 => "110110101001100001010111",
29695 => "111010110011100011101110",
29696 => "111110110000111011000001",
29697 => "000010110111110010100100",
29698 => "000101111100100110001000",
29699 => "000111111111011100101000",
29700 => "001010000101111010101101",
29701 => "001100010111111110111010",
29702 => "001101100001101000011100",
29703 => "001100010011010100101110",
29704 => "001000110100100000010101",
29705 => "000011101001110000011110",
29706 => "111111001001100010000001",
29707 => "111101001011100001110011",
29708 => "111100100001010110110001",
29709 => "111101100001111001110100",
29710 => "000000110110001010111101",
29711 => "000100101011011010101000",
29712 => "001000001101010010111011",
29713 => "001011000101111101110111",
29714 => "001101010100101010100110",
29715 => "001111111101010000000110",
29716 => "010010111101010000110110",
29717 => "010101111110011001110000",
29718 => "011001001000000011001011",
29719 => "011011001100000011110111",
29720 => "011010101011011001100111",
29721 => "011000000111101000111101",
29722 => "010100100111101100010100",
29723 => "010000100100001000110010",
29724 => "001100100000011010000100",
29725 => "001001001100001010001111",
29726 => "000110101110111101111011",
29727 => "000011000100100000111000",
29728 => "111011111011001101001101",
29729 => "110010100100001101110100",
29730 => "101001110001001111101100",
29731 => "100100000010001100101001",
29732 => "100010111110000010110101",
29733 => "100101010101000010000001",
29734 => "101001011001011110011010",
29735 => "101111100100100100010110",
29736 => "111000010011000100100100",
29737 => "000001011001001001000100",
29738 => "001000000101000101110011",
29739 => "001100111111011000011010",
29740 => "010001111010111110000110",
29741 => "010110011000011010101010",
29742 => "011000101010111111111111",
29743 => "010111100010100000100110",
29744 => "010010110100001110001100",
29745 => "001011110110001000100010",
29746 => "000100110100101101110110",
29747 => "111110100100111110111101",
29748 => "111001011101001111111011",
29749 => "110110111000000001110100",
29750 => "110111001110111100100100",
29751 => "111001101100100110100110",
29752 => "111100010101010101001000",
29753 => "111101100100100110111000",
29754 => "111110111111011101000111",
29755 => "000010010011101111000110",
29756 => "000110110110011010011001",
29757 => "001010000111111010010110",
29758 => "001010011011000111101010",
29759 => "001001010000001101111110",
29760 => "000110111110001101000110",
29761 => "000011001100001110010110",
29762 => "111111011001001010110011",
29763 => "111010011010101011011110",
29764 => "110100000001101000101000",
29765 => "110000011010010100000110",
29766 => "110000100010110110101100",
29767 => "110001111101111000110110",
29768 => "110011100111101111000010",
29769 => "110100000011110011111010",
29770 => "110011000001011011101110",
29771 => "110011100000000100000000",
29772 => "110101011111101110100001",
29773 => "110110001111101010011001",
29774 => "110110101001011111011111",
29775 => "110111110000010100010001",
29776 => "110111010111000000001011",
29777 => "110100110011001010110010",
29778 => "110001111100101010000100",
29779 => "101111000010000110101100",
29780 => "101011101001110110110100",
29781 => "101001101110110101010010",
29782 => "101001110111000001000110",
29783 => "101010111110001010010010",
29784 => "101101011100101010111110",
29785 => "110000110000101001101000",
29786 => "110011111110000010000100",
29787 => "110111001010011100100110",
29788 => "111001110101000101000110",
29789 => "111100000010010011010111",
29790 => "111111000101001111111000",
29791 => "000011010100011000100100",
29792 => "000101110101000110100101",
29793 => "000100000000001101101001",
29794 => "000000001000011011100011",
29795 => "111100110101110000011010",
29796 => "111010011110100100111001",
29797 => "111001000101110001101110",
29798 => "111000101000101011000001",
29799 => "111010000011111000000011",
29800 => "111101011101001010001011",
29801 => "000001010111001110011111",
29802 => "000101101011110001100001",
29803 => "001010000110111101001001",
29804 => "001101000110000011010100",
29805 => "001110101100001100100010",
29806 => "001111110000000001110010",
29807 => "001111011011000001010110",
29808 => "001101101101111011011100",
29809 => "001100011000101111010010",
29810 => "001011000101100010101011",
29811 => "001000101001011101011010",
29812 => "000101101011100010100011",
29813 => "000011011101010100100010",
29814 => "000010111100010100100110",
29815 => "000011100011101110011110",
29816 => "000011101011001101111100",
29817 => "000010011111001101000111",
29818 => "000000100101011100100011",
29819 => "111110111001100111111100",
29820 => "111101010010111111100000",
29821 => "111100000011111100000000",
29822 => "111100011011000111100101",
29823 => "111110111100100101010100",
29824 => "000011000100111010011010",
29825 => "000111000110010010101111",
29826 => "001001100101010010010100",
29827 => "001010011100100001100100",
29828 => "001010001001110110001111",
29829 => "001000101000011110001010",
29830 => "000101100011101100110110",
29831 => "000001110101010001001111",
29832 => "111110010010111111000100",
29833 => "111011100010011011111011",
29834 => "111010000111110000101000",
29835 => "111000111001110010001101",
29836 => "110111111110011100110100",
29837 => "111001001010101111101110",
29838 => "111100010001010010000110",
29839 => "111111011100111011101110",
29840 => "000001011010000100100101",
29841 => "000010100101000100000101",
29842 => "000011001001000101011101",
29843 => "000010011110000010101111",
29844 => "000001101110010101101100",
29845 => "000001100110001101101001",
29846 => "000001100110111110010010",
29847 => "000010001001101000010110",
29848 => "000011010101101101010100",
29849 => "000100011011110001000110",
29850 => "000100101111011001110110",
29851 => "000100111111111100100010",
29852 => "000101010001101110001100",
29853 => "000010110001001111100111",
29854 => "111100111000100010110101",
29855 => "110110111100011101111101",
29856 => "110011000011001111001110",
29857 => "110001000001000101111100",
29858 => "110000110101010111100110",
29859 => "110010101011001010011000",
29860 => "110110001000101000010100",
29861 => "111010100010100100101010",
29862 => "111111011001011100010010",
29863 => "000101000100100001110010",
29864 => "001011001110101000011000",
29865 => "010000000011111101000110",
29866 => "010010111011011001010100",
29867 => "010100000111011011011000",
29868 => "010011101001111010100100",
29869 => "010001100000110111011010",
29870 => "001101111010100110110000",
29871 => "001001011001010101001001",
29872 => "000011011101011101010101",
29873 => "111101100111010100000111",
29874 => "111010011010000000110110",
29875 => "110111001110000101100001",
29876 => "110010000100011100000010",
29877 => "101101010110101101110100",
29878 => "101010000101110100010010",
29879 => "101000010111011010111100",
29880 => "101000111110011111001100",
29881 => "101100011101010010011010",
29882 => "110010001100001010110110",
29883 => "111000001101010100010010",
29884 => "111101110000010101111110",
29885 => "000011100010000000110110",
29886 => "001001100101100111110100",
29887 => "001111001010011001010100",
29888 => "010011111000001111001110",
29889 => "010111100011000100011010",
29890 => "011001010011000101011101",
29891 => "011000111011011100011001",
29892 => "010110111110001111100010",
29893 => "010011110110010001000100",
29894 => "001111110101100000010110",
29895 => "001011001001101110100000",
29896 => "000111011101111010110110",
29897 => "000101110100011111101000",
29898 => "000100001011000010000101",
29899 => "000000101111000110101101",
29900 => "111100011000001000101011",
29901 => "111001110110001001110110",
29902 => "111010101100000011001110",
29903 => "111101001100001111110010",
29904 => "000000000111011000111111",
29905 => "000101000010111011100100",
29906 => "001100000100100100101010",
29907 => "010001111101010111010100",
29908 => "010100111000011000110000",
29909 => "010101000110110011010110",
29910 => "010010111000011110011110",
29911 => "001111011011000001100100",
29912 => "001010111110000111100011",
29913 => "000100101100000111001100",
29914 => "111101101101011100010101",
29915 => "111000000010000110001010",
29916 => "110011110110000001010000",
29917 => "101110110001111010110100",
29918 => "101000011001100110110000",
29919 => "100011111000101011101001",
29920 => "100010100010010100001001",
29921 => "100011110000010001110001",
29922 => "100110111111010011001011",
29923 => "101010111000001000101100",
29924 => "101110001111101101000000",
29925 => "110000100101011101100000",
29926 => "110010001111010000110110",
29927 => "110011101100011001110110",
29928 => "110100111111000111000110",
29929 => "110110010010001000110000",
29930 => "110111101001000101011000",
29931 => "111001000110011111100000",
29932 => "111001100010110011110001",
29933 => "111000001010001010000010",
29934 => "110111010011101101100110",
29935 => "111000111111111000100100",
29936 => "111100011011011100111011",
29937 => "000000001110100100111010",
29938 => "000100000110001100110000",
29939 => "001000000101001000111000",
29940 => "001011001000010110100100",
29941 => "001100011001000110100000",
29942 => "001011010001101001100100",
29943 => "000111001010101110001000",
29944 => "000001110001001011111101",
29945 => "111101010100110100111001",
29946 => "111001110110100010010010",
29947 => "110111101100010100100010",
29948 => "111000011011111111000110",
29949 => "111011111111010000000010",
29950 => "000001011111000111000111",
29951 => "001000011010100110101101",
29952 => "001110110101010011001000",
29953 => "010011111001011001001110",
29954 => "011000001100000011101101",
29955 => "011010111101110001101010",
29956 => "011011101000111001100101",
29957 => "011001100010011110111111",
29958 => "010100011101000001110000",
29959 => "001110011001011001010010",
29960 => "001001001010100110101110",
29961 => "000100101110001110101101",
29962 => "000000001100000011110110",
29963 => "111100001001010011010010",
29964 => "111001001110001100101011",
29965 => "110110010010001010101110",
29966 => "110011111001011010111000",
29967 => "110010010101101111011010",
29968 => "110000011010001010011010",
29969 => "101111100111100010011000",
29970 => "110001000010111111110010",
29971 => "110011000000000101101010",
29972 => "110100101100101001100010",
29973 => "110111100101111100011010",
29974 => "111100011010101000110011",
29975 => "000000001000111001011101",
29976 => "000000000010010010001011",
29977 => "111101110100000100011100",
29978 => "111100001101100111011011",
29979 => "111011110000001100110101",
29980 => "111011000111010011101000",
29981 => "111001000101010000110001",
29982 => "110110100110001001110010",
29983 => "110101110100111101110000",
29984 => "110110110111010100101100",
29985 => "111000000111010101100010",
29986 => "111001010100100010111110",
29987 => "111011110001001111101101",
29988 => "000000001011110110000100",
29989 => "000011101111100010100010",
29990 => "000011110001001110101101",
29991 => "000011001111110000110110",
29992 => "000100010111100100101001",
29993 => "000100110101110111010100",
29994 => "000011110010011001110000",
29995 => "000011011000101001000101",
29996 => "000101110000010101011010",
29997 => "001001010110000011011010",
29998 => "001010111111010011100000",
29999 => "001011001110100100011010",
30000 => "001100010100000000011000",
30001 => "001110010010001100110010",
30002 => "001111110100110101111110",
30003 => "010000000111001111001110",
30004 => "001110101110001000000010",
30005 => "001100010000001111110000",
30006 => "001010010010000110111101",
30007 => "001000110011100101011000",
30008 => "000111010111111011001011",
30009 => "000110001101101011101101",
30010 => "000101001000110101010001",
30011 => "000100011101101100110010",
30012 => "000100100011000100001110",
30013 => "000101100100011111010000",
30014 => "000110100011001011100010",
30015 => "000101101100110010110000",
30016 => "000100001111101000010111",
30017 => "000011000011000100000011",
30018 => "000000111100010000100101",
30019 => "111110001111011111101001",
30020 => "111010001100100101101110",
30021 => "110100100000100101011101",
30022 => "101111011001111001100000",
30023 => "101010011101111001110110",
30024 => "100101000001101111010000",
30025 => "100010001000011011001011",
30026 => "100010011101101010001101",
30027 => "100011011001000011101101",
30028 => "100101101001010011010111",
30029 => "101011011001101101110110",
30030 => "110011011000001100111000",
30031 => "111010110000010001010111",
30032 => "111111100001011111111001",
30033 => "000001101010101110011101",
30034 => "000010110001110000011001",
30035 => "000100000101010001010010",
30036 => "000101110111100111001111",
30037 => "000111011010111101111110",
30038 => "001000000000010100111100",
30039 => "000111011001101100010001",
30040 => "000110010010111011110000",
30041 => "000110001011010010011000",
30042 => "000111000011001000001111",
30043 => "001000001111001111100010",
30044 => "001001100100110100001110",
30045 => "001010111011101001010110",
30046 => "001100010011000010010100",
30047 => "001100010101001001110000",
30048 => "001001111011001110101011",
30049 => "000110001101000101010010",
30050 => "000011100111111001011010",
30051 => "000100010000101100101011",
30052 => "000110101010110110011111",
30053 => "001001000010000111110100",
30054 => "001100010010111011000000",
30055 => "001111111101101000010110",
30056 => "010010010010010111000100",
30057 => "010010011000011000010110",
30058 => "010000110011101100101100",
30059 => "001111101111101001001100",
30060 => "001111010111010111111010",
30061 => "001110001001111011011100",
30062 => "001100010011011110010010",
30063 => "001010000000110110001100",
30064 => "000110000010100010111010",
30065 => "111111111000001100011010",
30066 => "111000010000111110101101",
30067 => "110000000111111011101000",
30068 => "101001011011100001010110",
30069 => "100110000001101100101111",
30070 => "100101001100001010001111",
30071 => "100101010100100101000111",
30072 => "100110000100100000100101",
30073 => "100111100111010001000011",
30074 => "101010000000000011110000",
30075 => "101110001101010110101110",
30076 => "110011111100010110000110",
30077 => "110111111110110110010010",
30078 => "111001100101010000001111",
30079 => "111010001000011111000111",
30080 => "111000101010110110110111",
30081 => "110100111100100011001001",
30082 => "110000100001100000000010",
30083 => "101100101010100001000100",
30084 => "101010101101011011111000",
30085 => "101100010100001110001000",
30086 => "110001111110101010111000",
30087 => "111001100101010001011110",
30088 => "000001000110001100111001",
30089 => "000111101110000011101100",
30090 => "001011011111000100011011",
30091 => "001011011000010111101111",
30092 => "001001000111010101011010",
30093 => "000101101101101011100001",
30094 => "000000000011000110000010",
30095 => "111000111000010101100111",
30096 => "110011100001001101011100",
30097 => "110001010110010001011100",
30098 => "110010010110011011010110",
30099 => "110110010111011110011101",
30100 => "111100101000110001100011",
30101 => "000101000011101101000110",
30102 => "001110101000101010101010",
30103 => "010111001101000100010100",
30104 => "011100101101101111101011",
30105 => "011110011001011111101001",
30106 => "011110001100010110010011",
30107 => "011011111100111000011000",
30108 => "010101001110100010100110",
30109 => "001100000111010101001000",
30110 => "000100010001001111011110",
30111 => "111101110100111110001001",
30112 => "110111111100001011000101",
30113 => "110010100110111111011110",
30114 => "101110110101001100111000",
30115 => "101101111001011010100010",
30116 => "101110100000111111110100",
30117 => "101110011100001000100010",
30118 => "101110011010101010101100",
30119 => "101111110110001101010110",
30120 => "110010111110101110010000",
30121 => "110111011001110111000010",
30122 => "111011000101000101000010",
30123 => "111101000100011001101011",
30124 => "111111000111110111110000",
30125 => "000010011001100010111011",
30126 => "000101001000000010100010",
30127 => "000101000010110111011111",
30128 => "000011101100000110111011",
30129 => "000010110101011111110111",
30130 => "000000110000000011111000",
30131 => "111100011000110001100110",
30132 => "110111001100000110011011",
30133 => "110011011111010111101010",
30134 => "110010010000110111010110",
30135 => "110010010110001000000100",
30136 => "110010110011011011001110",
30137 => "110011100000011011110100",
30138 => "110101000010000100111001",
30139 => "110111010111011000011000",
30140 => "111001000011100101111010",
30141 => "111001111111101100101101",
30142 => "111011001101010100110110",
30143 => "111101010000101001110000",
30144 => "000000000111001100010000",
30145 => "000011001110110011000011",
30146 => "000110111100010011010001",
30147 => "001011011100101000101110",
30148 => "001111110101000000000000",
30149 => "010011100101101000010010",
30150 => "010110100110000101011100",
30151 => "011000001011110101010011",
30152 => "010111101111000000001010",
30153 => "010101110010111111101010",
30154 => "010011001111001001011110",
30155 => "001111110011100101100010",
30156 => "001011010011001010011010",
30157 => "000111000110001000100100",
30158 => "000101000000011111101011",
30159 => "000101000001101001010000",
30160 => "000110010000011100110100",
30161 => "001000010111101111001011",
30162 => "001011010100101010110101",
30163 => "001111001111101110100000",
30164 => "010010101001111010111110",
30165 => "010011100000101110000110",
30166 => "010010011010000101011110",
30167 => "010000111000010100011010",
30168 => "001111011100011011011000",
30169 => "001101100000001101001110",
30170 => "001010100001001001001100",
30171 => "000110110000111010011111",
30172 => "000001101111101101100111",
30173 => "111011110101111100010010",
30174 => "110111101110010111100101",
30175 => "110111001111101001111111",
30176 => "111001011101100010001101",
30177 => "111100100100101111100100",
30178 => "000000100001111110000011",
30179 => "000100010000001000001000",
30180 => "000100110100111111000100",
30181 => "000011000000111101111001",
30182 => "000010000001101001001111",
30183 => "000010010011111000100111",
30184 => "000010101011001010100101",
30185 => "000010110100011001110100",
30186 => "000010110001110101011011",
30187 => "000010100110101011001111",
30188 => "000010000000010011110000",
30189 => "111111010110001011001101",
30190 => "111011011111100000111010",
30191 => "111010010100111101001010",
30192 => "111011111111000111100010",
30193 => "111101011110010111010111",
30194 => "111100100110110101111110",
30195 => "111001101001100010000100",
30196 => "111000110111001100101100",
30197 => "111011111011101111010000",
30198 => "111110110001000010111110",
30199 => "111111111101100011110100",
30200 => "000001111010110010111110",
30201 => "000100110100101100101000",
30202 => "000111011111111101110100",
30203 => "001001110001100001001000",
30204 => "001011000101101110101110",
30205 => "001010010010111110110110",
30206 => "000111000111111011001111",
30207 => "000011100001100111000010",
30208 => "000010011011011001000101",
30209 => "000100001100010011010000",
30210 => "000110100001011011011010",
30211 => "000111000010100010001111",
30212 => "000110011010010001011100",
30213 => "000110101001010011010110",
30214 => "000100110011011110011110",
30215 => "111110101000110000100110",
30216 => "111000011000010000111101",
30217 => "110100010111101111000010",
30218 => "110001011001001010110110",
30219 => "101110110001101101100110",
30220 => "101011110001111101100000",
30221 => "101001010101101100101100",
30222 => "101001100011100001100000",
30223 => "101011111011101100100110",
30224 => "101110010101110111000100",
30225 => "110001010011111001110110",
30226 => "110111001010010001101010",
30227 => "111101101101010011100101",
30228 => "111111110011100010000011",
30229 => "111101010111010110001001",
30230 => "111010011010101001011010",
30231 => "111000000011100011000101",
30232 => "110101000111111110000101",
30233 => "110010111000111110010110",
30234 => "110010101100011000110000",
30235 => "110100000010011010100111",
30236 => "110111011001001011110010",
30237 => "111101001100000110010101",
30238 => "000011111011000000100111",
30239 => "001001011011101001100111",
30240 => "001100001111001101100110",
30241 => "001100100011100111101100",
30242 => "001100011100111100100110",
30243 => "001100110111110011110010",
30244 => "001011000100010101111011",
30245 => "000100111011010100010010",
30246 => "111100110101000110110100",
30247 => "110101111000111001110100",
30248 => "110001011001110010001000",
30249 => "101111110000000110001010",
30250 => "110000011100011001110110",
30251 => "110011000100101111111010",
30252 => "111000010100010011110001",
30253 => "111111100000111100110000",
30254 => "000101111111110100101001",
30255 => "001011011101011011001011",
30256 => "010000111110000000001110",
30257 => "010101001011110101010100",
30258 => "010110110100110101100110",
30259 => "010101000010010011001010",
30260 => "001111010011110010110000",
30261 => "000111110100010111110010",
30262 => "000000001101011001101011",
30263 => "110111101000111101101101",
30264 => "101110110001010101010010",
30265 => "101000100011001000000010",
30266 => "100101111000010111010101",
30267 => "100101001010000011011011",
30268 => "100110001110110000011000",
30269 => "101001100100010001111000",
30270 => "101110101001101011101000",
30271 => "110101001010100101010001",
30272 => "111011100110100101011000",
30273 => "111111111110110101001000",
30274 => "000010101100000110010011",
30275 => "000101011101001111111100",
30276 => "001000010111010010000000",
30277 => "001001011110000001101100",
30278 => "001000001001100011110011",
30279 => "000110000110011001010001",
30280 => "000100001101100101011100",
30281 => "000001100011100000100100",
30282 => "111101110000101100100100",
30283 => "111010010001001001001110",
30284 => "111000001111000100101100",
30285 => "110111011011011101100001",
30286 => "110111001110101100101011",
30287 => "110111001001111000001101",
30288 => "110111100110101111010000",
30289 => "111001010100110101000000",
30290 => "111011010100010011010111",
30291 => "111011111100110000111100",
30292 => "111100010010100110010000",
30293 => "111110001110010000010111",
30294 => "000000100101111101110000",
30295 => "000010000001101001010000",
30296 => "000011000111111101011110",
30297 => "000100011100001100101111",
30298 => "000110001000011110000100",
30299 => "000111100010010100101101",
30300 => "001000000010110001000100",
30301 => "001000100001010010000110",
30302 => "001001001101000001001000",
30303 => "001000111010101111111011",
30304 => "000111000011111010110100",
30305 => "000100101000000000010000",
30306 => "000010010100010010111111",
30307 => "111111010110011010101111",
30308 => "111011110000010000110100",
30309 => "111000101010010001111001",
30310 => "110110110010001010000000",
30311 => "110110001100000110110111",
30312 => "110110100100110111011001",
30313 => "111000001011001100110010",
30314 => "111011000110110101000101",
30315 => "111110101101111101011000",
30316 => "000010000011010100111101",
30317 => "000011110100011110001010",
30318 => "000011011110001101110010",
30319 => "000001000110001011111100",
30320 => "111100110110100001101101",
30321 => "111000101001000100001110",
30322 => "110111010001111110111010",
30323 => "111001000101000110100001",
30324 => "111011110000011010101000",
30325 => "111110000010010100101010",
30326 => "000000101111001110110001",
30327 => "000100001000001111000001",
30328 => "000111101000100110100110",
30329 => "001011000111001010111001",
30330 => "001101111011101101011000",
30331 => "001111011000110101101100",
30332 => "010000001100101001111000",
30333 => "010000100001000011111000",
30334 => "001111011000111010110010",
30335 => "001101011011001101101000",
30336 => "001011100011001010010100",
30337 => "001010010000100111010010",
30338 => "001010111000100001000000",
30339 => "001101010001011101000110",
30340 => "010000000110000100110110",
30341 => "010010101001111000001000",
30342 => "010011111100111011011100",
30343 => "010011011100001100011100",
30344 => "010001100101101000111010",
30345 => "001111100111111001001010",
30346 => "001110111010110111011000",
30347 => "001111011001000110111100",
30348 => "010000010100001110010100",
30349 => "010000011110001010010110",
30350 => "001110000100101010110010",
30351 => "001001110011111100110101",
30352 => "000110010011000010100011",
30353 => "000100000001001110011010",
30354 => "000001000100011100100111",
30355 => "111100000001100100100101",
30356 => "110110010011011010110010",
30357 => "110011010110001000001100",
30358 => "110011111100011101100010",
30359 => "110101001101000101111001",
30360 => "110101110101111011011001",
30361 => "110111000000011100110001",
30362 => "111001001100001010101010",
30363 => "111100111010000011101111",
30364 => "000010001111100100110011",
30365 => "000111000110011010000111",
30366 => "001000101010010000110100",
30367 => "000110000111101101010101",
30368 => "000001011011100101111001",
30369 => "111100100011110101001110",
30370 => "110111101101100101010010",
30371 => "110010100101011101110110",
30372 => "101101000001011111101000",
30373 => "100111100011011101001101",
30374 => "100011100100110000111001",
30375 => "100001110100000001101110",
30376 => "100001111100011101100101",
30377 => "100011111110010110111011",
30378 => "100111110000011111000011",
30379 => "101100011011010011011000",
30380 => "110010100111010010000010",
30381 => "111011010111101101000010",
30382 => "000100011111001111101001",
30383 => "001010110010011010111010",
30384 => "001101111011101001110000",
30385 => "001111001100110110011100",
30386 => "010000000111111101001000",
30387 => "010010010010101011110100",
30388 => "010101000110001000011100",
30389 => "010110110111011111001110",
30390 => "011000001100110101100001",
30391 => "011000101010111000111111",
30392 => "010110001111100011111100",
30393 => "010010010000111011111010",
30394 => "001110111110110010100000",
30395 => "001011100001011011110010",
30396 => "000110001000101011111100",
30397 => "111110111000001010111001",
30398 => "111000001011011110000100",
30399 => "110100101001000010111101",
30400 => "110100001001110110111011",
30401 => "110100010100000000111110",
30402 => "110100111000100110000000",
30403 => "111001011011001110001000",
30404 => "000010011001000010001000",
30405 => "001100000010101010111100",
30406 => "010100110110000001101000",
30407 => "011010101000111111011010",
30408 => "011010111010101110011100",
30409 => "011001000110011010010011",
30410 => "010110000001001111010000",
30411 => "001100111101110100111000",
30412 => "000000000000100000010100",
30413 => "110011101000110110111110",
30414 => "101000010010101101111000",
30415 => "100001110101001101110111",
30416 => "100001011101100111100000",
30417 => "100001011100101001011011",
30418 => "100000111100011011101001",
30419 => "100001011111011100000011",
30420 => "100001100000001111111001",
30421 => "100011100101100011001101",
30422 => "101010100100110011011010",
30423 => "110010100101111111100000",
30424 => "111000101110000111101100",
30425 => "111110101100110111110111",
30426 => "000100111001011111110010",
30427 => "001001001110111011100000",
30428 => "001010110000001011011100",
30429 => "001010000000001011010010",
30430 => "000111110100100011100011",
30431 => "000101001110100110000110",
30432 => "000010001011100100011011",
30433 => "111101001101100101101011",
30434 => "110110111101101111110110",
30435 => "110010100011000010100100",
30436 => "110001010010010101000010",
30437 => "110010101100011111110000",
30438 => "110110000010010110011110",
30439 => "111010011001001011111010",
30440 => "111111111010101100111010",
30441 => "000101110001000101100101",
30442 => "001001011101001111100100",
30443 => "001011001000011101010110",
30444 => "001011111001110100011110",
30445 => "001010100000010010001011",
30446 => "000110010010010001111011",
30447 => "000000111101101100100011",
30448 => "111100101101111110100110",
30449 => "111010100010011010101000",
30450 => "111010100111111111111011",
30451 => "111101010011100100010001",
30452 => "000001101000011110100011",
30453 => "000101101001111100010101",
30454 => "001000110000100111011011",
30455 => "001010101011001011110011",
30456 => "001010100001111101110010",
30457 => "001000000110000110111110",
30458 => "000011011011011011000110",
30459 => "111101010111010010000100",
30460 => "111000000100101100111010",
30461 => "110100001000001101101000",
30462 => "110000001011001100001110",
30463 => "101100100110001101101000",
30464 => "101011011001111010001000",
30465 => "101100010011101100010110",
30466 => "101100011111001011100010",
30467 => "101010111100101100101110",
30468 => "101001001100111001100010",
30469 => "101000010000010101010110",
30470 => "101000101010110001101000",
30471 => "101010100010111011000110",
30472 => "101101010100111000111000",
30473 => "110001101101000111001110",
30474 => "110111110101101101000110",
30475 => "111101110010010001101100",
30476 => "000010110110100001000010",
30477 => "000111010011001011100010",
30478 => "001010000101100110010011",
30479 => "001011001110111010011011",
30480 => "001100000000110010101110",
30481 => "001100000011010011001000",
30482 => "001010010011100111111001",
30483 => "000111001101100111011110",
30484 => "000011111101101010011100",
30485 => "000001011010000010010100",
30486 => "000000010000100000010010",
30487 => "000000111110011110100101",
30488 => "000010101110110110110101",
30489 => "000100110100001101100001",
30490 => "000111111100000010111110",
30491 => "001011001101111000111011",
30492 => "001100111000011011111010",
30493 => "001110011100001100110010",
30494 => "010001110010000111110100",
30495 => "010101101010000111001100",
30496 => "011000010101000001001111",
30497 => "011001100110101111011100",
30498 => "011010100000111000101011",
30499 => "011011100001110001111011",
30500 => "011010101011011110101111",
30501 => "010110011110010000000110",
30502 => "010000101111001010001110",
30503 => "001011101000110000010110",
30504 => "000111110110111101000001",
30505 => "000110001001110100011011",
30506 => "000110001101001110110111",
30507 => "000101101110101100000101",
30508 => "000100010100101010100111",
30509 => "000100010111110011010001",
30510 => "000101111000111101101010",
30511 => "000110111010011101001101",
30512 => "001000000111111100101110",
30513 => "001010010100101010110110",
30514 => "001100001111101011010010",
30515 => "001101000101101010001010",
30516 => "001011110010111100000111",
30517 => "000111111000101110100011",
30518 => "000011001011011110010011",
30519 => "111101110010010101000000",
30520 => "110110111001011100110011",
30521 => "110000010110001001000110",
30522 => "101010100000000101111100",
30523 => "100100110001101101010011",
30524 => "100001101111101101110001",
30525 => "100001110011110100110111",
30526 => "100001111111011001001001",
30527 => "100010000100000010001000",
30528 => "100010110000000000111001",
30529 => "100011111011100001111010",
30530 => "100111110101101100000010",
30531 => "101111110001110110001110",
30532 => "111001010101011011100010",
30533 => "000010011011111000010111",
30534 => "001001111010101100110010",
30535 => "001110001101011010110010",
30536 => "001111011110000001010010",
30537 => "001111001100100001100110",
30538 => "001110010000101000011010",
30539 => "001101011010001001101010",
30540 => "001100110111001010100100",
30541 => "001011100000010011001000",
30542 => "001000010011001011000010",
30543 => "000011101010111010100011",
30544 => "111111010010000001111100",
30545 => "111100001101001001000101",
30546 => "111001011110010111110011",
30547 => "110110000010110011111110",
30548 => "110010110100111011011010",
30549 => "110001001000101111100010",
30550 => "110001010011101010110110",
30551 => "110011001101110111100100",
30552 => "110110011110110110010110",
30553 => "111011011000101111111001",
30554 => "000011001100000101111101",
30555 => "001101001101000110100110",
30556 => "010110000001000001011110",
30557 => "011011011100101001001001",
30558 => "011101111000100111111110",
30559 => "011101100011011110011110",
30560 => "011010000101000100101111",
30561 => "010011110011100100111010",
30562 => "001011111111001100100000",
30563 => "000100110111110111011001",
30564 => "111111110100000100110111",
30565 => "111010111111000000100010",
30566 => "110100111001111101010101",
30567 => "101111011000101011011000",
30568 => "101011010101001011000000",
30569 => "100111110010011000000110",
30570 => "100101101101101111011111",
30571 => "100110010110011100010011",
30572 => "101001010011000011010110",
30573 => "101110110100001010010100",
30574 => "110110011010010011010001",
30575 => "111101011010111000010110",
30576 => "000011000000101010011100",
30577 => "001000110101111110100111",
30578 => "001111001111100000100000",
30579 => "010100101110000000010010",
30580 => "010111100011111010011100",
30581 => "010110100101011100000010",
30582 => "010010010011010010101000",
30583 => "001100011001110001111100",
30584 => "000101101100010011101101",
30585 => "111110101110011000010000",
30586 => "111000110001001110101001",
30587 => "110100100000101010101010",
30588 => "110010100100011100101110",
30589 => "110011101001110101111100",
30590 => "110110011101101000100000",
30591 => "111001110000011111111010",
30592 => "111110000010101111101101",
30593 => "000001111110111111100111",
30594 => "000011100101100001010000",
30595 => "000011101100010010010111",
30596 => "000011010010101000111011",
30597 => "000010010110000011101100",
30598 => "000001001001011010010011",
30599 => "111111101010001001100101",
30600 => "111110111100111000010011",
30601 => "000001000000101111100011",
30602 => "000100111001011111011101",
30603 => "001000000111001011100010",
30604 => "001010100011010001010010",
30605 => "001101010000100100110010",
30606 => "001111011110011111100000",
30607 => "001111100111111100011100",
30608 => "001101101111100101001100",
30609 => "001010000100010101100010",
30610 => "000100001101100000010100",
30611 => "111101101100000100111111",
30612 => "111000010000110101110001",
30613 => "110011101110101100011000",
30614 => "101111100100000110110110",
30615 => "101010100010000011001100",
30616 => "100100101110101111011111",
30617 => "100001100100111001101101",
30618 => "100001101110100001000011",
30619 => "100011010100011101101101",
30620 => "100111111001011011011010",
30621 => "110000000000001101100000",
30622 => "111000101000001001001101",
30623 => "111111111101111111000011",
30624 => "000101010101011001110100",
30625 => "001000100110011100100000",
30626 => "001010110011100111001010",
30627 => "001100001000100110111100",
30628 => "001100001101000010000000",
30629 => "001010011010001100101100",
30630 => "000101111111000100110110",
30631 => "000000011010101110101001",
30632 => "111011111001010111011110",
30633 => "111000101101111010001001",
30634 => "110110100100010000011110",
30635 => "110100111101000001000101",
30636 => "110100010000101000101111",
30637 => "110110000111101011101100",
30638 => "111001101110111101011110",
30639 => "111100100000000010110010",
30640 => "111110011011110110010000",
30641 => "000001000100001111000011",
30642 => "000100011001000110101111",
30643 => "000111010111001011001111",
30644 => "001001010110110100110001",
30645 => "001010011101001111001011",
30646 => "001010111011100010001111",
30647 => "001010101111010000001100",
30648 => "001001100010001101110000",
30649 => "000111100111001101000001",
30650 => "000101110100111010101000",
30651 => "000011101101100010111110",
30652 => "000000101000011101000111",
30653 => "111110010100100001011111",
30654 => "111110101000011000000110",
30655 => "000000111000101000001101",
30656 => "000011000011010011011100",
30657 => "000011101000000110010001",
30658 => "000010111111011100111000",
30659 => "000011001001010010111011",
30660 => "000101001011100000111101",
30661 => "001000000000001000001100",
30662 => "001010010011110100011011",
30663 => "001100000111111001001100",
30664 => "001100110010100100101000",
30665 => "001011001001111001101001",
30666 => "001001001100001100000101",
30667 => "001001010110000010101011",
30668 => "001001101110101000001100",
30669 => "000111110100001000001111",
30670 => "000100010000100100110000",
30671 => "000000011001101000010000",
30672 => "111100001000100010111000",
30673 => "110110101100011100010000",
30674 => "110000100011011001110000",
30675 => "101011001100010110111000",
30676 => "100111100011011010111111",
30677 => "100111001101111001010011",
30678 => "101011011011000011011010",
30679 => "110010011000111100010110",
30680 => "111010000101100011010100",
30681 => "000001110000000000000110",
30682 => "001000001010000100011100",
30683 => "001101010000101010010010",
30684 => "010001101001100001101010",
30685 => "010100000100111110000010",
30686 => "010011100010101111100010",
30687 => "010000010000100101000110",
30688 => "001011000100100101001111",
30689 => "000110010100011101110010",
30690 => "000010111011010101100100",
30691 => "111110101101110001110001",
30692 => "111001011011011001101010",
30693 => "110101100101101100011001",
30694 => "110011011000100010100110",
30695 => "110001010100010011001110",
30696 => "110000000110110110001000",
30697 => "110000010100110000100010",
30698 => "110000000111011110011100",
30699 => "101111000001101000001010",
30700 => "101111001001111110100100",
30701 => "110001101100000001010110",
30702 => "110110001011101101111011",
30703 => "111011010101010000010010",
30704 => "111111011111101001000100",
30705 => "000011000100011001001001",
30706 => "000111011111100001000100",
30707 => "001011110011001010000010",
30708 => "001110011111101001100100",
30709 => "001111001000010000110100",
30710 => "001100010111101110101100",
30711 => "000110110010101000100110",
30712 => "000001111010101010110110",
30713 => "111101111100101010101101",
30714 => "111000101101111011011100",
30715 => "110011101010100001011100",
30716 => "110000100000111001001110",
30717 => "101110100100101100111110",
30718 => "101101110011000100100010",
30719 => "101101101110100010100110",
30720 => "101101101101100010100010",
30721 => "101111100011000100101000",
30722 => "110100000001110110111100",
30723 => "111001010111010111100101",
30724 => "111110111011111011111000",
30725 => "000101000111010101001000",
30726 => "001011001100001111010010",
30727 => "001111111011101000110110",
30728 => "010010111011111001111010",
30729 => "010101010010111100101000",
30730 => "011000000100111011001001",
30731 => "011010100011001000011000",
30732 => "011010101010000100111101",
30733 => "010111010001011111010010",
30734 => "010001111010001001001000",
30735 => "001100000001011000011110",
30736 => "000101001010011110011010",
30737 => "111110010001110101111010",
30738 => "111001000110110010001111",
30739 => "110110000011011001110010",
30740 => "110110010010010011000100",
30741 => "111001110010100110100111",
30742 => "111110010111110010100010",
30743 => "000011101000111100110100",
30744 => "001000101001101100010101",
30745 => "001010110000101001110001",
30746 => "001010101101101000101111",
30747 => "001001111101101011010010",
30748 => "000111001100110000010100",
30749 => "000010101010001110001110",
30750 => "111110010001011101100000",
30751 => "111010101101111011111000",
30752 => "111000011100111011011110",
30753 => "110111101111101000111011",
30754 => "110111110100110010000101",
30755 => "111000100110010000101111",
30756 => "111011001100001011110001",
30757 => "111110111100000000010000",
30758 => "000001000110100110011001",
30759 => "000001010100100110001000",
30760 => "000000100000100001010010",
30761 => "111101001111011100001101",
30762 => "110111110100110110110101",
30763 => "110010000110111001111110",
30764 => "101010111001110101010000",
30765 => "100011111000001000000110",
30766 => "100010000010111101110111",
30767 => "100011110111010100100001",
30768 => "100101000000100010100101",
30769 => "100101101100110001001110",
30770 => "100110011111010000011101",
30771 => "101001000000101000001010",
30772 => "110000100110001010010100",
30773 => "111010110011011001100101",
30774 => "000010110011010010111111",
30775 => "001001000000110001000011",
30776 => "001110101111100000001000",
30777 => "010010111110111100011010",
30778 => "010100110110101110010110",
30779 => "010100011100010011101110",
30780 => "010010111001110001011010",
30781 => "010000010011000000010000",
30782 => "001011101011011101010001",
30783 => "000110101100111101011100",
30784 => "000010111101101011110110",
30785 => "111111111111001100001010",
30786 => "111110010111111011001011",
30787 => "111110000100010010011010",
30788 => "111110001000100100010101",
30789 => "111111011001001110011000",
30790 => "000001001100010000011111",
30791 => "000010000100100001000101",
30792 => "000011011100010100100100",
30793 => "000101110101000000111011",
30794 => "000111110101010011001000",
30795 => "001001001110010100111000",
30796 => "001010000000001111100110",
30797 => "001010001110111111110110",
30798 => "001010010101000110110101",
30799 => "001001101010111011011111",
30800 => "000111101010011001100000",
30801 => "000101011100011011110100",
30802 => "000100111111011101010000",
30803 => "000110000110000000011001",
30804 => "000110101000010100100110",
30805 => "000110101100110010000110",
30806 => "000110100100101001011100",
30807 => "000100010010011011010111",
30808 => "000000101100001010111011",
30809 => "111110000011100010000110",
30810 => "111011101110100100101001",
30811 => "111010001001001011001001",
30812 => "111010011111001100011010",
30813 => "111011000001110000000101",
30814 => "111010111111100001001100",
30815 => "111100000000011110010011",
30816 => "111110011001001000101101",
30817 => "000000111111110001011111",
30818 => "000011010101101001100111",
30819 => "000101110101000100011000",
30820 => "000111110111011001111010",
30821 => "000111111000111111000101",
30822 => "000101100101101011101001",
30823 => "000001100110010111010110",
30824 => "111100110100000101001001",
30825 => "111000010000111101010100",
30826 => "110100011001001100100000",
30827 => "110010000101010011001100",
30828 => "110010011110001010110000",
30829 => "110101100000110101001001",
30830 => "111010101111011111010110",
30831 => "000001000000100000010010",
30832 => "000111000000111110011100",
30833 => "001100110111001101001110",
30834 => "010010010000100101011000",
30835 => "010110101000101100100100",
30836 => "011001101010010100001111",
30837 => "011001101010110000111100",
30838 => "010111000010011010001010",
30839 => "010100001010000010000010",
30840 => "010000000011110101110000",
30841 => "001010011011010100011111",
30842 => "000110110011001111101100",
30843 => "000110000001000110101001",
30844 => "000110000000000010000110",
30845 => "000110011111011000111101",
30846 => "000110111110000111011011",
30847 => "000101011001101001011110",
30848 => "000010000011111001101100",
30849 => "111110111001101011011000",
30850 => "111011100111110010101000",
30851 => "111000010111101000010110",
30852 => "110111010110000110011011",
30853 => "110111100101011001010110",
30854 => "110111000000011101010010",
30855 => "110111001010000011000000",
30856 => "111000110100111010110011",
30857 => "111011011010011011000100",
30858 => "111111000110001110110101",
30859 => "000001011110001100000010",
30860 => "000000010010100000010010",
30861 => "111101010100011000111011",
30862 => "111001111011001001011000",
30863 => "110110010001101101111000",
30864 => "110010110111110110111010",
30865 => "101110110100000110101000",
30866 => "101001110101100001000000",
30867 => "100101111101000101010111",
30868 => "100100100001111110010111",
30869 => "100101000111001100010101",
30870 => "100110110010101100101000",
30871 => "101001010101010011101100",
30872 => "101101001101001110110010",
30873 => "110010110010101010110100",
30874 => "111001001111011010010001",
30875 => "111110100000011110010000",
30876 => "000010010010110101110101",
30877 => "000101111011100011011001",
30878 => "001000011101011110111101",
30879 => "001001000110010110001011",
30880 => "001010011101111011011100",
30881 => "001110000110110100111000",
30882 => "010001101110111100010110",
30883 => "010010001010101010101000",
30884 => "001111001011000111001000",
30885 => "001100000100101100001100",
30886 => "001010001110010011011010",
30887 => "000111010100001001100010",
30888 => "000011001111111010100011",
30889 => "000000011101010100111010",
30890 => "111111110110010100110101",
30891 => "000001001010101110000001",
30892 => "000011110010011010001110",
30893 => "000110010111101110000100",
30894 => "001000010001011110101100",
30895 => "001010001101101001101111",
30896 => "001100001111000000000010",
30897 => "001101000101001000001010",
30898 => "001100110110001011011100",
30899 => "001100001101011000101110",
30900 => "001001100111100011000011",
30901 => "000100101010010000101000",
30902 => "111111111100001001100010",
30903 => "111100101011011000000001",
30904 => "111010011110101101000101",
30905 => "111001101010101110000001",
30906 => "111001111101010000100010",
30907 => "111010101010101011010110",
30908 => "111011111101101011101011",
30909 => "111101101111000001111011",
30910 => "111111101100010100100100",
30911 => "000001100000001001001110",
30912 => "000001010000000101110000",
30913 => "111110000001101110011001",
30914 => "111001110010000110010101",
30915 => "110011101100101101010010",
30916 => "101010000100101110010000",
30917 => "100010100011100110000011",
30918 => "100001011110100000000111",
30919 => "100001111101111111101101",
30920 => "100001110011100110110100",
30921 => "100011000110110100100101",
30922 => "100100001111010010011011",
30923 => "100101111000100111010110",
30924 => "101011100000110110110100",
30925 => "110011010110011010010110",
30926 => "111011000001010100001001",
30927 => "000010111000000011000101",
30928 => "001001110100000011010110",
30929 => "001110110100010110110000",
30930 => "010001110010011010010110",
30931 => "010010001010000011100010",
30932 => "010000011110110100011110",
30933 => "001101100010011001111100",
30934 => "001001101010110000001010",
30935 => "000110011100111010011110",
30936 => "000100110000011011111100",
30937 => "000010111110000000001101",
30938 => "111111110001101001000000",
30939 => "111100001001111111000000",
30940 => "111001110000101111111011",
30941 => "111001100001011100000010",
30942 => "111011100000011111011110",
30943 => "111110011111101100000100",
30944 => "000001111001110101100010",
30945 => "000110110100010100000000",
30946 => "001011110011101010011000",
30947 => "001101111010000110001010",
30948 => "001101111000101011101110",
30949 => "001100111111100100011100",
30950 => "001010010110101001000011",
30951 => "000111001101110010110001",
30952 => "000101111000111110101001",
30953 => "000110010000001000110111",
30954 => "000111001101010001000100",
30955 => "000111110110000101101110",
30956 => "000111100000011111110000",
30957 => "000110001001110110101011",
30958 => "000011111000100000011010",
30959 => "000001011011101101011001",
30960 => "111111111011100001000110",
30961 => "111110101001110101010001",
30962 => "111011111100101101010011",
30963 => "111000100110011001011000",
30964 => "110110111110010111010011",
30965 => "110111100110111111110101",
30966 => "111001000110100010101000",
30967 => "111010001010100011110010",
30968 => "111011001000101010110110",
30969 => "111101010111101001001010",
30970 => "000000010000101011010111",
30971 => "000001101011010111101111",
30972 => "000001001110101010010001",
30973 => "111111010001110111010110",
30974 => "111100001010100110011100",
30975 => "111001100011000011110100",
30976 => "111000000101101111111110",
30977 => "110110110001000010001101",
30978 => "110101010110101101110000",
30979 => "110011100101100001001110",
30980 => "110001000101000110011110",
30981 => "101111010100011100110110",
30982 => "101111101000101100111000",
30983 => "110001000100110001000010",
30984 => "110011001010000000011000",
30985 => "110111011011111010000011",
30986 => "111101011111001010100001",
30987 => "000010010011010101011110",
30988 => "000101011011010001000011",
30989 => "000111100100110101110000",
30990 => "000111100110010001100110",
30991 => "000110011101100000100000",
30992 => "000101101111010011110110",
30993 => "000100001011101011010001",
30994 => "000010111001010100100001",
30995 => "000100001011111110010010",
30996 => "000101111111011010110001",
30997 => "000110101001010100110100",
30998 => "000111101000010100011100",
30999 => "001001000101101100101110",
31000 => "001010010101110000100111",
31001 => "001100000000001111110000",
31002 => "001101101011011100100010",
31003 => "001101011010101100111010",
31004 => "001010110110101011100101",
31005 => "000111000001100000011100",
31006 => "000010010101000011100010",
31007 => "111110011101010000001011",
31008 => "111101001110010001000010",
31009 => "111101100000011101001100",
31010 => "111111000111111110001101",
31011 => "000010110010111010011100",
31012 => "000110001110101011001001",
31013 => "001000100010000001001110",
31014 => "001010110001110000000110",
31015 => "001011100110110110101010",
31016 => "001010100001000001101111",
31017 => "001000010010100001011100",
31018 => "000100011110011000000100",
31019 => "000000101100000011111100",
31020 => "111110111111001111101010",
31021 => "111110010011000111111101",
31022 => "111101111101101111010111",
31023 => "111110100100100011001111",
31024 => "111111101110101101011010",
31025 => "000001001000011110111111",
31026 => "000010011101010100000111",
31027 => "000010000101100111011111",
31028 => "111110110011010111010010",
31029 => "111010001100010010110100",
31030 => "110110111011110100011101",
31031 => "110101101010010000110000",
31032 => "110110001001111011111010",
31033 => "111000101111111010111000",
31034 => "111101000110011100110110",
31035 => "000010010111001111001010",
31036 => "000111100000011110100110",
31037 => "001011111111001001010100",
31038 => "010000011110011101010110",
31039 => "010100001110101110111000",
31040 => "010101000011010001000100",
31041 => "010010111110111100111100",
31042 => "001111101010111000011110",
31043 => "001100010110111000000100",
31044 => "001001111000111001111000",
31045 => "000111101110011010100110",
31046 => "000100100011010001101000",
31047 => "000000111010110110101101",
31048 => "111111000011101010010111",
31049 => "111111011001101111011110",
31050 => "111111100111011000000000",
31051 => "111110010110010111001100",
31052 => "111100101100010000111100",
31053 => "111011101101010110011111",
31054 => "111100000000101101001011",
31055 => "111101110010111110111110",
31056 => "000000001100001100101011",
31057 => "000010011110000110001000",
31058 => "000101000110000100011100",
31059 => "001000101100100010000111",
31060 => "001100011000101010110110",
31061 => "001110100010010000111000",
31062 => "001110110100001011010000",
31063 => "001100110000110001101100",
31064 => "000111010111101000101001",
31065 => "111110011101011000110100",
31066 => "110010010000101011001000",
31067 => "100110101011101110001110",
31068 => "100001101101101111011101",
31069 => "100001101100000001111011",
31070 => "100001011101000010001101",
31071 => "100001010111111101110011",
31072 => "100010000100100011110010",
31073 => "100011001100111110000001",
31074 => "100111000001010011100110",
31075 => "101110001001101010101110",
31076 => "110111011000110101011100",
31077 => "000001110110011101111001",
31078 => "001011010011110011001000",
31079 => "010010011001101111111100",
31080 => "010111011000110011010010",
31081 => "011001011100001000000001",
31082 => "010111110110000001101010",
31083 => "010011011100110000100110",
31084 => "001110000001000101110000",
31085 => "001000100100110010001010",
31086 => "000010101010110010110010",
31087 => "111100110100000010000101",
31088 => "110111101111010110000100",
31089 => "110010000000001000000110",
31090 => "101011000011101001011010",
31091 => "100101001100001001100100",
31092 => "100011100000000101110111",
31093 => "100111011111001100101010",
31094 => "101111000010010000110110",
31095 => "110111001110111110000100",
31096 => "111111110000000010011111",
31097 => "001000001101110111010100",
31098 => "001110011111010111010000",
31099 => "010000111011011011111010",
31100 => "010000000000001000011110",
31101 => "001101000111110010100000",
31102 => "001000111110100100010011",
31103 => "000100111100011010011000",
31104 => "000010101111000100000001",
31105 => "000001100100100001100001",
31106 => "000000010111110000100100",
31107 => "111111011000111010111100",
31108 => "111110010001011010101011",
31109 => "111101100111011000100011",
31110 => "111110101110110101011010",
31111 => "000000101111010111111110",
31112 => "000010001011111010001100",
31113 => "000010011010001110101101",
31114 => "000000111011000011111101",
31115 => "111110011111001001010100",
31116 => "111100110110001101011110",
31117 => "111100110011100010110101",
31118 => "111101100101101000011011",
31119 => "111110010010010100011000",
31120 => "111111001011101001011110",
31121 => "000000011010100000001101",
31122 => "000001101000000101000001",
31123 => "000010110001001111100000",
31124 => "000011000011011111110111",
31125 => "000010001001110101010001",
31126 => "000001011111010001000000",
31127 => "000001101011011011101110",
31128 => "000010000101100100111010",
31129 => "000010000001010100110111",
31130 => "000000100000000100110000",
31131 => "111101001011101110111101",
31132 => "111000101111011000000101",
31133 => "110100001111111100111110",
31134 => "110000101001101010110010",
31135 => "101101101110101001010100",
31136 => "101011101010100100101000",
31137 => "101011111010110101101000",
31138 => "101110001101100010010010",
31139 => "110000111011110110000110",
31140 => "110011100000101001111110",
31141 => "110101010001111010010011",
31142 => "110110001100101001100000",
31143 => "110111111000110011000010",
31144 => "111010011010001100000100",
31145 => "111011100110010001010010",
31146 => "111011010000001010001010",
31147 => "111011100101000100011101",
31148 => "111101001000100101001011",
31149 => "111110101111010000101010",
31150 => "000000011101011110110001",
31151 => "000010011011101001101011",
31152 => "000011101111000100101101",
31153 => "000100101111010000100100",
31154 => "000101010100001100101101",
31155 => "000010101110111111000001",
31156 => "111101000110000001111001",
31157 => "111000011110010101000110",
31158 => "110101101000110101000100",
31159 => "110010100001101010010110",
31160 => "101111110100110000010010",
31161 => "101110111000111101100110",
31162 => "110000101101010100011000",
31163 => "110110111000110011101101",
31164 => "111111001000001110010101",
31165 => "000101100100000001011010",
31166 => "001011100000001010011011",
31167 => "010010000111110001001110",
31168 => "010110100011011010000100",
31169 => "010111001110010110111110",
31170 => "010100100011110101001000",
31171 => "010000100110010101101010",
31172 => "001110111110101011000010",
31173 => "001111001001100110100100",
31174 => "001101000100111100100110",
31175 => "001001011000010100000110",
31176 => "001000001010011010110100",
31177 => "001001100101011100101011",
31178 => "001010010011101010110001",
31179 => "001001010001001010001101",
31180 => "000111110110110011011101",
31181 => "000111001101000100100111",
31182 => "001000010101010100101101",
31183 => "001010000111111001111100",
31184 => "001001111111111010111101",
31185 => "001001101101011011000000",
31186 => "001011110101111001001011",
31187 => "001110101010000001111100",
31188 => "010001001110111110000010",
31189 => "010100010110111101100110",
31190 => "010111000110010000110010",
31191 => "011000010101000110010001",
31192 => "010110111011010011110000",
31193 => "010010001101000101101010",
31194 => "001011011011001011011101",
31195 => "000011110000010100000100",
31196 => "111100000011011101001101",
31197 => "110101010011000111010100",
31198 => "101111101010010000001100",
31199 => "101100000011000001000100",
31200 => "101011010110101000001100",
31201 => "101100100001110110111000",
31202 => "101110000001100010011010",
31203 => "101111000111001000100010",
31204 => "110001000110011111101010",
31205 => "110101101010111111111010",
31206 => "111011001101110101100011",
31207 => "111111011100001001011011",
31208 => "000010000001100111100010",
31209 => "000011010100111110010000",
31210 => "000100010011101110101110",
31211 => "000101010100001101111100",
31212 => "000110000000111100010111",
31213 => "000110001101101101100000",
31214 => "000100000111011111010011",
31215 => "111110111010000110100000",
31216 => "110111100011001111001100",
31217 => "101101101010010000101100",
31218 => "100100100100001011000110",
31219 => "100001110111111110110111",
31220 => "100011010011101000000011",
31221 => "100100001001010010110011",
31222 => "100100101110001000010101",
31223 => "100110000000110101110011",
31224 => "101001100110110111011110",
31225 => "110001010010101100111000",
31226 => "111011000100010001011001",
31227 => "000100101011001111100000",
31228 => "001101100101011101101010",
31229 => "010100101001100110010100",
31230 => "011001100001011101111011",
31231 => "011100000001100111111001",
31232 => "011011001000011000000101",
31233 => "010111111111011111100100",
31234 => "010100101110100100010000",
31235 => "010001011000000011101000",
31236 => "001110000011100001010010",
31237 => "001011101110110101011101",
31238 => "001001111001110000011111",
31239 => "000111100100011110001100",
31240 => "000100101011101011001101",
31241 => "000000110100111101000111",
31242 => "111100000000110110110100",
31243 => "111000010000000110110001",
31244 => "110111011101001011100000",
31245 => "111001111000110010010011",
31246 => "111111001100100101001101",
31247 => "000101111101010011010110",
31248 => "001011001110001101111100",
31249 => "001101101110000111111010",
31250 => "001111010101111000110110",
31251 => "010000100001001101001110",
31252 => "001111000100000000111010",
31253 => "001011100000011010011010",
31254 => "001000100010100101010011",
31255 => "000110101101110110010010",
31256 => "000101011000111011101111",
31257 => "000011010011000101011010",
31258 => "111111101111001111101111",
31259 => "111100111010101011001001",
31260 => "111100000011100001110100",
31261 => "111100001111011110011100",
31262 => "111101111111000001011101",
31263 => "000000011111011111101100",
31264 => "000001110011000000101011",
31265 => "000010101001100010011011",
31266 => "000010111100010000010110",
31267 => "000001010001111111100011",
31268 => "111111011100100110011001",
31269 => "111111010000001010000010",
31270 => "111111100101101000001100",
31271 => "111111111001000000110000",
31272 => "000000110011101000000111",
31273 => "000001100111110011011011",
31274 => "000001100011010001110011",
31275 => "000001101111100000000110",
31276 => "000010011010111010101111",
31277 => "000011010011010001010000",
31278 => "000110110110111110000110",
31279 => "001100100111010001011100",
31280 => "001111101000100111101100",
31281 => "001111011010001010111100",
31282 => "001101101010110101100000",
31283 => "001000110000000010001000",
31284 => "000000001001100011011001",
31285 => "110100110111010001100011",
31286 => "101000110111101101001100",
31287 => "100001101100010100100001",
31288 => "100001001001010000111111",
31289 => "100001110111101001110111",
31290 => "100001010100101010010010",
31291 => "100010101000100001001000",
31292 => "100111101001001001011011",
31293 => "101110111001011010111000",
31294 => "110110101011111000000000",
31295 => "111101111011010001100110",
31296 => "000011100010110111100001",
31297 => "000111000011110000101010",
31298 => "000111101100010100010011",
31299 => "000101010100001100011001",
31300 => "000011011110010011111011",
31301 => "000011111001100100101010",
31302 => "000011000000111011110100",
31303 => "000000011001100110001001",
31304 => "111110011111000110011101",
31305 => "111011101011001011101100",
31306 => "110110110011001110110011",
31307 => "110000111010101101001110",
31308 => "101001111000000100011100",
31309 => "100011111001100011111010",
31310 => "100010010000010111010100",
31311 => "100011001111011110101010",
31312 => "100100000010111111011001",
31313 => "100101001110001111101111",
31314 => "101000010111110010100110",
31315 => "101111000100111101010100",
31316 => "111001011100011001111011",
31317 => "000011111001010011010000",
31318 => "001011011001011111000010",
31319 => "010000111001100001111000",
31320 => "010100100110010111100010",
31321 => "010100101100101100100110",
31322 => "010001110001110011000100",
31323 => "001101100011111010100110",
31324 => "001000100111011000000110",
31325 => "000100010010110010101001",
31326 => "000001110000110101000011",
31327 => "000000010010011000001110",
31328 => "111111010000000010100001",
31329 => "111111001100001010110101",
31330 => "000000100011001110011001",
31331 => "000010100101111000100001",
31332 => "000011111111010110110010",
31333 => "000100100100001111110010",
31334 => "000101101010101110110110",
31335 => "001000110001100000110100",
31336 => "001100111010100101011010",
31337 => "001111100100010001000110",
31338 => "010001111100011110101010",
31339 => "010110101010101100110110",
31340 => "011011001100010100011100",
31341 => "011100010000101001001010",
31342 => "011011001111100000110111",
31343 => "011010011011011111011011",
31344 => "011001101100100001100111",
31345 => "010110100111000111110110",
31346 => "001111111000111001101010",
31347 => "001000100010000110111001",
31348 => "000011000111111111001010",
31349 => "111111010001100011000110",
31350 => "111101111000011110011100",
31351 => "111111001000100000010010",
31352 => "000000000001100111011111",
31353 => "000000001001010101010110",
31354 => "000001101001100110010000",
31355 => "000010111111110100100001",
31356 => "000001111011011011000011",
31357 => "000000011101100100111011",
31358 => "111111111011001010011111",
31359 => "111110001100110110000011",
31360 => "111010110001100111110010",
31361 => "110111100101000001110010",
31362 => "110101111110000001100001",
31363 => "110101010011000011100000",
31364 => "110011011010001001011000",
31365 => "110000100111010110100000",
31366 => "101110001111100100110100",
31367 => "101001110101100101010000",
31368 => "100100001000001010110011",
31369 => "100010011100110001001000",
31370 => "100011011111100110000000",
31371 => "100011100111100101011100",
31372 => "100100100100111001111011",
31373 => "100101110010111111101111",
31374 => "100110001010010011000110",
31375 => "101001101011010011101110",
31376 => "110000011111111001111100",
31377 => "110110100100101010010000",
31378 => "111011111111101101101001",
31379 => "000001101000001100001001",
31380 => "000110010011110010110011",
31381 => "001001101011000001010101",
31382 => "001010110001011010001111",
31383 => "001001000111000110111110",
31384 => "000111000010110101110110",
31385 => "000101111100101010100110",
31386 => "000100101111111000111001",
31387 => "000011101001110010101110",
31388 => "000100000111001001101100",
31389 => "000110000011000000100010",
31390 => "001000000001100000110110",
31391 => "001000111100101000011011",
31392 => "001000110001101000010010",
31393 => "000111111011011001111011",
31394 => "000110110100010110000000",
31395 => "000110101000010011000010",
31396 => "001000100001011100011100",
31397 => "001011010010011110111001",
31398 => "001100111101101111000000",
31399 => "001110000110011001010110",
31400 => "001111101101101000101010",
31401 => "010000001011000011111110",
31402 => "001101111011001101001110",
31403 => "001010110001110010100010",
31404 => "001001000110110101000000",
31405 => "001000011001000001000010",
31406 => "000111001110001100110001",
31407 => "000110000001101101110101",
31408 => "000101101111101010111010",
31409 => "000101100110100000100000",
31410 => "000100000000000111100010",
31411 => "000001101010100101111000",
31412 => "000001011010101000111111",
31413 => "000011110110110011010110",
31414 => "000110101001011010101111",
31415 => "001000001001111101010100",
31416 => "001000010110011110100010",
31417 => "000111001111101010100011",
31418 => "000101000001010100001100",
31419 => "000010100101000010100001",
31420 => "000000010011000100011010",
31421 => "111101100011001011110011",
31422 => "111010100110001001010100",
31423 => "111000101011010100000110",
31424 => "110111111100110010100111",
31425 => "110111011101100111110100",
31426 => "110110000101000000100010",
31427 => "110011111101001110110110",
31428 => "110011101010011001000100",
31429 => "110111001000011110101100",
31430 => "111101100001011101101010",
31431 => "000100110101011110000101",
31432 => "001010101110111001110110",
31433 => "001101110011100011101100",
31434 => "001101101000100001011010",
31435 => "001001010000111010001110",
31436 => "000001100111011110010110",
31437 => "111000111001000001001100",
31438 => "101111001001100101010100",
31439 => "100110000100001011100101",
31440 => "100001011100110111111001",
31441 => "100001011000001110100111",
31442 => "100010111100000110011101",
31443 => "100100010011010110110100",
31444 => "100110111000110010110000",
31445 => "101110001000110100100010",
31446 => "111001000100101000111110",
31447 => "000010111101000111011011",
31448 => "001001111110110001100000",
31449 => "001101111011000111111010",
31450 => "001110010001000101001010",
31451 => "001011110101111100010110",
31452 => "000111101011000111001000",
31453 => "000011001011011100000000",
31454 => "000000001010111110101101",
31455 => "111110101010000010101111",
31456 => "111101101000101110111010",
31457 => "111100001010000011011101",
31458 => "111001110100011111001000",
31459 => "110111101010001111001001",
31460 => "110110010110001010111010",
31461 => "110101010001011000011011",
31462 => "110011101111001010011000",
31463 => "110001111011000011001010",
31464 => "110001010111001110010000",
31465 => "110010100000011010011110",
31466 => "110100011001101011011001",
31467 => "110111011100111011001110",
31468 => "111011011010100110010010",
31469 => "111111100001100101111110",
31470 => "000101000000010001011000",
31471 => "001010110001100010011111",
31472 => "001101111001101101101110",
31473 => "001111000101000101001110",
31474 => "001111011010000110000110",
31475 => "001110010101000001111010",
31476 => "001100011101010011101110",
31477 => "001001111011001101010100",
31478 => "000110010110000100001011",
31479 => "000011000011111111100111",
31480 => "000001001001000110000100",
31481 => "000000010111000000001000",
31482 => "000000101100100000001001",
31483 => "000010000001100001001000",
31484 => "000011010001010011011000",
31485 => "000011011001001110101100",
31486 => "000010110001011000110011",
31487 => "000010010101010011100100",
31488 => "000010101110001110111001",
31489 => "000100100010010101100100",
31490 => "000110110001101110101111",
31491 => "001000001011100101100110",
31492 => "001010100001011010000101",
31493 => "001110110111010100101000",
31494 => "010010011110101100001000",
31495 => "010011101001001000101100",
31496 => "010011010110010100100000",
31497 => "010010001100111011111010",
31498 => "010000010010101010101000",
31499 => "001110001000011110110100",
31500 => "001011110101011100101011",
31501 => "001001000111011111000010",
31502 => "000110101010010010110100",
31503 => "000101100111110101011000",
31504 => "000101011101010100111001",
31505 => "000100110001100011000110",
31506 => "000011110100011111111010",
31507 => "000011101001010110101110",
31508 => "000100000111110111111111",
31509 => "000100000100000001111100",
31510 => "000010100000011011010100",
31511 => "111111101001011101101001",
31512 => "111100011011000001111101",
31513 => "111001110001110010000110",
31514 => "111000101100001001110101",
31515 => "111001101111000110100100",
31516 => "111100001001001001010111",
31517 => "111110001010110100011001",
31518 => "111111000010100111010110",
31519 => "111110100110001001101001",
31520 => "111011001100001011111000",
31521 => "110100101001011101101000",
31522 => "101110111110011101110000",
31523 => "101100100010100010010110",
31524 => "101011001101010110000000",
31525 => "101001111101101011111010",
31526 => "101001110010000010000100",
31527 => "101010001011101000011100",
31528 => "101010001110100101101110",
31529 => "101010100001000011111110",
31530 => "101100101001100011001000",
31531 => "110000101110010111000100",
31532 => "110011110011101011100110",
31533 => "110100010100010001000110",
31534 => "110100110011010100001010",
31535 => "110110011010111110111001",
31536 => "110111011000101111000000",
31537 => "111000001001110001110011",
31538 => "111010100111010110110101",
31539 => "111110000110000100010110",
31540 => "000001001010111110000100",
31541 => "000100001111111010000000",
31542 => "000111111010101000010111",
31543 => "001010111011111111100100",
31544 => "001011101011111010110110",
31545 => "001010101100011000100100",
31546 => "001001100000000010101100",
31547 => "001000101011011000110100",
31548 => "001000100110100000000111",
31549 => "001000101111110100110110",
31550 => "000110111011100110101001",
31551 => "000010111000001101010000",
31552 => "111111011011001110001101",
31553 => "111110010010000111111110",
31554 => "111101111101001100000010",
31555 => "111100101111111100110101",
31556 => "111100001011110000100000",
31557 => "111111001011011100011100",
31558 => "000100111111000110011010",
31559 => "001010001000000101001000",
31560 => "001101110000110110010110",
31561 => "010001000100101101101100",
31562 => "010011010010110110011100",
31563 => "010011010011010011010000",
31564 => "010010101100100100010000",
31565 => "010011010010010010101000",
31566 => "010011111001111011010000",
31567 => "010010100110000111100010",
31568 => "001111100000111010101010",
31569 => "001100001010110001111110",
31570 => "001001011011101001011000",
31571 => "000111000001111100011000",
31572 => "000100100001010111110110",
31573 => "000001101011001000110011",
31574 => "111110011001101110100110",
31575 => "111011100001000100101110",
31576 => "111001101000010010001000",
31577 => "110111110111101000011010",
31578 => "110101101110100111011000",
31579 => "110011111001100111000110",
31580 => "110011111000111110111010",
31581 => "110111100010000000011000",
31582 => "111110010111010111100111",
31583 => "000110001110010001100001",
31584 => "001101110100001100111010",
31585 => "010011011001110100100010",
31586 => "010101011011000101000110",
31587 => "010011100010010111001100",
31588 => "001101011001111000000000",
31589 => "000100011010011001100000",
31590 => "111001010110001010000011",
31591 => "101011110011110011011010",
31592 => "100010000001111101111010",
31593 => "100000111110110101010011",
31594 => "100001111110110010101111",
31595 => "100001011011101000111101",
31596 => "100010101111100011010111",
31597 => "100011111101111110100101",
31598 => "100101011110011101111110",
31599 => "101100110010000001100110",
31600 => "110111001000011101001100",
31601 => "111110101010010100100101",
31602 => "000011100010000000011100",
31603 => "000110010011111111110001",
31604 => "000110110000000111011000",
31605 => "000101011101101100110110",
31606 => "000010111010111101100001",
31607 => "000000101100000110110101",
31608 => "111111001000001110000110",
31609 => "111100101011111001011100",
31610 => "111010010111101000111100",
31611 => "111001011100000010101001",
31612 => "111000000010100001000010",
31613 => "110101110011000100110011",
31614 => "110101000110110111000010",
31615 => "110110010011100011101111",
31616 => "110111100110101110010001",
31617 => "111000110100011110110101",
31618 => "111010100000101000001001",
31619 => "111100001111011100011010",
31620 => "111110001011100000100001",
31621 => "000000000000100101010100",
31622 => "000000100100001111100110",
31623 => "000001011000000001011011",
31624 => "000011110010110000001011",
31625 => "000101111000111101010101",
31626 => "000111100101111011011100",
31627 => "001010001011110010011010",
31628 => "001100001111110110100010",
31629 => "001101000111011011100100",
31630 => "001101010100010101000100",
31631 => "001100010001101110101110",
31632 => "001010110101101011000001",
31633 => "001001111100000001110001",
31634 => "001000001001010111101110",
31635 => "000101010110111011101100",
31636 => "000010111110000111001111",
31637 => "000000100100001001001101",
31638 => "111101110000100100110100",
31639 => "111011110000110111111000",
31640 => "111010100110000010011011",
31641 => "111001000100101110001000",
31642 => "110111110110110111010000",
31643 => "111000010101110101101000",
31644 => "111010000111110011001011",
31645 => "111100101100110001111010",
31646 => "000000010011001110011110",
31647 => "000100010000011011010000",
31648 => "000111111100001100000110",
31649 => "001011000010001001110100",
31650 => "001100011110111011100010",
31651 => "001100001000010001011010",
31652 => "001010101011000010011101",
31653 => "001000000111101011000011",
31654 => "000101000011000100001101",
31655 => "000010100110100100111111",
31656 => "000001001111111010011001",
31657 => "000001001000010001110110",
31658 => "000001100111101100010001",
31659 => "000001111000110010101001",
31660 => "000010001100101110111001",
31661 => "000010011000110110010101",
31662 => "000001100101001010011011",
31663 => "111111111000010000110110",
31664 => "111101101100110001110011",
31665 => "111011000010111011111001",
31666 => "111000011100011111001000",
31667 => "110110101111100010001100",
31668 => "110110000000101010010000",
31669 => "110110000110101110100010",
31670 => "110111001010110000101010",
31671 => "111000000110100000100101",
31672 => "110111101101011010010101",
31673 => "110111001010001101010000",
31674 => "110111101010001001000111",
31675 => "111001010111101110110010",
31676 => "111100101000111101010011",
31677 => "111111111010111000100001",
31678 => "000001100000000111110011",
31679 => "000010011110010010101100",
31680 => "000010110010001101110100",
31681 => "000001011010101011000110",
31682 => "111111110100100111101111",
31683 => "111110110110011010001010",
31684 => "111110100111110101011101",
31685 => "000000100000001100101101",
31686 => "000011101111010001010101",
31687 => "000110010100001010010100",
31688 => "001000000111100101111011",
31689 => "001001010011101100001000",
31690 => "001010110000101001110011",
31691 => "001101111010011001000110",
31692 => "010001101110110011111110",
31693 => "010100011100010111011100",
31694 => "010101010001101111111110",
31695 => "010011100101011011100110",
31696 => "010000001011000110100100",
31697 => "001100101111101100110100",
31698 => "001010000111100100000011",
31699 => "001000011000010011000001",
31700 => "000110010010001010110110",
31701 => "000010111110010100000010",
31702 => "111111110001110100001010",
31703 => "111101001011110110010000",
31704 => "111010001011000010101110",
31705 => "110111000111011010001100",
31706 => "110101101111110010001101",
31707 => "110110101100101001111110",
31708 => "111000111010110111001100",
31709 => "111100100111100001101100",
31710 => "000011010110101110101010",
31711 => "001011110111110000110000",
31712 => "010010111001000000100000",
31713 => "010110101001001000100010",
31714 => "010111000011110001010000",
31715 => "010101101110010011100010",
31716 => "010100010010010101000110",
31717 => "010010101000010001011100",
31718 => "010000001011001001101100",
31719 => "001100000110001011101010",
31720 => "000110001010110100000010",
31721 => "000000101011011110100101",
31722 => "111101000101010000110011",
31723 => "111001110100110111001010",
31724 => "110110000111111001110110",
31725 => "110010111101001011000000",
31726 => "110001001011101000001000",
31727 => "110001000010011111001000",
31728 => "110010000111100100000010",
31729 => "110100000010111111011010",
31730 => "110110000011010000010000",
31731 => "110111100100000111101101",
31732 => "111010110100001010110010",
31733 => "000001001101101010001011",
31734 => "001000111111100100111111",
31735 => "010001011110000101000000",
31736 => "011000010010111011111100",
31737 => "011001110000001010100101",
31738 => "011000100011011001000000",
31739 => "010110101010101011011110",
31740 => "001111111001110001111000",
31741 => "000100111100110101110001",
31742 => "111001010001111010100110",
31743 => "101100011101011100111100",
31744 => "100010100100000100010011",
31745 => "100000110000101011111110",
31746 => "100010001111100101111111",
31747 => "100001110001101011100010",
31748 => "100001110010000111011111",
31749 => "100010101110110010010111",
31750 => "100010110101011111000110",
31751 => "100110100000111110011000",
31752 => "110001000011001110111000",
31753 => "111100110101000111110011",
31754 => "000101001111010101101110",
31755 => "001011100101000010111010",
31756 => "010000001000100000100100",
31757 => "010010000100110011111000",
31758 => "010001010000001100010100",
31759 => "001100100001100111000100",
31760 => "000101001001001000000010",
31761 => "111110011101111011000101",
31762 => "111000100000011011101010",
31763 => "110010100011000000101100",
31764 => "101101111110110010110010",
31765 => "101010101111010101011010",
31766 => "101000010001000011011000",
31767 => "100111111001001110100001",
31768 => "101001110010001000111010",
31769 => "101100010010010111011010",
31770 => "101111000100101011100000",
31771 => "110010011100100010111110",
31772 => "110101010100101001110001",
31773 => "110111011100111110100000",
31774 => "111010001000011111110000",
31775 => "111101010110110100011100",
31776 => "000000110000011001101011",
31777 => "000100101101010011110110",
31778 => "001000010010011101101100",
31779 => "001011010101110000011001",
31780 => "001111010100101001111100",
31781 => "010010111111000111011100",
31782 => "010100000011000110001100",
31783 => "010011001101110011010110",
31784 => "010001010011101110000110",
31785 => "001110000110001110010100",
31786 => "001010110101110110110111",
31787 => "001000011010100010101010",
31788 => "000101100110111111101101",
31789 => "000010000100111001101111",
31790 => "111110110001100111000000",
31791 => "111011110011001001111100",
31792 => "111001000001111001100000",
31793 => "110110011010010111011110",
31794 => "110011100001100100001100",
31795 => "110001110011011011100010",
31796 => "110011010001010111100000",
31797 => "110110010101100001000110",
31798 => "111000111011010110000010",
31799 => "111100100010000101110111",
31800 => "000010001101100010100101",
31801 => "001000010100100001011000",
31802 => "001100111100110110101000",
31803 => "001110110011000001001010",
31804 => "001110100111111101000010",
31805 => "001110011010011011100010",
31806 => "001101010010101110101100",
31807 => "001001110111000001101101",
31808 => "000101011010011111101000",
31809 => "000001001001110001110100",
31810 => "111101100011000111010001",
31811 => "111010110001110101011111",
31812 => "110111110100110011011010",
31813 => "110101000111110010110000",
31814 => "110100100010100111000100",
31815 => "110100110011111111110000",
31816 => "110010110010101011111100",
31817 => "101110111111000011000010",
31818 => "101100100011010011101000",
31819 => "101100001101000000010110",
31820 => "101100100111010111010110",
31821 => "101101010011000010001100",
31822 => "101110011001110100111000",
31823 => "110000000101000100110110",
31824 => "110001010001010110011100",
31825 => "110000110001111100101110",
31826 => "110000110100011111111100",
31827 => "110011011101000011110110",
31828 => "110110101011100010110000",
31829 => "111001010011110101011010",
31830 => "111100001010100010101001",
31831 => "111110010011001000000111",
31832 => "111110001110111100010001",
31833 => "111100000101110100100110",
31834 => "111001010111111010000000",
31835 => "111000000100010000101000",
31836 => "111000101111000010010010",
31837 => "111010101010001000100010",
31838 => "111101011111101000010001",
31839 => "000001001001000101010110",
31840 => "000101100101100000110000",
31841 => "001010011101111101001100",
31842 => "001110011011000110110000",
31843 => "010001010011010000000100",
31844 => "010100110101001000100000",
31845 => "011000110011101100011010",
31846 => "011010110000011110011111",
31847 => "011010001101010111000110",
31848 => "011000110000100010010011",
31849 => "010110010000110001001010",
31850 => "010001111000111010110000",
31851 => "001101100001100110010000",
31852 => "001011001011000011010111",
31853 => "001010100100010100010001",
31854 => "001011011110010110001101",
31855 => "001100110011010111110010",
31856 => "001100000111010001011000",
31857 => "001001100111110000100110",
31858 => "000111010011110010010110",
31859 => "000101101101101111101101",
31860 => "000101011101111000010110",
31861 => "000111001100110010110101",
31862 => "001001111001110111000100",
31863 => "001101000000011100011110",
31864 => "010000010110110001000110",
31865 => "010001101100110101100110",
31866 => "001111110000100111000000",
31867 => "001100110010000011000110",
31868 => "001010001011001100001100",
31869 => "000110110100110010100010",
31870 => "000001110110110001011001",
31871 => "111011011101000100010110",
31872 => "110101001101100000000110",
31873 => "110001010011111010001100",
31874 => "110000000110000101001000",
31875 => "110000000001011001000100",
31876 => "110000001011110010011100",
31877 => "110001110000001110010110",
31878 => "110101100110101110011100",
31879 => "111010100100111101101100",
31880 => "111110110011000001100101",
31881 => "000000011101001011111110",
31882 => "000000000010111101011011",
31883 => "000000001100111110011101",
31884 => "000001010000110101011100",
31885 => "000010110001001000101101",
31886 => "000101010110001111100111",
31887 => "001000000010000110100011",
31888 => "001001100101011101011110",
31889 => "001001100001000000011110",
31890 => "000111110100010011010010",
31891 => "000110001110101001010101",
31892 => "000100111110010011000100",
31893 => "000001100101000101111010",
31894 => "111011101010110101010010",
31895 => "110101101000011110110101",
31896 => "110001010010001000000000",
31897 => "101110010011101100010000",
31898 => "101011010110001111111000",
31899 => "100111111100111011001010",
31900 => "100101110100010100011111",
31901 => "100111101110011111101111",
31902 => "101101100010000010010000",
31903 => "110100100001010010010000",
31904 => "111100000100110010001111",
31905 => "000011111000000100001110",
31906 => "001001011111001101101101",
31907 => "001100100111100110111110",
31908 => "001111010000100000001000",
31909 => "010000111001100101100100",
31910 => "010000001000001010111000",
31911 => "001101100000100010001000",
31912 => "001000111100011001100101",
31913 => "000010110101111011010111",
31914 => "111110010101001101000100",
31915 => "111100000001001011101001",
31916 => "111001111000000100101000",
31917 => "111000011000111101111010",
31918 => "111000010011100001001110",
31919 => "111000111000111111001100",
31920 => "111010110111111110110000",
31921 => "111111000100110100000011",
31922 => "000011000000001100100000",
31923 => "000100000001010000100010",
31924 => "000011100101110001001110",
31925 => "000011001000011100011111",
31926 => "000010001011101011010001",
31927 => "000001101111000010101100",
31928 => "000001011010101001001001",
31929 => "000000101110111000010101",
31930 => "000010001100110101110010",
31931 => "000100111000001100001110",
31932 => "000110000000010010110001",
31933 => "000111010000000101000111",
31934 => "001001100110100000000010",
31935 => "001011100110001100110011",
31936 => "001100111100001000001010",
31937 => "001101001101011100110010",
31938 => "001011110010001011111010",
31939 => "001001110111001111111111",
31940 => "001000000010101011110010",
31941 => "000100010111011111101111",
31942 => "111110111111001110101001",
31943 => "111010001110101100110110",
31944 => "110101011100100111011000",
31945 => "110000010100000001111110",
31946 => "101100101111010011101010",
31947 => "101011001111100000101000",
31948 => "101100011011110100010110",
31949 => "110000001011110000101000",
31950 => "110100011100101001110010",
31951 => "111001010011110101101011",
31952 => "111111111101001110001001",
31953 => "000111111001111111000110",
31954 => "001111111100100110110110",
31955 => "010110101101001110010000",
31956 => "011010100111101001110001",
31957 => "011010100001100000011111",
31958 => "010111010110001001000110",
31959 => "010010011001010011110000",
31960 => "001011001101000110001111",
31961 => "000010100000001001101010",
31962 => "111010001000101111001001",
31963 => "110011100110011010100110",
31964 => "110000001001000011110010",
31965 => "101110010110000001111000",
31966 => "101100110010110110001100",
31967 => "101100110100000010000110",
31968 => "101110010001000101111100",
31969 => "101111101110000001100010",
31970 => "110000110111101001001010",
31971 => "110001101111101110111100",
31972 => "110010100101100100101000",
31973 => "110011110000001111000100",
31974 => "110101000101000000110010",
31975 => "110101001000011101011111",
31976 => "110011000000110110100000",
31977 => "110000011110000111100000",
31978 => "101111000101011100101010",
31979 => "101111010110100100100010",
31980 => "110001100101001111111010",
31981 => "110100001001110110001101",
31982 => "110101100000100100011001",
31983 => "110110001000011110011010",
31984 => "110110001100101111100110",
31985 => "110101011101000001000110",
31986 => "110100011011111001011110",
31987 => "110011101110101101101110",
31988 => "110011010111010011011000",
31989 => "110011011000011001111110",
31990 => "110011111101101101101000",
31991 => "110101100011000110010101",
31992 => "111000111001011010110011",
31993 => "111101001001001010011110",
31994 => "000000111011110001111111",
31995 => "000101100011010011110001",
31996 => "001011100111010101110101",
31997 => "010001000110110001001100",
31998 => "010100110010000111110000",
31999 => "010110011111100011010100",
32000 => "010101110111100011100110",
32001 => "010010110110100011010100",
32002 => "001110101011110001011100",
32003 => "001011001111101000000001",
32004 => "001001100101101001110011",
32005 => "001010011001100110110010",
32006 => "001100110101110101101000",
32007 => "001110100011000110111010",
32008 => "001111001001110001011000",
32009 => "001111010001011100101110",
32010 => "001110100111000111010110",
32011 => "001100111100000000000110",
32012 => "001010101110001110101101",
32013 => "001010011110111010000111",
32014 => "001101100010110100000010",
32015 => "010000100110110010000110",
32016 => "010000111111101101100100",
32017 => "001111100110011110100100",
32018 => "001101111110011111010100",
32019 => "001100101110001110000100",
32020 => "001011101001100001111010",
32021 => "001010111100010001100100",
32022 => "001010100000101100100010",
32023 => "001001100100111011101100",
32024 => "001000000110010111011010",
32025 => "000110001101011110001110",
32026 => "000100011110110000010001",
32027 => "000011110101001001001010",
32028 => "000011100111010110000010",
32029 => "000011000101001110101010",
32030 => "000010011010010110100110",
32031 => "000001101000100101110001",
32032 => "000000100111100000001001",
32033 => "111110100001001010011101",
32034 => "111010110010010100111011",
32035 => "110110101101100010111011",
32036 => "110100000111010001011011",
32037 => "110100000101011010100101",
32038 => "110110000000111101001101",
32039 => "110111101000110100000100",
32040 => "110111111100111110010010",
32041 => "111000001000000101110001",
32042 => "111000111101110110011101",
32043 => "111010001010111100101100",
32044 => "111011100001101111010010",
32045 => "111100011100110010011100",
32046 => "111011111011010011110000",
32047 => "111010011101001110111110",
32048 => "111001001110110111000110",
32049 => "110111110101011110101110",
32050 => "110101100101100011001000",
32051 => "110011000010111001011110",
32052 => "110000110101110100011110",
32053 => "101110111011110100111010",
32054 => "101101011001011011001000",
32055 => "101101001101011000010100",
32056 => "101111000000110110111100",
32057 => "110001010111011101110100",
32058 => "110011000100011001101000",
32059 => "110101011000010110111111",
32060 => "111001000001011110100111",
32061 => "111100111101111010000110",
32062 => "000000010111011100010101",
32063 => "000010010011100111010000",
32064 => "000010110010001111101010",
32065 => "000011001111111001101001",
32066 => "000011101101010000000000",
32067 => "000011011000100000100111",
32068 => "000010111110101100011000",
32069 => "000011100010000010010100",
32070 => "000101001011000000110100",
32071 => "000110111101000011010111",
32072 => "000111111111101100111100",
32073 => "001000011001011000011100",
32074 => "001000011101101010111000",
32075 => "001000001101011100110110",
32076 => "000110101010111101110100",
32077 => "000011010100000101100101",
32078 => "111111001011011011110111",
32079 => "111010000111000010011010",
32080 => "110100110111100011101100",
32081 => "110011000010101110001100",
32082 => "110101000111100001011100",
32083 => "111000110111000101111110",
32084 => "111101101011010101101110",
32085 => "000010100110110011100101",
32086 => "000110111011100010001011",
32087 => "001011110000010100110010",
32088 => "010000111001010000001000",
32089 => "010101001000110110101110",
32090 => "011000011011000100011011",
32091 => "011001100100000111100000",
32092 => "010110100001101010100110",
32093 => "010000111111110100111100",
32094 => "001100010100000100001010",
32095 => "000111111001011101101110",
32096 => "000001111111111111101110",
32097 => "111011011100011111000011",
32098 => "110101100111010000111110",
32099 => "110001110101010001010010",
32100 => "110000110110010000010000",
32101 => "110000011110100001010000",
32102 => "101111001101000110000100",
32103 => "110000001011101000011010",
32104 => "110101010100111111010100",
32105 => "111011100111011101010010",
32106 => "000001001110101001100011",
32107 => "000111011000110000000001",
32108 => "001110010011001000010010",
32109 => "010100000111100101101100",
32110 => "010110010000010101101110",
32111 => "010100100000011101001000",
32112 => "010001001111011010111100",
32113 => "001100111100011101010110",
32114 => "000110111100011001001101",
32115 => "000000100001011000110100",
32116 => "111011100101000010101111",
32117 => "111000111111000001111011",
32118 => "111000000110010001111010",
32119 => "110111100010111000110000",
32120 => "110111000011100011111011",
32121 => "110111101000000110111111",
32122 => "111001101111111011000110",
32123 => "111011110111101100101100",
32124 => "111100101011110001010001",
32125 => "111100110000000110110111",
32126 => "111011011101011100101000",
32127 => "110111011100000011010111",
32128 => "110001001010000110011010",
32129 => "101010010111000111101100",
32130 => "100101111110011101001000",
32131 => "100101111000110000100101",
32132 => "101000110100110010111010",
32133 => "101101110000010110000010",
32134 => "110100100110101111010001",
32135 => "111011111011011010101000",
32136 => "000001101100011001011000",
32137 => "000100101101101110011000",
32138 => "000101100111111110010010",
32139 => "000101100011011010011011",
32140 => "000011110100101011100010",
32141 => "000000011110111011101100",
32142 => "111101011000010011000010",
32143 => "111011010010110110110000",
32144 => "111010010010010100110101",
32145 => "111010010011011001101010",
32146 => "111011001000000101010110",
32147 => "111101011101101001001010",
32148 => "000001101001011110000001",
32149 => "000110111100110010100101",
32150 => "001011011011111001110101",
32151 => "001100001101110011010010",
32152 => "001001111001001010100100",
32153 => "000111100000000111111110",
32154 => "000101011011110110101000",
32155 => "000100000001000101001101",
32156 => "000100011010011011011011",
32157 => "000110010101011000111011",
32158 => "001001001001100110000101",
32159 => "001011101100000100010010",
32160 => "001100110011011101111000",
32161 => "001100000110000101001100",
32162 => "001000110101101000101101",
32163 => "000011110001010000111101",
32164 => "111111001011110101111001",
32165 => "111100111110010111001010",
32166 => "111101110011000001000111",
32167 => "000000010101100000000101",
32168 => "000011001101110110100001",
32169 => "000101010000001111011100",
32170 => "000101000111101101111000",
32171 => "000100011111100101101010",
32172 => "000101011010101101101000",
32173 => "000110101000111101011010",
32174 => "000110110100011001100000",
32175 => "000110001111000111001110",
32176 => "000101011000111100001010",
32177 => "000100010010000110111000",
32178 => "000011100011101000010010",
32179 => "000100010000000111101011",
32180 => "000101100111010001111001",
32181 => "000111000001100000001000",
32182 => "001000101011110010101100",
32183 => "001001001110110010100100",
32184 => "000111010010110100000100",
32185 => "000011000010111100111010",
32186 => "111110000101011101110001",
32187 => "111001110000100010110101",
32188 => "110110001111100100001011",
32189 => "110101100011001010110000",
32190 => "111001001110110011001110",
32191 => "111111010110000001010100",
32192 => "000101101010010011101100",
32193 => "001011000010110001000001",
32194 => "001111111111100011011110",
32195 => "010100011111101111110010",
32196 => "010110001010100001111100",
32197 => "010100110110100010110110",
32198 => "010001110100110111011100",
32199 => "001101011110110011111010",
32200 => "001000100011000101010100",
32201 => "000010100000111100001011",
32202 => "111011111000111010111010",
32203 => "110110000111010111001010",
32204 => "110000111111010000111100",
32205 => "101100111101001010100110",
32206 => "101001001010000110011110",
32207 => "100100110010110001010001",
32208 => "100010001111101100111111",
32209 => "100010011001101111110001",
32210 => "100011111100011010101001",
32211 => "100100100110001000000000",
32212 => "100101100010101100010101",
32213 => "101100011111110110110100",
32214 => "110111000000000000000001",
32215 => "111110110010001111010110",
32216 => "000101000010000110101111",
32217 => "001001110111010001100111",
32218 => "001100010001001111010100",
32219 => "001100111011000011010010",
32220 => "001010010101000100101100",
32221 => "000101111110010011001101",
32222 => "000010100011000101101100",
32223 => "000000000011011100110111",
32224 => "111111000000000001101000",
32225 => "111110011011001110111111",
32226 => "111101000110101000000010",
32227 => "111011010000101110100100",
32228 => "111001011100111000010000",
32229 => "111000110011001001111010",
32230 => "110110111000010111010100",
32231 => "110001111000001000010110",
32232 => "101101101100100100001110",
32233 => "101100001100111111110010",
32234 => "101100111110110100000010",
32235 => "110000010011101010101010",
32236 => "110101010010000110000110",
32237 => "111100011011111001011111",
32238 => "000101110011001111101111",
32239 => "001111010000110101011010",
32240 => "010111101101000101000010",
32241 => "011101001001110001100000",
32242 => "011110010001111100010001",
32243 => "011101011111111000110100",
32244 => "011100010111111010110101",
32245 => "011000101001110101110100",
32246 => "010000110100001001000000",
32247 => "001000100001111110111001",
32248 => "000010110011000010111111",
32249 => "111100100100000110111101",
32250 => "110101010011000110001000",
32251 => "110001011111000010100010",
32252 => "110001100010110011101110",
32253 => "110010010010100010010110",
32254 => "110010011000011101111110",
32255 => "110010001101111010011010",
32256 => "110011101001001000111110",
32257 => "111000100101101101100010",
32258 => "000000000110101010010100",
32259 => "000111001100011000011011",
32260 => "001101000001100000110010",
32261 => "010011101001110100101000",
32262 => "011010010011000110011011",
32263 => "011101000001100101110101",
32264 => "011011110110000110110101",
32265 => "011000100011001110010010",
32266 => "010010100100000001000010",
32267 => "001010110010000000111000",
32268 => "000010001001001100001110",
32269 => "111001000011001000001111",
32270 => "110010110011100111110110",
32271 => "110000001100010000100010",
32272 => "101110010010011011110100",
32273 => "101100111001000000100110",
32274 => "101101101111011000101110",
32275 => "110001010110110100101100",
32276 => "110101100110110011010100",
32277 => "110111101001110000110110",
32278 => "110111110111001011001010",
32279 => "110111000000001001111010",
32280 => "110011100110011000100100",
32281 => "101100111011111101010010",
32282 => "100110010101010010100011",
32283 => "100100011000011100011010",
32284 => "100101101110000011110011",
32285 => "101000001010111001010000",
32286 => "101110101100010011100100",
32287 => "111000001100001111111000",
32288 => "000000000110100000000010",
32289 => "000101101001111101110000",
32290 => "001000100100111101110101",
32291 => "001001000100101000110101",
32292 => "001000001011110101011000",
32293 => "000101100011001001011100",
32294 => "000001101101110111011101",
32295 => "111101011111000010110100",
32296 => "111001000110001001101011",
32297 => "110101001100001000001000",
32298 => "110001110101100100000010",
32299 => "110000011000111111011110",
32300 => "110010101110110000001100",
32301 => "110111110101011000100111",
32302 => "111101011010011100010101",
32303 => "000010001111100101001100",
32304 => "000110000010001010101100",
32305 => "001000010110111001111110",
32306 => "001000110011111111111011",
32307 => "001000011000011101011011",
32308 => "001000101111100111100011",
32309 => "001010101111000101000101",
32310 => "001101010101010010000100",
32311 => "001110110001100101010100",
32312 => "001110110010010000000100",
32313 => "001101101000101100001000",
32314 => "001011010111101110101100",
32315 => "000111111100000011111010",
32316 => "000011110111011100001100",
32317 => "000001010111010010001100",
32318 => "000000100010000000001111",
32319 => "111111001101010011010011",
32320 => "111110011010000010101100",
32321 => "111111011111000000010000",
32322 => "000000010100110000011110",
32323 => "111111001100001110011111",
32324 => "111101011101111101001100",
32325 => "111101010101110110100000",
32326 => "111110010010100011011000",
32327 => "111110010110101100011001",
32328 => "111101100101001010010000",
32329 => "111101010110101110101111",
32330 => "111110010010011100101100",
32331 => "111111100001101001001011",
32332 => "000001000110000110010101",
32333 => "000100010101111101000010",
32334 => "001000001010011000101010",
32335 => "001010101100100110001110",
32336 => "001011110000010010001100",
32337 => "001010101000110011101011",
32338 => "000111010111000011011000",
32339 => "000011001100010100101001",
32340 => "111110111101010110111010",
32341 => "111011101000000110011100",
32342 => "111010001100001000000111",
32343 => "111011010000101100010110",
32344 => "111110101000010010011100",
32345 => "000011010101000100100111",
32346 => "001000111010111001111100",
32347 => "001110100010100101001100",
32348 => "010010110110110000001110",
32349 => "010101001111111000010000",
32350 => "010101100110011111101010",
32351 => "010100111110000001001010",
32352 => "010100011010110100101100",
32353 => "010011100000100101011000",
32354 => "010001100101011000010100",
32355 => "001110010100100100101100",
32356 => "001001110111011101101001",
32357 => "000100100110010010010110",
32358 => "111110110100011100000000",
32359 => "111001011010110100100110",
32360 => "110101000101010010011011",
32361 => "110010001010011010010000",
32362 => "110000110100100101001000",
32363 => "110000110010101000111010",
32364 => "110010101111000011010010",
32365 => "110111010001100100100110",
32366 => "111110000111101100111110",
32367 => "000110001111100000011110",
32368 => "001100101100011100011110",
32369 => "010000001010010001100110",
32370 => "010010000110010010101110",
32371 => "010010001110011100001110",
32372 => "001111101111001001010110",
32373 => "001010101010010100111000",
32374 => "000011011011001110000101",
32375 => "111100111000100101000001",
32376 => "111001010111001010010001",
32377 => "110111011011101100111100",
32378 => "110100111011100011010000",
32379 => "110010010111001100110110",
32380 => "110001010001011110111110",
32381 => "101111111010001100101000",
32382 => "101101000000101001010000",
32383 => "101010111000110111011000",
32384 => "101001000100110011010000",
32385 => "100110111100010010001000",
32386 => "100111101110010010010101",
32387 => "101011011000011010001000",
32388 => "101111100101001011110110",
32389 => "110100100101001000110000",
32390 => "111010110010111111110000",
32391 => "000010101100000100100110",
32392 => "001011111001001001011110",
32393 => "010011011011001100101000",
32394 => "010111101110101101100010",
32395 => "011010000111110011111111",
32396 => "011010000101011001101000",
32397 => "010101011101110110010100",
32398 => "001110000000101010110000",
32399 => "000110011100110101101101",
32400 => "111110000110110000111011",
32401 => "110110011111100000000001",
32402 => "110001110101111111110110",
32403 => "101110001111101011010010",
32404 => "101100010010001000001100",
32405 => "101110001110101111010100",
32406 => "110001100100111011010010",
32407 => "110011111111011100111110",
32408 => "110111001011111010111100",
32409 => "111100110111111001100000",
32410 => "000011001111110001011001",
32411 => "001000100100101001001100",
32412 => "001110011100000010001110",
32413 => "010100000000010100010100",
32414 => "010111011010000000110100",
32415 => "011010001100010011001001",
32416 => "011011101001010100000111",
32417 => "011010111101010111100001",
32418 => "011001001010111100001111",
32419 => "010011110101101100000100",
32420 => "001011101000111100011111",
32421 => "000101000000000101101010",
32422 => "111111001010011001011001",
32423 => "111000011101000010001100",
32424 => "110010010001110000100100",
32425 => "101110010100010101111000",
32426 => "101101101010100100100010",
32427 => "101111101010001111011100",
32428 => "110011011000100101001100",
32429 => "111000010000111010110110",
32430 => "111100100111101100110101",
32431 => "111110110000110000011100",
32432 => "111101001011110011101011",
32433 => "111000000100101001110100",
32434 => "110001110011010100110000",
32435 => "101100010100111110010010",
32436 => "101001010110011110011000",
32437 => "101001001100010101001100",
32438 => "101010111111110010101010",
32439 => "101111001111001000010000",
32440 => "110100011010001000111010",
32441 => "110111100111110111100100",
32442 => "111001010110001010000011",
32443 => "111011010001101100111110",
32444 => "111101111010010101100111",
32445 => "000000010010111101001110",
32446 => "000000111111101101011111",
32447 => "000000100000010001100111",
32448 => "111110110101000001011011",
32449 => "111010011111000000011101",
32450 => "110100110101010101011110",
32451 => "110001001101011001111010",
32452 => "110000101011011111100000",
32453 => "110010001100000011000010",
32454 => "110100110100100010000110",
32455 => "111000010001011010101110",
32456 => "111011101110100101111111",
32457 => "111110011010100000011100",
32458 => "000000110110000111001010",
32459 => "000011010101110110110000",
32460 => "000101101111000100111100",
32461 => "001001000010111011111010",
32462 => "001101011010011110010100",
32463 => "010000110010110000011000",
32464 => "010010000110101000101000",
32465 => "010001011011111000111110",
32466 => "001110010010011101000010",
32467 => "001000101011001110010001",
32468 => "000010000111011101110101",
32469 => "111101001011000001100000",
32470 => "111011010110101101000011",
32471 => "111011101001101100000011",
32472 => "111100011001100011010010",
32473 => "111100101011100100010101",
32474 => "111100011101000110010000",
32475 => "111100001110111101101110",
32476 => "111100001000010101010000",
32477 => "111100100000010001001001",
32478 => "111101101111111011001100",
32479 => "111111010000101100111001",
32480 => "000000010011010001100111",
32481 => "000000100000010110011101",
32482 => "000000001111011100110111",
32483 => "000000000011110100111111",
32484 => "000000000101001010011101",
32485 => "000001000101101101000100",
32486 => "000011000110110000100001",
32487 => "000100110010100110101100",
32488 => "000101011000001111001000",
32489 => "000100001101011001000101",
32490 => "000001000010110001011001",
32491 => "111100100010100110110001",
32492 => "110111110101111000100000",
32493 => "110101000001110010110111",
32494 => "110100111100010000100110",
32495 => "110110100010101000101010",
32496 => "111001001001010101111111",
32497 => "111100101001110000000111",
32498 => "000000111011001101110111",
32499 => "000100011001010000100000",
32500 => "000101110000010000011000",
32501 => "000110100111111101100001",
32502 => "001000000010001010101001",
32503 => "001001010100101110010100",
32504 => "001010001001010101010100",
32505 => "001010010100110010100011",
32506 => "001010101001101101000100",
32507 => "001011010100100011010011",
32508 => "001011010000011001000100",
32509 => "001010000001101000011000",
32510 => "000111010001110111111000",
32511 => "000011100011110001100011",
32512 => "111111011110100111100100",
32513 => "111010001111101110001101",
32514 => "110100100000111000000000",
32515 => "101111101011110111111000",
32516 => "101100110000101010000000",
32517 => "101101001101010100101100",
32518 => "110001001111100100000010",
32519 => "111000001111100001101111",
32520 => "000001000000000011000010",
32521 => "001001010101011111110100",
32522 => "001111010110010111010000",
32523 => "010001100011110010000110",
32524 => "010001000100101000001110",
32525 => "001111110111110100100100",
32526 => "001100110000110001011000",
32527 => "000111101010010101110110",
32528 => "000010101011111100111001",
32529 => "111110111011001011010000",
32530 => "111101101001101110010011",
32531 => "111111001111101001001010",
32532 => "000010000110110000111001",
32533 => "000100100111101111100110",
32534 => "000110000011100111000010",
32535 => "000110001100111110101100",
32536 => "000100011111111011010100",
32537 => "000001110101110101111010",
32538 => "111111111001001100111100",
32539 => "111101100110011000110010",
32540 => "111010100011101000111111",
32541 => "111000110011000000001010",
32542 => "111001001100000111001010",
32543 => "111011011010100001101110",
32544 => "111110111000111110011101",
32545 => "000010110110010010101100",
32546 => "000110010011101100110000",
32547 => "001000001001001101001111",
32548 => "001000010000000100111011",
32549 => "000111000011100111011110",
32550 => "000101000110101110000111",
32551 => "000011000010000101001010",
32552 => "000001000100101110001011",
32553 => "111111100010000101101110",
32554 => "111101101111101101011111",
32555 => "111011100101100001111011",
32556 => "111011011111100100100110",
32557 => "111101101100111100010000",
32558 => "111111101110100101001011",
32559 => "000001100010011011110010",
32560 => "000100001101110100111001",
32561 => "000110101001110110001001",
32562 => "000111101100101000011111",
32563 => "001000001110010111000011",
32564 => "001000010110000100011101",
32565 => "000111010101111101010010",
32566 => "000110101110011101111000",
32567 => "000111000001111011110000",
32568 => "000111000100100110101101",
32569 => "001000000111100001101000",
32570 => "001010111100101010101101",
32571 => "001101001101011111111110",
32572 => "001101011011110101011010",
32573 => "001101010000000110100110",
32574 => "001110001111110011001110",
32575 => "001110011110101111101010",
32576 => "001011100111100111001010",
32577 => "000111000010110010101100",
32578 => "000011111101110010010111",
32579 => "000011101001001001101011",
32580 => "000011111110010110010001",
32581 => "000011101000000100010111",
32582 => "000011101111110001000001",
32583 => "000011001001001010110010",
32584 => "111111100101010000110000",
32585 => "111001011000011011110001",
32586 => "110010001110001000110110",
32587 => "101100100111100011011100",
32588 => "101001111100111001100110",
32589 => "101001100001000011110100",
32590 => "101011000000100000010010",
32591 => "101110100000000000110100",
32592 => "110011001101011011000010",
32593 => "110111100101111001011000",
32594 => "111010110010101001000110",
32595 => "111101100011111100000010",
32596 => "000001011001001011000000",
32597 => "000110110110001110001010",
32598 => "001011100011101101000010",
32599 => "001101011111101100011100",
32600 => "001101100100110000010100",
32601 => "001011010010100001000100",
32602 => "000101111010011010111010",
32603 => "111110110111111001001000",
32604 => "110111111011001001110110",
32605 => "110011100001010001111000",
32606 => "110000110000101101010110",
32607 => "101100110000101100011110",
32608 => "101010000010001001000000",
32609 => "101010010010011010000000",
32610 => "101010111001000101101100",
32611 => "101011110101011001110000",
32612 => "101111100101100011010110",
32613 => "110110110010101011000101",
32614 => "111110110011001001111010",
32615 => "000101110101100001000110",
32616 => "001100100111000110000110",
32617 => "010000100110111110101000",
32618 => "001111101110100011011000",
32619 => "001100011001000101011100",
32620 => "000111101000100100011111",
32621 => "000001110110000111010111",
32622 => "111101001101100010000011",
32623 => "111010011001011100110000",
32624 => "111000100111001101010111",
32625 => "110111101000101110110101",
32626 => "110111010111010001000101",
32627 => "110110011101111001101000",
32628 => "110101000100110110001100",
32629 => "110101111110110011000100",
32630 => "111001100111000111100101",
32631 => "111110010101000100001010",
32632 => "000010010111111000010010",
32633 => "000011011001001000010011",
32634 => "000010110000001100110100",
32635 => "000011001101011011000000",
32636 => "000011011101101110110011",
32637 => "000010110101010111010110",
32638 => "000010111001001111011011",
32639 => "000011011100001111000111",
32640 => "000010101101100101001011",
32641 => "000000001110011111111010",
32642 => "111101011111001011101110",
32643 => "111011000011100101001000",
32644 => "111000100011100010100011",
32645 => "110111010100010000000011",
32646 => "111000001001010100010100",
32647 => "111010000000110000110110",
32648 => "111100011011000011101010",
32649 => "111111100010110000010110",
32650 => "000010110111110101010000",
32651 => "000101010101011010101000",
32652 => "000110010010011000111010",
32653 => "000110000110010010000010",
32654 => "000110001011110011111100",
32655 => "000111010000111010110000",
32656 => "000111101100101100101100",
32657 => "000110100110000011010011",
32658 => "000101011010111011000001",
32659 => "000100111001001100110000",
32660 => "000100101000110000010011",
32661 => "000100010010011010110101",
32662 => "000011010111100010010110",
32663 => "000001111000010100100000",
32664 => "000000001011111100101000",
32665 => "111101111111101001010110",
32666 => "111010100110111010011010",
32667 => "110110011111100101111101",
32668 => "110010100000100110110010",
32669 => "101110101000100110011010",
32670 => "101100001011001001111100",
32671 => "101100110110001101010000",
32672 => "101111110001100011110110",
32673 => "110011011000001011000010",
32674 => "110111010011110111011101",
32675 => "111011111001111001010111",
32676 => "000000001000001000010011",
32677 => "000001101010000000000111",
32678 => "000000111110100001110010",
32679 => "111111101101010010000011",
32680 => "111101101000100010010010",
32681 => "111011110100101100011010",
32682 => "111011010011111101101000",
32683 => "111011000111110111000101",
32684 => "111011101100001111001100",
32685 => "111110010100001001110010",
32686 => "000001111010111010011010",
32687 => "000100010101111011001010",
32688 => "000101100111000001110110",
32689 => "000110100100111111000010",
32690 => "000110011110010011110010",
32691 => "000101110010110111011001",
32692 => "000101100000111000001001",
32693 => "000011111101011111110110",
32694 => "000001000100011111101110",
32695 => "111110111101001000010011",
32696 => "111101101000010110010001",
32697 => "111100101111001111001100",
32698 => "111101010110111000101100",
32699 => "000000010110100100001101",
32700 => "000110000110010100011010",
32701 => "001101110000100011010010",
32702 => "010100000111000001101010",
32703 => "010110111100111111010010",
32704 => "010111110111101101010000",
32705 => "011000000100011100110111",
32706 => "010111000000101001010000",
32707 => "010100100111001110101000",
32708 => "010000010010101010101000",
32709 => "001011001100010000101000",
32710 => "001000001001111110101110",
32711 => "000110001000101101110100",
32712 => "000010101111000100101111",
32713 => "111111000001101001001110",
32714 => "111101101001101110101101",
32715 => "111111010110111011011100",
32716 => "000001001110011100100000",
32717 => "000000100001100100011101",
32718 => "111101111001010001011101",
32719 => "111011000011001001100100",
32720 => "111001110101110010100001",
32721 => "111010010110010110100010",
32722 => "111011001000111101101100",
32723 => "111101001110101010011011",
32724 => "000001010000011001110100",
32725 => "000101101000000101110111",
32726 => "001001111100111111100001",
32727 => "001101110100111101110100",
32728 => "001111111001110111101100",
32729 => "001111110010101111000100",
32730 => "001101100110100111001110",
32731 => "001010000110110101100011",
32732 => "000110110011011111111111",
32733 => "000011100000111011000110",
32734 => "111111000010100010100010",
32735 => "111001111111011111011000",
32736 => "110011111110000101010110",
32737 => "101011011111010100101000",
32738 => "100100000100100100100110",
32739 => "100001100110101010110001",
32740 => "100001110101111001111001",
32741 => "100010011111111000001110",
32742 => "100011110100100000101001",
32743 => "100110111011000110001001",
32744 => "101101110010111010001010",
32745 => "110110010010000001101000",
32746 => "111011110010111111111000",
32747 => "111111101100001100001100",
32748 => "000101100010111011111110",
32749 => "001100000010111000100100",
32750 => "010000010110000001100000",
32751 => "010010010111011010010010",
32752 => "010010101001101010101100",
32753 => "010000111101011010010000",
32754 => "001101000101101100111110",
32755 => "000111001010000001011110",
32756 => "000001100100110111100001",
32757 => "111110010110001010100101",
32758 => "111010101010111010100110",
32759 => "110101010010001011000100",
32760 => "110001011110101001011100",
32761 => "110000001111000011110110",
32762 => "101111100011010101101110",
32763 => "101110100100101000001000",
32764 => "101111000110111001010010",
32765 => "110011101101010011110100",
32766 => "111011111111110011000111",
32767 => "000101010010101011001100",
32768 => "001101000100011111110110",
32769 => "010010010111111100010010",
32770 => "010101100000111010111100",
32771 => "010101011101110010011000",
32772 => "010010001100000101000010",
32773 => "001110111110101000110100",
32774 => "001101101001100111010000",
32775 => "001100011101100000011000",
32776 => "001001011101000101110001",
32777 => "000101001010101000111001",
32778 => "000001000001001011001000",
32779 => "111100110100101011100111",
32780 => "111001010010111100111110",
32781 => "110111100100011101110001",
32782 => "110110010100010110111110",
32783 => "110101001101001101001000",
32784 => "110101110000110011111101",
32785 => "111000011001001101111100",
32786 => "111100001011111000000101",
32787 => "111111000010111000011111",
32788 => "111111100101110011010111",
32789 => "111111011110011101001010",
32790 => "000001000101111101100000",
32791 => "000011010101110100010110",
32792 => "000011001000010100011110",
32793 => "000001100000111010100011",
32794 => "000001010110100001001110",
32795 => "000001010110101011110100",
32796 => "111111101010111101011110",
32797 => "111101110001100001001101",
32798 => "111110101010101011100110",
32799 => "000011001101011000010101",
32800 => "001000010001100111001010",
32801 => "001011100000111000101010",
32802 => "001101101110010101001000",
32803 => "001111000010111100101100",
32804 => "001110100011001100011000",
32805 => "001100000011011010001000",
32806 => "001000010111100111101010",
32807 => "000100001101101111011000",
32808 => "000000000100101110101010",
32809 => "111101000101010111001000",
32810 => "111011001100000011110000",
32811 => "111010010000100011011101",
32812 => "111011111101111000001001",
32813 => "111111110110000011000110",
32814 => "000100000001000010101111",
32815 => "001000010001011110011000",
32816 => "001011110011000110111110",
32817 => "001101000111010100110010",
32818 => "001011101100000011111100",
32819 => "001000000110000000101100",
32820 => "000011011000010110000110",
32821 => "111110001011001011000000",
32822 => "111001011011100100111100",
32823 => "110101001100010111100110",
32824 => "110000011111100000110100",
32825 => "101100000100000110001000",
32826 => "101000011111011001000100",
32827 => "100101100010000011101001",
32828 => "100100001100010001000111",
32829 => "100101000110100000111110",
32830 => "100111100100000001010011",
32831 => "101001111000010110001110",
32832 => "101010111001101011110110",
32833 => "101100100001010110000100",
32834 => "110000101100101101011010",
32835 => "110101111010100110010010",
32836 => "111001110111111011010000",
32837 => "111100001111010100010000",
32838 => "111101010011111011001111",
32839 => "111101101111001100011000",
32840 => "111111000110100111111101",
32841 => "000000110110100100010110",
32842 => "000001011101010111000000",
32843 => "000001111001010011100010",
32844 => "000001011111010010000111",
32845 => "111111000111111100101011",
32846 => "111101001011100011101100",
32847 => "111011011100111011111011",
32848 => "110111110011001010011011",
32849 => "110011111011000100100100",
32850 => "110001110010001111010110",
32851 => "110001111100000000011000",
32852 => "110101000100101111110101",
32853 => "111010011011110011010111",
32854 => "000000101011101100101010",
32855 => "000111110001101100000010",
32856 => "001111010011110000001010",
32857 => "010101111001000101110000",
32858 => "011011001011010101011101",
32859 => "011110011111110101010000",
32860 => "011110101111000111000100",
32861 => "011101101011010100010001",
32862 => "011011100010011010100101",
32863 => "010101101010100000101000",
32864 => "001110011010011001101010",
32865 => "001001010111011001000001",
32866 => "000101010011000110111010",
32867 => "000001101101101110011001",
32868 => "000000010100110000011111",
32869 => "000001101001110100111100",
32870 => "000100100010011001100110",
32871 => "000111011000010100010111",
32872 => "001001011100101111110010",
32873 => "001010110000110010100011",
32874 => "001100111000100000100000",
32875 => "010000100011001100010010",
32876 => "010010110110101110111010",
32877 => "010011011000101101111000",
32878 => "010101000110000000010000",
32879 => "010111001000111111100000",
32880 => "010110110111111110010000",
32881 => "010011101111101110000100",
32882 => "001110001100011000011110",
32883 => "001000001100000110110000",
32884 => "000011010110111110100010",
32885 => "111110011100000000011001",
32886 => "111000101010110001010010",
32887 => "110010000101011100001100",
32888 => "101001100101111011000100",
32889 => "100010100000011001111011",
32890 => "100001010111101001110101",
32891 => "100010001010000100000001",
32892 => "100001011000110010111111",
32893 => "100001101100100100101111",
32894 => "100010011001000101000101",
32895 => "100100010010000110010011",
32896 => "101011010011100001110110",
32897 => "110011110101011000001010",
32898 => "111001010000000011100001",
32899 => "111101001100110110100001",
32900 => "000000111010011111001110",
32901 => "000100000010100100100110",
32902 => "000110011101101111101011",
32903 => "000111101000000101001110",
32904 => "000111000101010010001101",
32905 => "000100101001100001001100",
32906 => "000000111000111111111010",
32907 => "111100111110111010010000",
32908 => "111001101010000101110000",
32909 => "110111000011011010001010",
32910 => "110101000100110101001110",
32911 => "110011101000101000101100",
32912 => "110010001110000100010100",
32913 => "110000110110111000001010",
32914 => "110000010000111101100010",
32915 => "110000010001101011100110",
32916 => "110001010100110100010000",
32917 => "110100101010101111010000",
32918 => "111010101011110110010011",
32919 => "000011001011010010001010",
32920 => "001100010111001100110000",
32921 => "010011100100001110010010",
32922 => "010111000111011010111000",
32923 => "010110010111010110001010",
32924 => "010011011001110111110010",
32925 => "010001001110111100011110",
32926 => "001111101010011101001000",
32927 => "001101011000100011000110",
32928 => "001010011101110011110001",
32929 => "000111110010100100000000",
32930 => "000101111110111101110101",
32931 => "000100010110010010111110",
32932 => "000001011001111100111110",
32933 => "111101000101010010010110",
32934 => "111010000000111000110110",
32935 => "111010001001101111101001",
32936 => "111011111000001001100110",
32937 => "111101011101010101101100",
32938 => "111110111100000101011110",
32939 => "000001000111001000001010",
32940 => "000100010011110111011110",
32941 => "000110110000110110011100",
32942 => "000111101000110000110000",
32943 => "001000010101001010100000",
32944 => "001000110100000110000010",
32945 => "000111111011101000010110",
32946 => "000100100110000101100100",
32947 => "111110111000111011011111",
32948 => "111001000101000110111000",
32949 => "110100110000101110010111",
32950 => "110010111001111101110100",
32951 => "110100100000010010001110",
32952 => "111000011100000010111000",
32953 => "111101001100010000110001",
32954 => "000010000111101100011110",
32955 => "000110001000101101111000",
32956 => "000111110100010001010100",
32957 => "000110011100001110111111",
32958 => "000011010000011001111011",
32959 => "111111110101100100011100",
32960 => "111100100001010100111101",
32961 => "111001101000110100111000",
32962 => "110111001001101110000011",
32963 => "110101101101101001110100",
32964 => "110110111111101111100110",
32965 => "111010010011011000001111",
32966 => "111101111000000011110001",
32967 => "000001111111000101111001",
32968 => "000110111010011101111001",
32969 => "001011011000010100100010",
32970 => "001110010110011101010000",
32971 => "001111011100001001000100",
32972 => "001101101101000010111110",
32973 => "001001110001000110001000",
32974 => "000101101101001000110001",
32975 => "000000111001001100010010",
32976 => "111010011111111000101110",
32977 => "110011111011001110001000",
32978 => "101101011001000111110010",
32979 => "100111011011001001001010",
32980 => "100100011101010111011001",
32981 => "100100100111111100000110",
32982 => "100101100010001011100111",
32983 => "100111001011101111100011",
32984 => "101011011100100010100000",
32985 => "110001000000110001010110",
32986 => "110110000110001111110000",
32987 => "111011101111011011100110",
32988 => "000000101010101000011001",
32989 => "000010100000010110001110",
32990 => "000010011000110100000000",
32991 => "000001100101111101111011",
32992 => "000000011111000010101000",
32993 => "111111101001000011111111",
32994 => "111111001011100110011111",
32995 => "111111011011101110010110",
32996 => "000000011111101011100011",
32997 => "000001111101101110000111",
32998 => "000010110001000000001011",
32999 => "000001111011001011111101",
33000 => "000000111010101011000010",
33001 => "000000001000100100111110",
33002 => "111101100101110111100101",
33003 => "111010010111111111001100",
33004 => "111000101001100011101100",
33005 => "111000000100000111111110",
33006 => "111000110011110001101110",
33007 => "111011100000111010000010",
33008 => "111111001101010001001110",
33009 => "000011011110000101001001",
33010 => "001000111111100110011011",
33011 => "001110111100111011110100",
33012 => "010100001110000111110000",
33013 => "011000110110010101011100",
33014 => "011011011111010111110001",
33015 => "011011001110010110000011",
33016 => "011001000111110100100000",
33017 => "010100101110011010000000",
33018 => "001110100011110010001100",
33019 => "001010000000001111001010",
33020 => "000111110101100010100110",
33021 => "000110010111110000010000",
33022 => "000101101001001100011000",
33023 => "000110011100000100101010",
33024 => "001000000011001010111001",
33025 => "001001100111110000011101",
33026 => "001011010111110111011100",
33027 => "001101000101011000010000",
33028 => "001110111001000100010000",
33029 => "010001100111111011111100",
33030 => "010100100101000010000100",
33031 => "010111010001011001011010",
33032 => "011001011110011011010010",
33033 => "011001001000111001111101",
33034 => "010101111010001111001100",
33035 => "010010000010011101011100",
33036 => "001110101001111000010000",
33037 => "001010111110001010110000",
33038 => "000110010000110001100001",
33039 => "000001011011001111110100",
33040 => "111100111001110010010010",
33041 => "110111101000010101001100",
33042 => "110001101101111101100010",
33043 => "101100111010010010000110",
33044 => "101011100011101111100100",
33045 => "101101110001111010101110",
33046 => "110000010110000100010010",
33047 => "110010001001101000100010",
33048 => "110100100010101010100101",
33049 => "110110100011110001000110",
33050 => "110110100011101111111000",
33051 => "110101001011111101011101",
33052 => "110100101101110101111001",
33053 => "110110001011000100100111",
33054 => "111000000110101010001001",
33055 => "111001011000100110100010",
33056 => "111010000010000001111000",
33057 => "111001111100010110100111",
33058 => "111000110101001101011011",
33059 => "110110011000000001110010",
33060 => "110011111110011010110100",
33061 => "110100010000101010000100",
33062 => "110110101111111101011010",
33063 => "110111110110010110000000",
33064 => "110101111111111100101100",
33065 => "110011011000001010011110",
33066 => "110001101100001111100000",
33067 => "110000010110011101110010",
33068 => "101111001111100101000000",
33069 => "101111110000111110001000",
33070 => "110011010111101100001110",
33071 => "111000111001001110101101",
33072 => "111101100101010111010100",
33073 => "000001110110001110011010",
33074 => "000110010001010010110011",
33075 => "000111101111110010011110",
33076 => "000101001100110010000001",
33077 => "000010100001100000011110",
33078 => "000011010100011001110100",
33079 => "000110001101110111001001",
33080 => "000111100011111101001010",
33081 => "000111011111010011110010",
33082 => "001000000011001001111001",
33083 => "001000010100111111111101",
33084 => "000110011110110000010110",
33085 => "000011011001010000101100",
33086 => "000001100000001010010010",
33087 => "000000110101101011000100",
33088 => "000000011001011101001011",
33089 => "000001000101011010011011",
33090 => "000010001111110110101100",
33091 => "000010010011000011011011",
33092 => "000010101011101011110100",
33093 => "000100011111001111101001",
33094 => "000110111011111010100101",
33095 => "001001110011111100101000",
33096 => "001100001001101010110110",
33097 => "001100000001001011000110",
33098 => "001001011000100101011000",
33099 => "000110000011100011011011",
33100 => "000010011111001110101100",
33101 => "111110100111111011000101",
33102 => "111100100000111100010000",
33103 => "111101001110011000011010",
33104 => "111111000111001101001010",
33105 => "000000110001100101001000",
33106 => "000010010011010101101100",
33107 => "000100111000011011011011",
33108 => "001000010011001000010111",
33109 => "001010010011011001001001",
33110 => "001010011000011100000000",
33111 => "001001011010111110001010",
33112 => "000111011100000101101010",
33113 => "000100110001100000011110",
33114 => "000010000110101001011110",
33115 => "111111010101111100000011",
33116 => "111011111101100101001101",
33117 => "111000100010111000100010",
33118 => "110110110100110000001000",
33119 => "110110111101101000010001",
33120 => "110111110011111000100000",
33121 => "111001011000100101101110",
33122 => "111100000000100010101110",
33123 => "111111010010101001010100",
33124 => "000010110111101011101000",
33125 => "000101111110101000110001",
33126 => "000111011101111011100000",
33127 => "000111011001010100110111",
33128 => "000101101110110111000011",
33129 => "000001001101100001000010",
33130 => "111010000010001010010111",
33131 => "110001000100001110101010",
33132 => "100111101110110011011101",
33133 => "100010011110010000101101",
33134 => "100010011010001001110001",
33135 => "100011100000000001011000",
33136 => "100100010000001000000100",
33137 => "100100110110011001010110",
33138 => "100110100101001001100011",
33139 => "101100100011101100111100",
33140 => "110100110100000100010000",
33141 => "111011100001011011111110",
33142 => "000001000110010111010011",
33143 => "000100110101110100010000",
33144 => "000101100101110100110101",
33145 => "000100011101101101010000",
33146 => "000001001011110011001101",
33147 => "111100110010010100110011",
33148 => "111010111000110001001011",
33149 => "111011011001011001011110",
33150 => "111011111111001001111101",
33151 => "111101001101111111001011",
33152 => "111111001011100110011010",
33153 => "111111111100100010010111",
33154 => "111111101111001111001001",
33155 => "111111011101001101111100",
33156 => "111110010010011100001000",
33157 => "111100100101000011101100",
33158 => "111011001110100010101101",
33159 => "111001110110011011000001",
33160 => "111001100100101101101110",
33161 => "111100011011000010101011",
33162 => "000001001000100111000111",
33163 => "000101100101011110001100",
33164 => "001010111000101000111111",
33165 => "010001001011010010101110",
33166 => "010101110011011001010110",
33167 => "011000001100010100111111",
33168 => "011000100100110010001011",
33169 => "010110011101100000011100",
33170 => "010011000110100100010000",
33171 => "001110011001100101011110",
33172 => "000111111000010000101001",
33173 => "000011000101111111011100",
33174 => "000001111000010001110110",
33175 => "000001011110110111000001",
33176 => "000000010110110111110110",
33177 => "111111001010010110100101",
33178 => "111110101001111111001100",
33179 => "111111011110001000111111",
33180 => "000000110010000100101001",
33181 => "000000110110111000001000",
33182 => "000001010000001100110000",
33183 => "000100111110010110110000",
33184 => "001001011001111110000100",
33185 => "001010001000110011110101",
33186 => "001000110001011110111110",
33187 => "001000100011000011110010",
33188 => "001000111011100101001110",
33189 => "001000001100011110111101",
33190 => "000110001100101100010000",
33191 => "000011101010001111001101",
33192 => "111111101011100010010011",
33193 => "111000100100001111101110",
33194 => "101111101011110110000000",
33195 => "101001000111111110101110",
33196 => "100111011111001101100001",
33197 => "101010000100000100111100",
33198 => "101111000110000110010000",
33199 => "110101010101001111111111",
33200 => "111011100100000110101111",
33201 => "000001000011000001111000",
33202 => "000100101000100010110000",
33203 => "000101001010110100100111",
33204 => "000100001011001001101000",
33205 => "000011001101101011010010",
33206 => "000001111010010110000110",
33207 => "000001000011011010100001",
33208 => "000001010110011000010010",
33209 => "000001101111101110101001",
33210 => "000010010011110000100000",
33211 => "000100001010111100011100",
33212 => "000111010010110010001111",
33213 => "001010110110110101111000",
33214 => "001101110011010110101000",
33215 => "001110101111111111010100",
33216 => "001101001110111011100110",
33217 => "001010000001110110011001",
33218 => "000101101101110011010110",
33219 => "000000111011101111101001",
33220 => "111101000011111111001001",
33221 => "111010111011100111110000",
33222 => "111010001011001001011111",
33223 => "111010100111101010010111",
33224 => "111101001100001110111011",
33225 => "000001000100101011101010",
33226 => "000010011001110000011100",
33227 => "111111011111101011000011",
33228 => "111011000001110010100111",
33229 => "111000011000010000110010",
33230 => "111001001001011011111011",
33231 => "111011110011110001100110",
33232 => "111101110001010011110000",
33233 => "111111000101101110011101",
33234 => "000000111111001011100110",
33235 => "000011101100100101010011",
33236 => "000110100100111100001100",
33237 => "001000100101110011000101",
33238 => "001001100111111001011110",
33239 => "001010001011001011000100",
33240 => "001010001011010111111000",
33241 => "001000111111010111111101",
33242 => "000110010110000111010100",
33243 => "000011110000010000110000",
33244 => "000010000101000101111001",
33245 => "111111110111110111011101",
33246 => "111101100000101100101100",
33247 => "111100111110010011111100",
33248 => "111101100011100100110100",
33249 => "111101010000100101101010",
33250 => "111011110000111001100000",
33251 => "111010000011110101111101",
33252 => "111001010011010000000110",
33253 => "111010100101001110011010",
33254 => "111110010110000001101111",
33255 => "000011000100101011110101",
33256 => "000111000011101100010001",
33257 => "001011001001110001010101",
33258 => "010000001100110111111110",
33259 => "010100001101010111001100",
33260 => "010101010010011000011110",
33261 => "010100000001010101110110",
33262 => "010001110101111101111010",
33263 => "001111110001100110000110",
33264 => "001101100100001011010100",
33265 => "001001111010000001010101",
33266 => "000101000101110011000001",
33267 => "000000011111100010110111",
33268 => "111100011010011101001010",
33269 => "111001001011111101010010",
33270 => "110110101110010100000000",
33271 => "110100011010101101011001",
33272 => "110011100111100100010100",
33273 => "110101010001001011110010",
33274 => "110111110100010110011111",
33275 => "111010110011110001110110",
33276 => "111110111111011011101100",
33277 => "000011111000001010001110",
33278 => "001001010101000010100101",
33279 => "001111010110111011101000",
33280 => "010011011100101101001000",
33281 => "010011001011000111110010",
33282 => "001111000001010011001010",
33283 => "000111101111101110111001",
33284 => "111101111111111000100011",
33285 => "110011000110101011100110",
33286 => "101000011111110110111110",
33287 => "100001111010100101101101",
33288 => "100001010000010110011011",
33289 => "100001110110100110101011",
33290 => "100001011001010100000101",
33291 => "100001111011111111110101",
33292 => "100010100001011001111001",
33293 => "100011111001010011101111",
33294 => "101001011111010111101000",
33295 => "110001011110111000110110",
33296 => "111000011101010100011100",
33297 => "111101101011100100010011",
33298 => "000000000011001110011010",
33299 => "111111110101011110101111",
33300 => "111110111111011010111100",
33301 => "111101111110101111100010",
33302 => "111101011001101111101100",
33303 => "111110001100010100100011",
33304 => "111111010100011110111110",
33305 => "111111101000001111110110",
33306 => "111110111110011011101101",
33307 => "111101001111100011011000",
33308 => "111011101010010011001100",
33309 => "111100000010110010010011",
33310 => "111101011011111000010101",
33311 => "111101100001010001011010",
33312 => "111100010010101011000110",
33313 => "111011000001110110010100",
33314 => "111010010111111000011111",
33315 => "111011011010101110111101",
33316 => "111110101110000010010000",
33317 => "000010111000001001000110",
33318 => "000111010101100000000100",
33319 => "001100010110111101001110",
33320 => "010000101110011010111010",
33321 => "010011101101101010111100",
33322 => "010101000000000110001010",
33323 => "010100000000001010111010",
33324 => "010010100001101001101010",
33325 => "010001100100011010000100",
33326 => "001110111001000010010010",
33327 => "001010101011111000101100",
33328 => "000111011010101110100010",
33329 => "000101000011110000001101",
33330 => "000010110111111111010000",
33331 => "000001100101010011000111",
33332 => "000001011101110100010011",
33333 => "000001101111100001111100",
33334 => "000010010111101010110011",
33335 => "000011111010010011110110",
33336 => "000101001110101111101010",
33337 => "000100100101110101100010",
33338 => "000010001111000100010111",
33339 => "111111100100110010001111",
33340 => "111101110001101000101001",
33341 => "111100111100001001101001",
33342 => "111100011011111111000010",
33343 => "111100100001001110011010",
33344 => "111100011010001111100101",
33345 => "111001000000010001100110",
33346 => "110001110001100011001100",
33347 => "101010101011000110101100",
33348 => "100111000101111001100011",
33349 => "100110110010010001101100",
33350 => "101000001110100111000010",
33351 => "101011101010110001101100",
33352 => "110001101000001000001100",
33353 => "110111110110110000000100",
33354 => "111011101001011000111110",
33355 => "111101000011100011100011",
33356 => "111101010100101001110111",
33357 => "111100110100011011100111",
33358 => "111011010010010100101100",
33359 => "111001000101110001101111",
33360 => "110111010101100000000100",
33361 => "110110010100100011001101",
33362 => "110101111010111011000100",
33363 => "110110011111000010110011",
33364 => "111000011111010100101110",
33365 => "111101011101101000011100",
33366 => "000101110000110110100111",
33367 => "001101011000111010100100",
33368 => "010001000001000011111010",
33369 => "010010000110001111011000",
33370 => "010010001010111010111000",
33371 => "010000001000110011000100",
33372 => "001011011000100100101111",
33373 => "000101111110000001010011",
33374 => "000010011111111000000101",
33375 => "000000110111101010000000",
33376 => "111111100000111001101100",
33377 => "111110100001010010111110",
33378 => "111110111111101010111111",
33379 => "000000111101000011101100",
33380 => "000011001111000110001001",
33381 => "000101001111010010110110",
33382 => "000111111010001001110101",
33383 => "001100000101001111110110",
33384 => "010001000000110101011100",
33385 => "010100111101111011011100",
33386 => "010110100110110110100000",
33387 => "010101110010011011101000",
33388 => "010011000011110010011010",
33389 => "001111101100101010000010",
33390 => "001101010010010000111000",
33391 => "001011010100110110111110",
33392 => "001000011110000111110001",
33393 => "000101011100110000101110",
33394 => "000010111101000001001111",
33395 => "000000011101111110101001",
33396 => "111101110101100010001110",
33397 => "111010011001010011011100",
33398 => "110110001110101111000110",
33399 => "110011011101001101001110",
33400 => "110010000001010011110000",
33401 => "110000000011111011100010",
33402 => "101110100101111001100110",
33403 => "101110111000100101100110",
33404 => "101111111100000110010110",
33405 => "110001110111000101011100",
33406 => "110101110001001010111001",
33407 => "111011011000111100010111",
33408 => "000001101100001001011111",
33409 => "000111101111010111000011",
33410 => "001100110110001001001000",
33411 => "010000011000100101010010",
33412 => "010001110011000011010000",
33413 => "010000111011001101000010",
33414 => "001101100110101001011000",
33415 => "000111111100001111001110",
33416 => "000000110110101010110100",
33417 => "111010000010111000100010",
33418 => "110101100011011111101010",
33419 => "110011011101010111001010",
33420 => "110010001100110101010100",
33421 => "110001101111111111001000",
33422 => "110010101110000010011000",
33423 => "110101010010100101011001",
33424 => "111001100111010101010010",
33425 => "111110001011010101110001",
33426 => "000001010100000010000110",
33427 => "000100001010110100010100",
33428 => "001000100010001110010100",
33429 => "001101100011111000010100",
33430 => "010001001101010010111000",
33431 => "010011110110111110011010",
33432 => "010110100110111101000010",
33433 => "011000001111000101101111",
33434 => "010111011101011011100100",
33435 => "010011101001001001101010",
33436 => "001100101111000001001110",
33437 => "000100101100011101000101",
33438 => "111100011010101000000010",
33439 => "110011100111100110111110",
33440 => "101011101110001001111110",
33441 => "100101011100110111001000",
33442 => "100001101000111100011101",
33443 => "100001100011110011100110",
33444 => "100010101010101101000101",
33445 => "100011110011100101111011",
33446 => "101000101100000111100110",
33447 => "110001001111101110101010",
33448 => "111001100101011110010011",
33449 => "000000101011001100000100",
33450 => "000110001100011111111010",
33451 => "001001000111100011001000",
33452 => "001010010111110011111000",
33453 => "001011000001101110100100",
33454 => "001001101100000111000110",
33455 => "000101001111111010011011",
33456 => "000000011100100001010101",
33457 => "111110010101111001000110",
33458 => "111101001110100100011011",
33459 => "111010111110000100110111",
33460 => "111001001110100001010110",
33461 => "111000111011100100001100",
33462 => "111001010101000010010000",
33463 => "111010110101001011011110",
33464 => "111100110101010000010010",
33465 => "111101101101011011101011",
33466 => "111101110010011110110111",
33467 => "111101100000101000100011",
33468 => "111100100011111100100011",
33469 => "111100100001000100000011",
33470 => "111111010000000101101010",
33471 => "000011011111001101100111",
33472 => "000110111000101100001111",
33473 => "001001111100110100111100",
33474 => "001110000101000001100000",
33475 => "010010000100101010011110",
33476 => "010100010011000111101110",
33477 => "010100110110000010100110",
33478 => "010100100100001000100110",
33479 => "010100101100111101101110",
33480 => "010100101011001010110000",
33481 => "010010010001010000110000",
33482 => "001110011011010110000110",
33483 => "001011001111001001000000",
33484 => "001000010011011110000101",
33485 => "000101100001100100111111",
33486 => "000010110011001100000010",
33487 => "111111111000100001111000",
33488 => "111110100110101100110010",
33489 => "111110010100111110110010",
33490 => "111011011000000001101100",
33491 => "110110110011110100010100",
33492 => "110101000100010101010110",
33493 => "110101111111001101001100",
33494 => "110110100100001011001100",
33495 => "110111011111111001001011",
33496 => "111010010001111000100110",
33497 => "111011110110110001100110",
33498 => "111001010100100110100010",
33499 => "110100000100111101010000",
33500 => "101111000000000101011010",
33501 => "101100101110010111111010",
33502 => "101101100010111111010000",
33503 => "101111011111001100000110",
33504 => "110010011110010000010000",
33505 => "110110101001000101111111",
33506 => "111010000010101111100000",
33507 => "111011110100101011110000",
33508 => "111100000111010001011010",
33509 => "111010111100010011000111",
33510 => "111001001101101101110110",
33511 => "110111010011010100101010",
33512 => "110101000100100000110100",
33513 => "110010111101000011111010",
33514 => "110000101101000100100100",
33515 => "101110011101011101001010",
33516 => "101110000011000100011110",
33517 => "110000100101001001100000",
33518 => "110101011111111011001111",
33519 => "111011110101001010011110",
33520 => "000010100001100101101111",
33521 => "001000010101101111000100",
33522 => "001011101100101001010111",
33523 => "001011111111110011010110",
33524 => "001010110101111110010111",
33525 => "001001101000100010010000",
33526 => "000111111010001001001101",
33527 => "000101000001000000010100",
33528 => "000001001101010011110111",
33529 => "111101100010100101000010",
33530 => "111010101111011111101000",
33531 => "111000010000000010101010",
33532 => "110101011100000111011100",
33533 => "110011110001001100011010",
33534 => "110110001101101110011010",
33535 => "111100100101001110100100",
33536 => "000011011101010001101111",
33537 => "001010001110110001111110",
33538 => "010001100110111110100100",
33539 => "010111010111111111011100",
33540 => "011001101100000101111011",
33541 => "011001001111010011101011",
33542 => "010111100111111110111110",
33543 => "010101100011010100010000",
33544 => "010001111111111111000010",
33545 => "001100110011110011101100",
33546 => "000111100010001011111000",
33547 => "000011010111101111001100",
33548 => "000000111100111001100101",
33549 => "000000001010100001001001",
33550 => "000000011110001101011111",
33551 => "000001110111000100100010",
33552 => "000100010011001010011111",
33553 => "000111010001010110110100",
33554 => "001001000111000010100100",
33555 => "000111110101101101110110",
33556 => "000100001001000001101110",
33557 => "000001000000110011001000",
33558 => "000000010011100000010110",
33559 => "000001101011010000011101",
33560 => "000100001100001111001101",
33561 => "000110100010010101011111",
33562 => "000111101010011110010001",
33563 => "001000111111101111111010",
33564 => "001011011011111111101010",
33565 => "001100001110000000101100",
33566 => "001001010110011000101010",
33567 => "000100001000100010001110",
33568 => "111110010000001001010100",
33569 => "111000000101011110101000",
33570 => "110001110101010001110110",
33571 => "101101001111101011101110",
33572 => "101011101001111111110000",
33573 => "101011110100001010111000",
33574 => "101100100101001101100010",
33575 => "101110100100001000000010",
33576 => "110010011100010101000010",
33577 => "110111011101101001101001",
33578 => "111100001001110000001010",
33579 => "000000010000010000010101",
33580 => "000011101010111001000011",
33581 => "000110000110100100010010",
33582 => "001000110110110011000100",
33583 => "001100010111011010011000",
33584 => "001110100110111010111010",
33585 => "001110001000010101110100",
33586 => "001011011101101101000000",
33587 => "001000100100001000111111",
33588 => "000110011000010110011111",
33589 => "000010111111110101011011",
33590 => "111101001000000111010011",
33591 => "110110010001111111110100",
33592 => "110000011001000100001110",
33593 => "101100011110011011000000",
33594 => "101001111010000110100100",
33595 => "100111000101000111011001",
33596 => "100100011100001000010101",
33597 => "100100011001110110010001",
33598 => "101000001010111001110110",
33599 => "101101110011101011111100",
33600 => "110010010110100101110010",
33601 => "110110100111111011110101",
33602 => "111101000101111000110101",
33603 => "000011110010111001001111",
33604 => "000111111000010001001100",
33605 => "001010100000010110100010",
33606 => "001101000011101101111100",
33607 => "001110000111100111011110",
33608 => "001100000111100101010000",
33609 => "000111111101110101101010",
33610 => "000011101001101011100001",
33611 => "000000010010101011010010",
33612 => "111110010110111111100100",
33613 => "111101001100000101001101",
33614 => "111100101001111001110111",
33615 => "111101110010000011010101",
33616 => "111110110110100010011110",
33617 => "111110111001000000000101",
33618 => "000000101011001010101101",
33619 => "000011011010110101110001",
33620 => "000100000001011101110111",
33621 => "000011110100100111101001",
33622 => "000100100110101001110101",
33623 => "000101001111100010001110",
33624 => "000101000001011101110011",
33625 => "000100101011111010000100",
33626 => "000100110010101000101011",
33627 => "000101111010100110000111",
33628 => "001000010011011001111011",
33629 => "001001111101000100110111",
33630 => "001001111000111011100010",
33631 => "001010011011100110000110",
33632 => "001100000110011111110000",
33633 => "001100111110111000101000",
33634 => "001011110111011101010110",
33635 => "001000101001110111110100",
33636 => "000101101010100000011110",
33637 => "000101000010001001000100",
33638 => "000100010111111110001010",
33639 => "000001000000011110000010",
33640 => "111100111101111111000010",
33641 => "111010101101010111111111",
33642 => "111000100010111000111110",
33643 => "110101001110010000010101",
33644 => "110010101111011001101110",
33645 => "110010001100101000111000",
33646 => "110011100110111100001110",
33647 => "110110111001010101000110",
33648 => "111010110100101001010100",
33649 => "111110011110101111101101",
33650 => "000000101011101110000001",
33651 => "000000001001000001000111",
33652 => "111110001010101011011110",
33653 => "111100010000000001001010",
33654 => "111010001101111110110011",
33655 => "111000001111010101111011",
33656 => "110110111001110101110100",
33657 => "110110010101111001100001",
33658 => "110110000000010100010111",
33659 => "110101100000100110111111",
33660 => "110101001001110000100011",
33661 => "110101100101101000100010",
33662 => "110111101111011111101100",
33663 => "111010110001001000001110",
33664 => "111100111100000111111001",
33665 => "111110110101110000000100",
33666 => "000000001111100011010100",
33667 => "111111110100101101010101",
33668 => "111110111001000011101011",
33669 => "111110001100001101001000",
33670 => "111101101101000110011011",
33671 => "000000000000000010111010",
33672 => "000101001001110000100000",
33673 => "001001001010010111010000",
33674 => "001010110001011001110110",
33675 => "001011110001101011011010",
33676 => "001100000110100011011110",
33677 => "001001111110000100010010",
33678 => "000110000111010011111010",
33679 => "000100000101000000101010",
33680 => "000100100101010111110111",
33681 => "000100100111000011101111",
33682 => "000010111000100001011110",
33683 => "000000100000011010011110",
33684 => "111101110010101101100101",
33685 => "111010001111001011101111",
33686 => "110110101101010010100100",
33687 => "110101111011111100000001",
33688 => "111001000010101110011011",
33689 => "111110000000110010001001",
33690 => "000011000001010110010111",
33691 => "000111110000101101011010",
33692 => "001100001000101111011100",
33693 => "001111001011000100001010",
33694 => "001111110000100111000000",
33695 => "001110101001100110010000",
33696 => "001100111010100001110010",
33697 => "001010101001000101011100",
33698 => "001000010100000100010110",
33699 => "000101101000101110100001",
33700 => "000010000100010110001001",
33701 => "111111001101100110100000",
33702 => "111110011100011001010010",
33703 => "111110101011101000000011",
33704 => "111111001011001010010011",
33705 => "000001000111101011000001",
33706 => "000100001000000011100101",
33707 => "000101110011000101111111",
33708 => "000101111100110101011111",
33709 => "000101010000011000111100",
33710 => "000011100110110100001001",
33711 => "000010100100111010011111",
33712 => "000011011010111111001101",
33713 => "000101001011101100100001",
33714 => "000110111010100101110100",
33715 => "001000011001100010010011",
33716 => "001001001100000000010100",
33717 => "001000100111001001101000",
33718 => "000111101101111110001100",
33719 => "000111110011100101001110",
33720 => "000111101111011100100101",
33721 => "000111000100110101000101",
33722 => "000101111000001001000110",
33723 => "000011100100111000111010",
33724 => "000010001000011001110101",
33725 => "000010010110000111000011",
33726 => "000010001000000001001001",
33727 => "000001101011001110101011",
33728 => "000001110100010111100010",
33729 => "000001110000010001100010",
33730 => "000001010100111000101101",
33731 => "000000110101000000111001",
33732 => "000000001000001111000011",
33733 => "111111101011100110010110",
33734 => "000000110101111100100111",
33735 => "000010010001111110000111",
33736 => "000000110110101001001100",
33737 => "111110000001101011001110",
33738 => "111100001011011111011000",
33739 => "111010011111011110001000",
33740 => "111001100010110010101001",
33741 => "111001101100111111110100",
33742 => "111001101101010111010111",
33743 => "111010010101111111011100",
33744 => "111100000011110001001110",
33745 => "111101011101101110000101",
33746 => "111101101101000010100110",
33747 => "111100110001010100101011",
33748 => "111011101001001100000101",
33749 => "111010011101101111101000",
33750 => "110111001110001111100010",
33751 => "110001001011111110011110",
33752 => "101010011000000011110100",
33753 => "100101010011111111011101",
33754 => "100011001001001101010001",
33755 => "100010111000110111111000",
33756 => "100011110011001111100110",
33757 => "100111000111001111001101",
33758 => "101100100011001101111010",
33759 => "110001110010011100000100",
33760 => "110110010001101001000100",
33761 => "111010100110000001110110",
33762 => "111110101100110001101010",
33763 => "000010100000010110010010",
33764 => "000101010100111110100000",
33765 => "000110100000110001000100",
33766 => "000111000101110110111010",
33767 => "001000100011101011001101",
33768 => "001010011000101001001010",
33769 => "001011001000111011110000",
33770 => "001011010011011001000010",
33771 => "001011000100101101100111",
33772 => "001001001100110110000110",
33773 => "000110110110001011111001",
33774 => "000101110011000100111001",
33775 => "000100101011100111000101",
33776 => "000001110011100111110010",
33777 => "111101111011101000100000",
33778 => "111011011001000011001101",
33779 => "111011101111011101001000",
33780 => "111110000110110010010111",
33781 => "000000110010000010100111",
33782 => "000100010010010111100001",
33783 => "001010000111100001100010",
33784 => "010000010001011011011100",
33785 => "010100010001101010100110",
33786 => "010111100111001000111010",
33787 => "011010101011011000110111",
33788 => "011011111011110000011001",
33789 => "011011001000111110100001",
33790 => "010111011001010110000100",
33791 => "010001011011111010100110",
33792 => "001100000010010101111000",
33793 => "000110100010111111010001",
33794 => "111111011000010100011001",
33795 => "111000010101011010011111",
33796 => "110011100111000100010100",
33797 => "110000011011000001001010",
33798 => "101101010101000110011110",
33799 => "101011010100111100110100",
33800 => "101011010000000110110000",
33801 => "101101001100001110110010",
33802 => "110001001101001000110100",
33803 => "110100111000100010110010",
33804 => "110110101010101010110001",
33805 => "110111001111110111100100",
33806 => "110110010010011101100001",
33807 => "110100111010000101110000",
33808 => "110100100011001000011010",
33809 => "110100010000011010101001",
33810 => "110011101110001011100000",
33811 => "110010111111111010101010",
33812 => "110010010010010010110010",
33813 => "110010001101101000000010",
33814 => "110001111100111000010110",
33815 => "110001110001111111011010",
33816 => "110011011111011110111000",
33817 => "110110111000000111100110",
33818 => "111010001000010101101010",
33819 => "111100000111000001000010",
33820 => "111101111100010011110101",
33821 => "000000011010001110000110",
33822 => "000001001111111111110111",
33823 => "111111111011000010100000",
33824 => "111111001100101100010000",
33825 => "000000011001100101000010",
33826 => "000010011100011111110100",
33827 => "000011010111111100100111",
33828 => "000010001010101100100101",
33829 => "000000010111010110000101",
33830 => "111111010110011010011011",
33831 => "111110101001000011101011",
33832 => "111110110001111011000010",
33833 => "000001000100000101001010",
33834 => "000101000100111100011001",
33835 => "001001000110111000010001",
33836 => "001010110111010110101100",
33837 => "001001011001110000110110",
33838 => "000110000001000110010100",
33839 => "000001100010010111001111",
33840 => "111101000010000101111010",
33841 => "111010110111111111011010",
33842 => "111011110000010001110100",
33843 => "111110100101010101001100",
33844 => "000001111110010111000101",
33845 => "000100110000011000010111",
33846 => "000110100000000100110000",
33847 => "000110111111111101111001",
33848 => "000110011111011011010001",
33849 => "000101001011111011000101",
33850 => "000011000100100111100010",
33851 => "000001000111000001101110",
33852 => "111111010111000010001110",
33853 => "111101001110000011011011",
33854 => "111011011001000111101000",
33855 => "111001111000000100100011",
33856 => "111000110000100100100100",
33857 => "111001010011100000111111",
33858 => "111011010110101101010000",
33859 => "111101101111000101100111",
33860 => "111111011110011000001001",
33861 => "111111101010000001110000",
33862 => "111110001000111000000000",
33863 => "111011110000010101010000",
33864 => "111001011110101101011111",
33865 => "110111110000010100010100",
33866 => "110111111001110011111010",
33867 => "111011000100001001100110",
33868 => "111111000010001010011000",
33869 => "000010001000001110100011",
33870 => "000101100100000011011011",
33871 => "001000110010111001000111",
33872 => "001010000010001011011100",
33873 => "001001100011100000110100",
33874 => "001000110110101010011100",
33875 => "001000110100001111010001",
33876 => "001000111101111000100000",
33877 => "001000101101110010010011",
33878 => "001000001101111000010010",
33879 => "000111110101010001000110",
33880 => "000111100111101110101110",
33881 => "000110101011110110101000",
33882 => "000101000011000011111001",
33883 => "000100001001110100101100",
33884 => "000100000000001011100100",
33885 => "000100011100011111000100",
33886 => "000101110000011101110110",
33887 => "000110111001111000111110",
33888 => "001000101000011001000001",
33889 => "001100011011000011001100",
33890 => "010000100001000000011110",
33891 => "010011101111100010000010",
33892 => "010110110100111000001000",
33893 => "011001000101001011010101",
33894 => "011001101101010010111001",
33895 => "011000101011000011101011",
33896 => "010110000000010111001110",
33897 => "010010100111100000101010",
33898 => "001111111100110001001110",
33899 => "001101111001110110110010",
33900 => "001010011000011110001011",
33901 => "000101011001101010011001",
33902 => "000000111011101001000101",
33903 => "111100010010010100000010",
33904 => "110111010100000001000101",
33905 => "110001110110101101101010",
33906 => "101001100010001110001110",
33907 => "100010010110000110101101",
33908 => "100001010011110100110011",
33909 => "100010010111000100111000",
33910 => "100010100011000101110101",
33911 => "100011100010111011101011",
33912 => "100110011110011101001011",
33913 => "101100101101111101000000",
33914 => "110101001000000010100010",
33915 => "111101100000111001011010",
33916 => "000101011111011111111110",
33917 => "001011100100100001110100",
33918 => "001111000110000010110100",
33919 => "010000100001101010110110",
33920 => "010000000101000001000010",
33921 => "001110101101010100100010",
33922 => "001100011111011111001100",
33923 => "001001011001010100001100",
33924 => "000101000111111110111000",
33925 => "111111100101011010011000",
33926 => "111011000100110001000100",
33927 => "110111110011110001000010",
33928 => "110100111110100000000110",
33929 => "110011010001001010010110",
33930 => "110001011110111100100010",
33931 => "110000110011000100011110",
33932 => "110011010000001111110100",
33933 => "110110110101101111110111",
33934 => "111011100101011010011001",
33935 => "000010010001110011101001",
33936 => "001001000011000011100110",
33937 => "001110101110000110000000",
33938 => "010011000111000101010110",
33939 => "010111010111001000010110",
33940 => "011011001000111111000001",
33941 => "011100001011101011001110",
33942 => "011011011011111011100111",
33943 => "011001111001111000100010",
33944 => "010110011110011110011000",
33945 => "010000101010010101000000",
33946 => "001000111100111111111010",
33947 => "000010000110000000110100",
33948 => "111101101111101110110010",
33949 => "111010011110101100001100",
33950 => "110111100111101110010010",
33951 => "110101001110110000100011",
33952 => "110011111011010000101010",
33953 => "110100000101101110110000",
33954 => "110100111101110101101001",
33955 => "110110100101110111000000",
33956 => "111000101011111110000001",
33957 => "111011100011111110001001",
33958 => "111110111001001000100000",
33959 => "111110101001100111101011",
33960 => "111010110011110011100000",
33961 => "111000000100111000110010",
33962 => "110111011101010101000010",
33963 => "110111101110100101001101",
33964 => "110111100111011111100110",
33965 => "110110011001100100010011",
33966 => "110101011010111001011010",
33967 => "110100110100011111110110",
33968 => "110011100011010110110100",
33969 => "110010010100110000100100",
33970 => "110010100111100000111000",
33971 => "110100010111000000100001",
33972 => "110101100100110100011000",
33973 => "110101110110000100000110",
33974 => "110110011111001100110001",
33975 => "110110111110100000100101",
33976 => "110110010111010101010011",
33977 => "110101000000110011101111",
33978 => "110100000111101011010000",
33979 => "110101001001011101100010",
33980 => "110111010010111010101000",
33981 => "111000110001111010111101",
33982 => "111001111010001111000010",
33983 => "111010101100111110000000",
33984 => "111010101101110110111100",
33985 => "111011100010111000111001",
33986 => "111110001110011010110010",
33987 => "000010001001001100110111",
33988 => "000111000101111010111010",
33989 => "001011101100100010001100",
33990 => "001101111010011000111000",
33991 => "001101100111011101000010",
33992 => "001010101010000111100101",
33993 => "000101000000101111100110",
33994 => "111110100111111010101001",
33995 => "111001010100001011101100",
33996 => "110110000100000010001010",
33997 => "110101010000100010110000",
33998 => "110110001001011001001111",
33999 => "111000001011001100010111",
34000 => "111011010101000001001101",
34001 => "111110111101111010000011",
34002 => "000010000111100010011001",
34003 => "000101000000101001101100",
34004 => "001000011110011110000000",
34005 => "001010111101100001101001",
34006 => "001010000110011110011011",
34007 => "000110100001110110011100",
34008 => "000010011101101100111010",
34009 => "111111010111110001010010",
34010 => "111101011101110010110100",
34011 => "111100010001011010100110",
34012 => "111100001001001100110010",
34013 => "111101001100100011011111",
34014 => "111110001011010010110100",
34015 => "111110000001000010010011",
34016 => "111100010110000011101011",
34017 => "111001100100001010010100",
34018 => "110110110101110001111011",
34019 => "110100111101111000000110",
34020 => "110100101001111001010000",
34021 => "110110011111110100110000",
34022 => "111001110110000110110010",
34023 => "111101101010100100011000",
34024 => "000001000100101101110101",
34025 => "000011001000011001000010",
34026 => "000011111110100101010000",
34027 => "000100001001001000000010",
34028 => "000011100010010010000001",
34029 => "000010100000001011101000",
34030 => "000001010011101100011010",
34031 => "111111101011101101001111",
34032 => "111101110101110100111001",
34033 => "111100010000011000110001",
34034 => "111011010011101001101111",
34035 => "111010111110011010100101",
34036 => "111010111010011000110000",
34037 => "111011001011110110101011",
34038 => "111011111110001011110001",
34039 => "111101011010001100101011",
34040 => "111111010010100011110100",
34041 => "000001000001110010100001",
34042 => "000011000100100001110111",
34043 => "000110001100000100111001",
34044 => "001010000101001110100010",
34045 => "001110001000001100011110",
34046 => "010010010000110011100100",
34047 => "010110100101001111100100",
34048 => "011001110000001100101101",
34049 => "011010101001010110101011",
34050 => "011010010011101001011001",
34051 => "011000110011111000001011",
34052 => "010101100000110100111100",
34053 => "010001100110011000011110",
34054 => "001101101110101010010010",
34055 => "001001010010001101001101",
34056 => "000100000100000010011100",
34057 => "111110111011100111100100",
34058 => "111011000001011111010000",
34059 => "110111111011010010111101",
34060 => "110101000000110011101101",
34061 => "110010001011101011111010",
34062 => "101110111000010100111000",
34063 => "101100010001000111100110",
34064 => "101100101000100110100000",
34065 => "110000000000100010011010",
34066 => "110100011111101111110000",
34067 => "111000111110011001001111",
34068 => "111110011011010011100101",
34069 => "000100111110011111111000",
34070 => "001010100100001111111001",
34071 => "001110011000000010010110",
34072 => "010000100001110101110100",
34073 => "010000101000111111000110",
34074 => "001111000010001011100110",
34075 => "001011101101000100111101",
34076 => "000101110000101110010100",
34077 => "111110000001000100100111",
34078 => "110111001011110111101001",
34079 => "110010001100011101101110",
34080 => "101110010010111001100100",
34081 => "101011110100011101111000",
34082 => "101010010000100011000100",
34083 => "101001100101100110001110",
34084 => "101100001011100111111000",
34085 => "110001000101110111110000",
34086 => "110101100100011100010110",
34087 => "111001111110000101010100",
34088 => "111101111101100100011101",
34089 => "000001011101110001101011",
34090 => "000110100110010100101011",
34091 => "001100100101111000000110",
34092 => "010000111100111000001110",
34093 => "010100100111100010110010",
34094 => "011001000010111111100010",
34095 => "011011101110110010001101",
34096 => "011010011000100000110011",
34097 => "010110110110000111000000",
34098 => "010010111111100000100010",
34099 => "001110111001111010101000",
34100 => "001001010000001011100001",
34101 => "000000101101110100110101",
34102 => "111001011000110000110110",
34103 => "110111101010000101110010",
34104 => "111000001000001101100110",
34105 => "110110111111101000001110",
34106 => "110110011011000111010110",
34107 => "111001011001000100000110",
34108 => "111110001110111010100101",
34109 => "000001101001011110110101",
34110 => "000100101011010001001001",
34111 => "001000100100111100100010",
34112 => "001011000010101011001111",
34113 => "001010010101001010000000",
34114 => "000110100000010010000010",
34115 => "000010010001000101001110",
34116 => "000000001110100001110010",
34117 => "111110110000010011001011",
34118 => "111101101101000100011110",
34119 => "111110010100101110011010",
34120 => "111110011001001001111010",
34121 => "111101000010110011100101",
34122 => "111011100001110110001100",
34123 => "111010001001110100010010",
34124 => "111001010110111100011111",
34125 => "111001000101011000100101",
34126 => "111001010000010100110100",
34127 => "111010101000110100101110",
34128 => "111101010000001110111111",
34129 => "111111111110100000011010",
34130 => "000001011101100110101000",
34131 => "000010001110001011000101",
34132 => "000011100100110001100101",
34133 => "000100101101101011110111",
34134 => "000100011000000110100110",
34135 => "000010010100010011001001",
34136 => "111111011111100110100100",
34137 => "111101011001101101110001",
34138 => "111010111010110000101011",
34139 => "110111000100111011000000",
34140 => "110101010001101111111111",
34141 => "111000010011011010110000",
34142 => "111101111011101100111101",
34143 => "000010101000111110100101",
34144 => "000110010001000010100111",
34145 => "001010001010100101010000",
34146 => "001100010000100001011000",
34147 => "001001001111100110111111",
34148 => "000010010000110011010011",
34149 => "111011010010111001100001",
34150 => "110101111100010010111010",
34151 => "110001100110010000101100",
34152 => "101111000011010010111110",
34153 => "101111100100101100001010",
34154 => "110010010101101000100100",
34155 => "110110000100000011111110",
34156 => "111010001100101011100011",
34157 => "111110010100001101000110",
34158 => "000010010011110010010101",
34159 => "000101101010110000011000",
34160 => "000111000111001100011100",
34161 => "000101101010110101111111",
34162 => "000001101100101000010000",
34163 => "111101001010100000000100",
34164 => "111010001100101100010010",
34165 => "111001010101001010000001",
34166 => "111001000100000001001111",
34167 => "110111101111000000000101",
34168 => "110110010110101010111010",
34169 => "110110011110101001110000",
34170 => "110110110111011000110000",
34171 => "110110001110001100011110",
34172 => "110101011010001100111110",
34173 => "110101011110100000010001",
34174 => "110110111101010101001000",
34175 => "111001110101100100001101",
34176 => "111101010010101010001101",
34177 => "000000111011100111010010",
34178 => "000100011101111100011110",
34179 => "000110100000011010110011",
34180 => "000110101010110111101111",
34181 => "000110000110001000101010",
34182 => "000100100101100011011101",
34183 => "000001111000111010101110",
34184 => "111111100000010001010000",
34185 => "111101111001010001000010",
34186 => "111100010101010100000010",
34187 => "111011001010011011110110",
34188 => "111010110010000101010110",
34189 => "111010111100101001101100",
34190 => "111011111100011001011010",
34191 => "111101101010010000101111",
34192 => "111110111101101010100000",
34193 => "000000001111010000110101",
34194 => "000010011000100110001110",
34195 => "000011010100001100110110",
34196 => "000001101010101100101011",
34197 => "111111111011110100100111",
34198 => "000000000010110000111111",
34199 => "000001110011101111100001",
34200 => "000100011111110011101000",
34201 => "000110111101101100111011",
34202 => "001001000000110101011110",
34203 => "001010100111101110101000",
34204 => "001010110110100000010101",
34205 => "001010001100100000010100",
34206 => "001001101000111111111000",
34207 => "001000101010011110110100",
34208 => "000110111101011001111110",
34209 => "000100110011011100001010",
34210 => "000010100010101101010000",
34211 => "000000011000100010110100",
34212 => "111101101001001011010110",
34213 => "111010010000011110001100",
34214 => "110111000000000011011000",
34215 => "110100000010001011110100",
34216 => "110001100011010110000010",
34217 => "101111011110000110011100",
34218 => "101101111110100101011110",
34219 => "101110011010110010101000",
34220 => "110001001000011110111100",
34221 => "110101100110010110010111",
34222 => "111010111101101101011110",
34223 => "000000010100110101010100",
34224 => "000110100101000010110101",
34225 => "001101000110011101011010",
34226 => "010000111111000111110110",
34227 => "010010000000101001110000",
34228 => "010001100110011110111110",
34229 => "010000011001000101010100",
34230 => "001110011010101001101100",
34231 => "001011011111011011010111",
34232 => "001000000101111100010110",
34233 => "000100101100011111010101",
34234 => "000010001110001111011011",
34235 => "000000111100101100010010",
34236 => "111111101011000010001101",
34237 => "111111011100111001110101",
34238 => "000000101011110110111110",
34239 => "000001101011011110101110",
34240 => "000011010000011110001101",
34241 => "000100111110111101110110",
34242 => "000101010000010111010011",
34243 => "000101010001010010100011",
34244 => "000101010101000001011000",
34245 => "000101001100010011111110",
34246 => "000100111010000001001110",
34247 => "000011100100110110100011",
34248 => "000001110011001001100101",
34249 => "000001001010100101100111",
34250 => "000010110100001101010010",
34251 => "000101010100111101110111",
34252 => "000101100100011001110101",
34253 => "000100011011101011101100",
34254 => "000100000101000111001110",
34255 => "000100011011110010101100",
34256 => "000100011100001110110001",
34257 => "000010010101110000100110",
34258 => "111111110111111101100111",
34259 => "111111110000101100110100",
34260 => "000000000100100100111101",
34261 => "111111001001111101110001",
34262 => "111101111001000010111011",
34263 => "111101101110001011011000",
34264 => "111110010100101110001000",
34265 => "111100110110100100011000",
34266 => "111001010000111100000010",
34267 => "110101001100010010000111",
34268 => "110000111110110100111100",
34269 => "101101101011100011110000",
34270 => "101011001110001101110100",
34271 => "101010101000010101010100",
34272 => "101110100010011111101000",
34273 => "110101110001011111100010",
34274 => "111101100001010010101001",
34275 => "000011011110001000110110",
34276 => "000110100100101101111101",
34277 => "001000101101011010000101",
34278 => "001010011001111100010110",
34279 => "001010010111100100000101",
34280 => "001000100100100100010100",
34281 => "000110000001101001101001",
34282 => "000100001001111010101000",
34283 => "000010111110001110010100",
34284 => "000010000101001000100101",
34285 => "000001101010000111111001",
34286 => "000001000010001110010111",
34287 => "000000110111000110011101",
34288 => "000001110000000000011010",
34289 => "000001111111110000000010",
34290 => "000001000001110000011010",
34291 => "111111011110011011110101",
34292 => "111101100010100100111110",
34293 => "111011101100011110001110",
34294 => "111010111100101101101011",
34295 => "111100101110111010101111",
34296 => "000001001111100111111001",
34297 => "000110111000010110011011",
34298 => "001011110000110101101110",
34299 => "001110111000101010100100",
34300 => "010000010000110010011110",
34301 => "001111010111111011101110",
34302 => "001011011100100100110010",
34303 => "000100101110010001000101",
34304 => "111100011010001100000011",
34305 => "110101000101101101101110",
34306 => "110000001110010101101010",
34307 => "101100111100111110110000",
34308 => "101011000011010111001010",
34309 => "101010101110000101010000",
34310 => "101100001001010111111000",
34311 => "101111100110001000100110",
34312 => "110011110110100101000000",
34313 => "110111111011111000111010",
34314 => "111100000101110110111011",
34315 => "111111101110110101111010",
34316 => "000001001111110110000100",
34317 => "000000001111110110000011",
34318 => "111110111101010100100001",
34319 => "111110100000110011110110",
34320 => "111101010001110101001101",
34321 => "111011010001001111101000",
34322 => "111001010111011101010100",
34323 => "110111000110011101010110",
34324 => "110101000010011100111110",
34325 => "110011011100010111101010",
34326 => "110001101010110010010100",
34327 => "110001000110101110111000",
34328 => "110011001000000110010010",
34329 => "110110111101100111110010",
34330 => "111011111110001100000101",
34331 => "000010001000111001010110",
34332 => "001000100111110100101111",
34333 => "001101100000001110101110",
34334 => "001111101000010100110000",
34335 => "001111100111101000111010",
34336 => "001110001111000100111000",
34337 => "001011111101011111001100",
34338 => "001000010111000010001000",
34339 => "000010110111001000111010",
34340 => "111110101010000010011000",
34341 => "111110100101000000000001",
34342 => "000000000010101101100011",
34343 => "000000111110111000101011",
34344 => "000010010110000000011000",
34345 => "000100101001100001101010",
34346 => "000111010001010110111110",
34347 => "001000100011001010011110",
34348 => "000111110101101011000001",
34349 => "000110100010000111110000",
34350 => "000110001100001000001110",
34351 => "000110111000101110011011",
34352 => "000111001001101000111001",
34353 => "000111011011100000011000",
34354 => "001001010111100111010101",
34355 => "001100011101011000010100",
34356 => "001111101011001011111100",
34357 => "010000101100000110000010",
34358 => "001110010111110011001010",
34359 => "001011111100010101001010",
34360 => "001010010011110110001001",
34361 => "001000001001111010001100",
34362 => "000101100100111100110111",
34363 => "000010011000101001010100",
34364 => "000000000110110100011001",
34365 => "111111110010011101010111",
34366 => "111111110011111101010001",
34367 => "111111000001111010001000",
34368 => "111100010101111110101111",
34369 => "111000101100111010110110",
34370 => "110101011010101100001011",
34371 => "110000100101010011111100",
34372 => "101011001000011100010100",
34373 => "100111110010010100111001",
34374 => "100110001110100011011011",
34375 => "100110001100100111111111",
34376 => "100111111100101011011001",
34377 => "101011110101100100011010",
34378 => "110001100100011000111000",
34379 => "110111111010011001110010",
34380 => "111110111110011110101000",
34381 => "000100111111111000101100",
34382 => "000111101111110111001010",
34383 => "001001001110000000010100",
34384 => "001001101110110010111001",
34385 => "000111011001001000011110",
34386 => "000100000101101111001100",
34387 => "000010000100000000001011",
34388 => "000000110000011101000110",
34389 => "111111111110000011111110",
34390 => "000000011100011011101000",
34391 => "000010000110000000010100",
34392 => "000100001010101111001100",
34393 => "000110000110011101011011",
34394 => "000111011111110000010100",
34395 => "001000100100010100010111",
34396 => "001001111010000010111000",
34397 => "001010010100101000110100",
34398 => "001000011000011110010110",
34399 => "000110100011010111101110",
34400 => "000110110010101011000100",
34401 => "000110110110010000000101",
34402 => "000111010101110000110110",
34403 => "001010010111001111010010",
34404 => "001101101110111101011000",
34405 => "010001000000000110000110",
34406 => "010100111000000100100110",
34407 => "010110110111110100110000",
34408 => "010110111111011011101110",
34409 => "010111100000100011001100",
34410 => "010111100111100000010010",
34411 => "010100111110011001111110",
34412 => "010000000100011101100000",
34413 => "001011001001001100001000",
34414 => "000110010101110000001011",
34415 => "000010100010010010101001",
34416 => "000000001000000100011010",
34417 => "111011110111011011010100",
34418 => "110101110011010010011110",
34419 => "101111111111100011111010",
34420 => "101010110111001111100000",
34421 => "100111110000010111011101",
34422 => "100100111110000011100000",
34423 => "100001110101101101101111",
34424 => "100001011001001101000011",
34425 => "100011000100110011001110",
34426 => "100111001111001111010101",
34427 => "101110110011101011111010",
34428 => "110111100011011100101100",
34429 => "000001100100000111000000",
34430 => "001010110111110010001010",
34431 => "001111101001011100011010",
34432 => "010000101010110010110100",
34433 => "001111110110010110011010",
34434 => "001110011111110001100000",
34435 => "001010011111110011110000",
34436 => "000001100000110011010110",
34437 => "111000111010100111011010",
34438 => "110100100001011010011001",
34439 => "110001111000100111011000",
34440 => "101111010111100011010010",
34441 => "101101010011000111111010",
34442 => "101110110010100111010110",
34443 => "110101010000101010001110",
34444 => "111100000101011110011111",
34445 => "111111101101001111011000",
34446 => "000001000111111100011100",
34447 => "000010010101100001011110",
34448 => "000011101101110101000101",
34449 => "000100111101110100111100",
34450 => "000110111001000111000100",
34451 => "001010000101011000010100",
34452 => "001110100010010101011010",
34453 => "010010011000101111010100",
34454 => "010011000001110011100100",
34455 => "010001111100110110010100",
34456 => "010000010010110011101000",
34457 => "001011100100100001101100",
34458 => "000011110101010110001111",
34459 => "111011111100111101011000",
34460 => "110101110111101010011110",
34461 => "110001110110111101010010",
34462 => "101111010100101100001110",
34463 => "101110001000111011000100",
34464 => "101110010010111011101100",
34465 => "101111101000100011010100",
34466 => "110001111100111000011010",
34467 => "110101101100010100111101",
34468 => "111011100000100100001011",
34469 => "000000110000101010000000",
34470 => "000010110010010100100101",
34471 => "000011011000001000110111",
34472 => "000011101110101111111001",
34473 => "000011000000110000011011",
34474 => "000001001010001010000101",
34475 => "111101111100101011111101",
34476 => "111010000000000100001000",
34477 => "110110101111011100100110",
34478 => "110011111111110010111100",
34479 => "110001010010001011001010",
34480 => "101110111101001010011100",
34481 => "101101001011001100010000",
34482 => "101100001000111100011000",
34483 => "101101000110010001111110",
34484 => "110001010000100001010010",
34485 => "110111010000111011111110",
34486 => "111101000001111011111101",
34487 => "000010101001111000110010",
34488 => "000111011011111010100011",
34489 => "001001011010010110111000",
34490 => "001000111100000100011110",
34491 => "000110111010011001001101",
34492 => "000011111110110011100000",
34493 => "000001111000001101100111",
34494 => "000000001101011011010100",
34495 => "111101110011100101000000",
34496 => "111100011100010100100111",
34497 => "111101011100000101100001",
34498 => "111111110111000100110101",
34499 => "000010100000111111010111",
34500 => "000100110110101111100001",
34501 => "000111011010111011010010",
34502 => "001010001101010100100100",
34503 => "001011100110001001100001",
34504 => "001010011111101110001000",
34505 => "001000011000111001101111",
34506 => "000111011111100011110000",
34507 => "000110111101111000111001",
34508 => "000101011000001111001000",
34509 => "000011111101111010111001",
34510 => "000011011011010010001001",
34511 => "000011100111110111110010",
34512 => "000100101000001100110011",
34513 => "000101000101111111110011",
34514 => "000100111010001000100101",
34515 => "000101100101001000111000",
34516 => "000110011101110010000011",
34517 => "000110010111101111111001",
34518 => "000101100100110111010001",
34519 => "000100011011100110111111",
34520 => "000011100100000111100000",
34521 => "000011011001101001100000",
34522 => "000010111001000111010100",
34523 => "000001000100010111111001",
34524 => "111110001100001100001010",
34525 => "111010111000011010011100",
34526 => "110110111111111111100111",
34527 => "110001111010010011111100",
34528 => "101100100001001001011110",
34529 => "101000000011111111010100",
34530 => "100101000010111010111010",
34531 => "100100100111001111010111",
34532 => "100101011111101011110101",
34533 => "100110011110110001000111",
34534 => "101010011110101110100110",
34535 => "110000101011010101101000",
34536 => "110110001000100101111100",
34537 => "111011111011001100100111",
34538 => "000000111110011101001011",
34539 => "000100011000000100000100",
34540 => "000111011001001011010101",
34541 => "001000010001010010111011",
34542 => "000111010000001011010001",
34543 => "000110001010001010000110",
34544 => "000011111111001000111100",
34545 => "000001010000001111011110",
34546 => "111111011100100001000010",
34547 => "111110110001010110010011",
34548 => "111110101111110110110000",
34549 => "111111001010011110110001",
34550 => "000000011001111001000110",
34551 => "000000111010000111011100",
34552 => "000001000010000000101001",
34553 => "000010101011111110110111",
34554 => "000011001111101000001110",
34555 => "000010101000110001111001",
34556 => "000011110000111001111011",
34557 => "000110001011100010100111",
34558 => "001010011110110110010110",
34559 => "001111111101111101001110",
34560 => "010100100001110110101100",
34561 => "011001101001010100100111",
34562 => "011101110110010100000101",
34563 => "011110100110000101111000",
34564 => "011110001101011000110011",
34565 => "011101101001111101100001",
34566 => "011100100100010111000001",
34567 => "011011001111000100111011",
34568 => "010111000111101101101000",
34569 => "001111010101011001001110",
34570 => "000111110101000110111001",
34571 => "000011010011110100110111",
34572 => "000001000101011001110001",
34573 => "111111101011011100011001",
34574 => "111110011001100101011011",
34575 => "111101111101111001111000",
34576 => "111101100111011000011001",
34577 => "111011010011101111011011",
34578 => "111000011110110000000110",
34579 => "110111010000011010111110",
34580 => "111000000110101001110010",
34581 => "111011111011001001001100",
34582 => "000001011110100100111010",
34583 => "000110110011000011111010",
34584 => "001011110000100111011101",
34585 => "001111101111011111001110",
34586 => "010010100000000101100100",
34587 => "010011000010111000101110",
34588 => "001111001101100011001010",
34589 => "000111011011110010010111",
34590 => "111101110001011110110101",
34591 => "110101001111111000101100",
34592 => "110000000110110110011010",
34593 => "101100110100100000111010",
34594 => "101010011010011101100000",
34595 => "101010001101101001111100",
34596 => "101101011101100010001010",
34597 => "110100011111000011110110",
34598 => "111100100110100110101110",
34599 => "000010100110001010010011",
34600 => "000110010010110011101001",
34601 => "001000000111110000010000",
34602 => "000111101010010000100011",
34603 => "000101100011101101101110",
34604 => "000100000110110000000011",
34605 => "000100001101001001000010",
34606 => "000100000000010111101010",
34607 => "000010010110000001100000",
34608 => "111111111110000110100011",
34609 => "111101100010100111000011",
34610 => "111010011010110100101111",
34611 => "110101111111011000101101",
34612 => "110001101111000000001000",
34613 => "101111110000010010101000",
34614 => "110000110000001101000100",
34615 => "110011011000011011000100",
34616 => "110101000010000100010001",
34617 => "110101101111010000110000",
34618 => "110111110110100111000101",
34619 => "111011010110101000110110",
34620 => "111110001010110000011110",
34621 => "111111111010110010010000",
34622 => "000010000001100101001001",
34623 => "000100010000111111001110",
34624 => "000100100100011110010001",
34625 => "000010001001011000110111",
34626 => "111110110000011000000111",
34627 => "111101010100000011010110",
34628 => "111101101100100001100011",
34629 => "111100110111000011101001",
34630 => "111010011001111110001000",
34631 => "111000001111011000111110",
34632 => "110111010011100110011010",
34633 => "110111000111101101001100",
34634 => "110110011010001100110000",
34635 => "110101001001100000110000",
34636 => "110100110100001100000000",
34637 => "110111001101010010001000",
34638 => "111100100000011111010000",
34639 => "000010100000001111110011",
34640 => "001000100100110100001010",
34641 => "001110110010100000010010",
34642 => "010010110000010101001000",
34643 => "010011010101001101100010",
34644 => "010000111011001010110000",
34645 => "001011100110110100011100",
34646 => "000100011100100100000110",
34647 => "111101000000100101101110",
34648 => "110110110011000010011100",
34649 => "110010011100000111000110",
34650 => "101111110010110000111100",
34651 => "101111010101001010001000",
34652 => "110000111000000010101100",
34653 => "110100000110101000001010",
34654 => "111000110010100100111100",
34655 => "111101100100101000000110",
34656 => "000001111100010000110100",
34657 => "000101100010011010011000",
34658 => "000111001100101010101111",
34659 => "000111000111100011100110",
34660 => "000101110011111001111111",
34661 => "000011101101000000000111",
34662 => "000001101100001000100101",
34663 => "000000000000000101111101",
34664 => "111110101010111010101110",
34665 => "111101100100011011110110",
34666 => "111100110111101100011100",
34667 => "111101010000010000011010",
34668 => "111110001011001100100011",
34669 => "111111100110110001101000",
34670 => "000010010000010111100110",
34671 => "000100110000010001101001",
34672 => "000110010010011011000110",
34673 => "000111110101100011111000",
34674 => "001001000000101111010000",
34675 => "001000101101010110111000",
34676 => "000110101001111111010001",
34677 => "000011001110101011111101",
34678 => "111111011101100110101101",
34679 => "111011111101111010111010",
34680 => "111000011111110001010100",
34681 => "110100101110001011011001",
34682 => "110001000111011000110110",
34683 => "101110110111001011110110",
34684 => "101101110010010101101010",
34685 => "101101010000000111100100",
34686 => "101110001001100110001110",
34687 => "110000001101100100011110",
34688 => "110001111000010110101000",
34689 => "110011010111101100011000",
34690 => "110101101010001100001001",
34691 => "111000100001110001011011",
34692 => "111011001110111101000111",
34693 => "111101110111010110011110",
34694 => "000000010111101100011111",
34695 => "000010010000101111001100",
34696 => "000100011000110101111100",
34697 => "000110001010111001101001",
34698 => "000101011001101111011110",
34699 => "000010111100111011011100",
34700 => "000000010110100100101110",
34701 => "111101101101011100110100",
34702 => "111011101111101000010011",
34703 => "111010111010001101100000",
34704 => "111011010011100100000001",
34705 => "111100100010001100101110",
34706 => "111110001000011010100001",
34707 => "111111101101100111001100",
34708 => "111111110101100011000001",
34709 => "111111110000110010000001",
34710 => "000001001101000000110100",
34711 => "000010001010011011101010",
34712 => "000010101001010001000100",
34713 => "000011010011000111001111",
34714 => "000011011011111101010110",
34715 => "000100100011011110111110",
34716 => "000110010110011010011110",
34717 => "001000001000001100000011",
34718 => "001011010000011000101001",
34719 => "001110110011111010010100",
34720 => "010001101111111101101010",
34721 => "010011110110110100110000",
34722 => "010100011001011000011100",
34723 => "010010101010100100000000",
34724 => "001101111000110011111000",
34725 => "001000001110110110010110",
34726 => "000011010101001101010111",
34727 => "111110011100001001110011",
34728 => "111011111011011010101110",
34729 => "111100001000110101010011",
34730 => "111100100001101010110011",
34731 => "111100101111010011100110",
34732 => "111011010001111100100010",
34733 => "111000010111001101110110",
34734 => "110110111101111010010100",
34735 => "110111101101100100111110",
34736 => "111010011110100100001000",
34737 => "111110011100110001001101",
34738 => "000010110101010110110100",
34739 => "001000000010110011010110",
34740 => "001100101001110100101100",
34741 => "001111110110100100000100",
34742 => "010010101001110001011010",
34743 => "010100111011110010100010",
34744 => "010101100101111111110010",
34745 => "010011100111010101110110",
34746 => "010000000011110001100000",
34747 => "001100011100001011001010",
34748 => "001000000100101001011110",
34749 => "000010111001011111100111",
34750 => "111110101011110011000011",
34751 => "111101110010011101111010",
34752 => "000000011100110110101000",
34753 => "000011011111011010001000",
34754 => "000100111111111001101100",
34755 => "000101011100110011011111",
34756 => "000101000011101010001000",
34757 => "000011111000100100001011",
34758 => "000010000010011010111000",
34759 => "111111111100010101100001",
34760 => "111101011101001101010000",
34761 => "111001111000111001101101",
34762 => "110110001010101001001100",
34763 => "110011110011011000000010",
34764 => "110011011001100000011100",
34765 => "110100001000011011000011",
34766 => "110100000110000101101000",
34767 => "110011011101111010000110",
34768 => "110100101000010000010100",
34769 => "111000100110101000010111",
34770 => "111101100110001011010000",
34771 => "000001000110101110110001",
34772 => "000010101110101010001111",
34773 => "000011001101000110111011",
34774 => "000010100101101101100010",
34775 => "000000101100100001000011",
34776 => "111101101100110000011001",
34777 => "111010001010111001001011",
34778 => "110101111111010100110000",
34779 => "110001010010011111110000",
34780 => "101110000000010001111110",
34781 => "101101001101000001011010",
34782 => "101110001111100101010110",
34783 => "110000101101111010001000",
34784 => "110100001011101001001001",
34785 => "111000010011001001101100",
34786 => "111101000100011010011111",
34787 => "000001101101111111110101",
34788 => "000100111111000001111100",
34789 => "000110010010101111110011",
34790 => "000110000111100101100000",
34791 => "000101110100100010000111",
34792 => "000110110000000011001110",
34793 => "001000110111001101111001",
34794 => "001011010000100001100101",
34795 => "001101100001011101101010",
34796 => "001111001010001000101100",
34797 => "001111111000011101111010",
34798 => "010000001110011001001010",
34799 => "001111111000011111000000",
34800 => "001101101001100100110110",
34801 => "001001101110001101110100",
34802 => "000101101101000101001000",
34803 => "000010001100100110100111",
34804 => "111110111110011100111000",
34805 => "111100110001011001001001",
34806 => "111100010001000101101001",
34807 => "111101010011011000001000",
34808 => "111111011101001101101000",
34809 => "000010010100100100101101",
34810 => "000110001101100011100100",
34811 => "001010111111001001100000",
34812 => "001111000011101110001000",
34813 => "010001001110011001000010",
34814 => "010001011000011100110100",
34815 => "010000000001000100111110",
34816 => "001101011100000100100000",
34817 => "001001010010101011100100",
34818 => "000011111000111111100000",
34819 => "111110101100111000100110",
34820 => "111010101111001001101001",
34821 => "110111011001100011101111",
34822 => "110100001000001001011000",
34823 => "110001111111100101110010",
34824 => "110001110100111110010010",
34825 => "110011010010011111001100",
34826 => "110101100101111011011011",
34827 => "111000000110100010100100",
34828 => "111011001100001101101001",
34829 => "111110100100101111100010",
34830 => "000000110011011111101011",
34831 => "000001001101101110111100",
34832 => "111111101010110000000001",
34833 => "111100101000101110010001",
34834 => "111001001001011100010101",
34835 => "110110001111011110011001",
34836 => "110100100101111101001001",
34837 => "110011001011111011011000",
34838 => "110001111101101111101100",
34839 => "110010100001111101101010",
34840 => "110100001011101101111001",
34841 => "110101111010010100110010",
34842 => "110111111100100011101000",
34843 => "111001011101111000000000",
34844 => "111001101110110111100101",
34845 => "111000110011101001000000",
34846 => "110111011000110111100100",
34847 => "110110011111001011011000",
34848 => "110110000100011100001110",
34849 => "110101101010101001110110",
34850 => "110101100011000000010010",
34851 => "110110110111100000110010",
34852 => "111001011011000000110010",
34853 => "111011000011110000001001",
34854 => "111011101100010010011101",
34855 => "111100101001000111001100",
34856 => "111110011100110110011011",
34857 => "000001100100010010011101",
34858 => "000100011100101111100001",
34859 => "000101101011100111001001",
34860 => "000111001001110100001000",
34861 => "001001110101011000101111",
34862 => "001011101110101011000111",
34863 => "001011101011111110110000",
34864 => "001011010100010011110010",
34865 => "001011001100010111011110",
34866 => "001001001011100011110000",
34867 => "000101100010000000110111",
34868 => "000010011101000101000000",
34869 => "111111101000011100111001",
34870 => "111100001011111101001110",
34871 => "111001001000110111010010",
34872 => "111000100010100101111111",
34873 => "111010110111111100010011",
34874 => "111110010100110011000101",
34875 => "000010010101010001111101",
34876 => "000111100111110011100100",
34877 => "001100111110001111010010",
34878 => "001111101111000101010110",
34879 => "001110111111110011110100",
34880 => "001101000000001110110100",
34881 => "001011101001010000011001",
34882 => "001001101011111111110101",
34883 => "000101001100110001010110",
34884 => "111110001011110110101010",
34885 => "110111001100111110001100",
34886 => "110001100011110000100110",
34887 => "101011000010000011011100",
34888 => "100100011100100010011101",
34889 => "100010001000000101001010",
34890 => "100100010110011101110111",
34891 => "101001001000101000001100",
34892 => "101111110001111100010000",
34893 => "110110011100100000011101",
34894 => "111100001000110100100101",
34895 => "000001111011100111111101",
34896 => "000111100001100011010110",
34897 => "001100010010010111011110",
34898 => "010000000110100101111110",
34899 => "010010000010100111110100",
34900 => "010010001110111001011100",
34901 => "010001111000110100010110",
34902 => "010001100011000111101110",
34903 => "010000001011100110000110",
34904 => "001100100001011010001100",
34905 => "001001001000110101000100",
34906 => "001000011001111011011000",
34907 => "000111110110001101011000",
34908 => "000110001001010101100100",
34909 => "000100011011000101000110",
34910 => "000011010110001000001010",
34911 => "000011010101101000110001",
34912 => "000010111111100101101001",
34913 => "000010000011010000100111",
34914 => "000011010101101010110110",
34915 => "000111001000111101000001",
34916 => "001010010111010010111111",
34917 => "001010111101001000011000",
34918 => "001010000001010111010001",
34919 => "001001000010100101101111",
34920 => "000111010100111000001011",
34921 => "000100100111011111110111",
34922 => "000001110010110100101000",
34923 => "000000011101001101100101",
34924 => "000001100010010000101110",
34925 => "000010110111001101011110",
34926 => "000011110000110101000111",
34927 => "000101011010110010011010",
34928 => "000110010011110110111111",
34929 => "000101001111011110100011",
34930 => "000010000101010111011110",
34931 => "111100110111111111001100",
34932 => "110110000101110001111000",
34933 => "101101000110001011000100",
34934 => "100100101001010000011101",
34935 => "100001011010111110001111",
34936 => "100001111010001011011110",
34937 => "100010101000000111000101",
34938 => "100100000011000001100111",
34939 => "101000010010110010100100",
34940 => "101111100010101001001000",
34941 => "110111110000010101001111",
34942 => "111111110010000000100000",
34943 => "000110001111100110000100",
34944 => "001001001011011100000101",
34945 => "001001011011111011101000",
34946 => "001000100110000100000101",
34947 => "000111011101111011000001",
34948 => "000110110100001011100000",
34949 => "000110000100001011000101",
34950 => "000100110111100111010001",
34951 => "000011111011010000011100",
34952 => "000011100111001011110011",
34953 => "000011010010001100011011",
34954 => "000001011100011010101111",
34955 => "111110011000001001101011",
34956 => "111011110100001000001111",
34957 => "111010000101101101011101",
34958 => "111001000000011101100110",
34959 => "111000110001010001110110",
34960 => "111001110010000011000011",
34961 => "111100000100010000010110",
34962 => "111111000010101011000001",
34963 => "000010111111111001000011",
34964 => "000111101101111111001110",
34965 => "001011100011110101010010",
34966 => "001110010101110100000100",
34967 => "010000011100111111010100",
34968 => "010000111100010010010000",
34969 => "001111110010011110111000",
34970 => "001110011001110110110110",
34971 => "001101011010000100010110",
34972 => "001011111100101110000000",
34973 => "001001000100001010110100",
34974 => "000101001011011100101010",
34975 => "000001011010101101111001",
34976 => "111110001010010001001100",
34977 => "111011001000000010010111",
34978 => "111000000111110110000010",
34979 => "110101110111111011101010",
34980 => "110101011011011010001110",
34981 => "110110111101001011110100",
34982 => "111010010010011110110010",
34983 => "111110100000110000101000",
34984 => "000010001010011101111101",
34985 => "000101001110011010011010",
34986 => "000111101111000001100001",
34987 => "001000111001000111110100",
34988 => "001000100000000101100100",
34989 => "000110001110100000000100",
34990 => "000010000111001110101010",
34991 => "111101100101000101000110",
34992 => "111001111101101001000111",
34993 => "110111010111100110011000",
34994 => "110101000101100100001110",
34995 => "110011100111001011000100",
34996 => "110011101111110110101000",
34997 => "110100100001001000100101",
34998 => "110101001111000010110110",
34999 => "110101110010001111010111",
35000 => "110110001111001000111110",
35001 => "110111000110000001111010",
35002 => "110110110100010111100100",
35003 => "110100001100010001010100",
35004 => "110001100000010100010110",
35005 => "110001000110001000100000",
35006 => "110010100101011110000000",
35007 => "110011111101000101110110",
35008 => "110101000101101111110100",
35009 => "110111100000101000100110",
35010 => "111010101111100010011011",
35011 => "111110010111101010011000",
35012 => "000010011010011011101100",
35013 => "000101111100011100111111",
35014 => "001001111001011011010111",
35015 => "001110101001100111100010",
35016 => "010001100000110101110100",
35017 => "010001001001010101010000",
35018 => "001111001111010001101100",
35019 => "001101111001011010110110",
35020 => "001101011110001001001100",
35021 => "001100111010011101100110",
35022 => "001011001100000000100011",
35023 => "001000000110010101100110",
35024 => "000101000000001001101010",
35025 => "000010111110000101011100",
35026 => "000001110010100110000011",
35027 => "000001001010101100110110",
35028 => "000000011010011110100100",
35029 => "111111110111011110101010",
35030 => "000001010000001100000001",
35031 => "000100110001101011110000",
35032 => "001000111001110101001110",
35033 => "001100010001001010110000",
35034 => "001110111101001011000110",
35035 => "010001001101111000001010",
35036 => "010010011010110111101000",
35037 => "010010100100110011010010",
35038 => "010000111111011111110110",
35039 => "001100100000010100101000",
35040 => "000101101111101100110001",
35041 => "111100110011111100101011",
35042 => "110001111111000101110110",
35043 => "101000101000110011010110",
35044 => "100100001110010011100001",
35045 => "100100010100111011001101",
35046 => "100110001000011000011001",
35047 => "101001100000110010100010",
35048 => "101111011110100011011100",
35049 => "110101111101111111111100",
35050 => "111011011101101100110100",
35051 => "111111110110101010110010",
35052 => "000010011110110000000001",
35053 => "000100000001111101110010",
35054 => "000100111000101011001111",
35055 => "000100010010110010101100",
35056 => "000010100010100011111011",
35057 => "000000000001011101111101",
35058 => "111101100010001010001011",
35059 => "111100101110100001111000",
35060 => "111110001111010000001111",
35061 => "000000110100100111000001",
35062 => "000010001000101100100100",
35063 => "000001001101001001101110",
35064 => "111111001100111011001111",
35065 => "111101011010101101000011",
35066 => "111100000100111001011000",
35067 => "111010100110111100110101",
35068 => "111001101000100010100100",
35069 => "111011010001011100001011",
35070 => "111111011100000011111010",
35071 => "000011010011001011100001",
35072 => "000101101111111100100010",
35073 => "000111111000001100111101",
35074 => "001001000000111010010011",
35075 => "001000000111101110101111",
35076 => "000110011101010010010001",
35077 => "000100101010011100100001",
35078 => "000011001011100011000110",
35079 => "000011010110100001111110",
35080 => "000100001111000111111011",
35081 => "000101010110001100111000",
35082 => "001000010001000000001011",
35083 => "001011101000100101010011",
35084 => "001101010000100110001000",
35085 => "001101011111101011011100",
35086 => "001100010010001010011100",
35087 => "001001100010001101010010",
35088 => "000110001000010101100010",
35089 => "000010000001000101100101",
35090 => "111101001001110010110110",
35091 => "111000011010001100011010",
35092 => "110100111000010000010100",
35093 => "110011110110001110011110",
35094 => "110101010010101011001110",
35095 => "110111101100100100110001",
35096 => "111010010101000011010011",
35097 => "111101011100111000101101",
35098 => "000000101111111100101110",
35099 => "000010101000010100001000",
35100 => "000010100011100011111100",
35101 => "000010010101011101101111",
35102 => "000010110000110011011000",
35103 => "000011011010010010110110",
35104 => "000011111010100001101100",
35105 => "000010101000111010100000",
35106 => "111111001100100000011111",
35107 => "111011000111000010101101",
35108 => "110111001111000011101001",
35109 => "110100100011011001101100",
35110 => "110011010000110000101100",
35111 => "110010010101111100101100",
35112 => "110001100100011100011010",
35113 => "110001011000101000101110",
35114 => "110011000010101111101100",
35115 => "110110101111000011011100",
35116 => "111010110000110101010000",
35117 => "111110101000010111101001",
35118 => "000010001101100100000011",
35119 => "000101000011110100010001",
35120 => "000111010001001110011100",
35121 => "001000010110111001011000",
35122 => "001000010001000110011001",
35123 => "000110111011111101111001",
35124 => "000011110100110000001001",
35125 => "111111111100111001111100",
35126 => "111101000001001101010111",
35127 => "111100000010000100111010",
35128 => "111100000000111010011110",
35129 => "111010111110111000111110",
35130 => "111001111001101010010100",
35131 => "111010010101011001001110",
35132 => "111011011110110101101111",
35133 => "111100001001110101100101",
35134 => "111100000000011011111110",
35135 => "111100011110101100101111",
35136 => "111110110100101010101101",
35137 => "000001101011011001111100",
35138 => "000011100101110001101110",
35139 => "000100111001000110100101",
35140 => "000110010101101010000110",
35141 => "000111000100100000000001",
35142 => "000110011111001111010000",
35143 => "000110001101011000101100",
35144 => "000110000011100011000001",
35145 => "000100010001001100110101",
35146 => "000001000000100101101010",
35147 => "111101100001000111110101",
35148 => "111011100110110011000011",
35149 => "111011100001010110110001",
35150 => "111100000110000101011000",
35151 => "111110000001011011000001",
35152 => "000001000101110000001010",
35153 => "000011111110111111001111",
35154 => "000110100011000000000100",
35155 => "000111110011101110100010",
35156 => "000111100011100000011011",
35157 => "000110011000111111011101",
35158 => "000011101000111100010010",
35159 => "111111111100100100011010",
35160 => "111100010110110001000110",
35161 => "111000000010010111111011",
35162 => "110010011011010100111010",
35163 => "101100100001110000011010",
35164 => "101000110001010101011110",
35165 => "101000111010000110001000",
35166 => "101100001011010100000100",
35167 => "110000111011100111010100",
35168 => "110101110011011101001100",
35169 => "111010110101001001000100",
35170 => "000000110100110111100010",
35171 => "000110001000011111000010",
35172 => "001001011110110011100000",
35173 => "001100011100110101111100",
35174 => "001110001011001110011010",
35175 => "001100101001010000000010",
35176 => "001010000000001111011110",
35177 => "001000101100110001010110",
35178 => "001000100101001110101100",
35179 => "001000011110110011111000",
35180 => "000110011110111001110000",
35181 => "000010110101001110111111",
35182 => "000000010001100100110011",
35183 => "111111010010111111110100",
35184 => "111110000010101010111110",
35185 => "111011111100101000001001",
35186 => "111010100000000011000010",
35187 => "111010010011110111011001",
35188 => "111010010101001101000000",
35189 => "111011010110101000100000",
35190 => "111110110101010001011000",
35191 => "000011101100001100011001",
35192 => "001000010101100101100011",
35193 => "001011101010101110000000",
35194 => "001100100000010001111000",
35195 => "001010001000101011100001",
35196 => "000100001101001100111001",
35197 => "111011111111011001101010",
35198 => "110100110100110100101011",
35199 => "110000110010000101100010",
35200 => "101111001100100000010010",
35201 => "101111100100110011011000",
35202 => "110010010011000010000010",
35203 => "110110010110010001110010",
35204 => "111010001110101010101010",
35205 => "111101010000010100100100",
35206 => "111111100100010000111110",
35207 => "000010010001101000100111",
35208 => "000100101011111011110110",
35209 => "000100110000000010011101",
35210 => "000010111110111010000010",
35211 => "000001011110001110100011",
35212 => "000001110000100111000001",
35213 => "000011000101101010101101",
35214 => "000011101011010101001001",
35215 => "000101001011110110110001",
35216 => "001000101100010011001100",
35217 => "001011000111101001011110",
35218 => "001010010010000101111100",
35219 => "000110011011010111011110",
35220 => "000001100000001001011101",
35221 => "111101011111111001101110",
35222 => "111001110111100111101111",
35223 => "110110111111101101011010",
35224 => "110111000010010110100001",
35225 => "111001100000100101011011",
35226 => "111100000100100010100010",
35227 => "111101110110101100011110",
35228 => "111111011110011011100111",
35229 => "000000111011110111000100",
35230 => "000001010001110100011000",
35231 => "000000011101010001110111",
35232 => "111111101001101001101100",
35233 => "111111111011010000000011",
35234 => "000000111001001000111101",
35235 => "000001011110010000110101",
35236 => "000001111001110010110100",
35237 => "000010101101000010011000",
35238 => "000011100101000111010110",
35239 => "000100011111001010010100",
35240 => "000101011101100110010001",
35241 => "000101110100111010111000",
35242 => "000100110000000111011110",
35243 => "000010010110110111000111",
35244 => "111111011111100011111001",
35245 => "111101010001101010001001",
35246 => "111100110101101010111000",
35247 => "111101111100000100110111",
35248 => "111111101011010011100100",
35249 => "000001110010101011011000",
35250 => "000011100000110011010101",
35251 => "000100010100011010100111",
35252 => "000100101011110000001101",
35253 => "000100110001000100000100",
35254 => "000100100011110010101010",
35255 => "000100001111111011011101",
35256 => "000100101011010100000000",
35257 => "000110111111111011010100",
35258 => "001010110000110011010110",
35259 => "001110011101100001101110",
35260 => "010001010100000110001100",
35261 => "010011010101000000000100",
35262 => "010100010010101111100110",
35263 => "010011011100010001110010",
35264 => "010000111000110010111100",
35265 => "001101011011010011011010",
35266 => "001001011100000100111010",
35267 => "000101100111110101111100",
35268 => "000010101010100110101011",
35269 => "000000110101011111011100",
35270 => "000000001101110101110100",
35271 => "000000010101100110010111",
35272 => "000000111110101111100001",
35273 => "000001111111110110001111",
35274 => "000010100011111011100110",
35275 => "000010100010000111011100",
35276 => "000010010001011000011100",
35277 => "000001000100001111001100",
35278 => "111101111101011000010011",
35279 => "111001010111101000110110",
35280 => "110100100001000110011011",
35281 => "110000000111000001011110",
35282 => "101101001011001000001100",
35283 => "101101000011000010000100",
35284 => "101111001100100111001100",
35285 => "110001101101001101000000",
35286 => "110011110000100001101010",
35287 => "110110000010100100101000",
35288 => "111000111111101100010001",
35289 => "111011111110100011101110",
35290 => "111110101110000110100101",
35291 => "000001000011100000100001",
35292 => "000010000110110011101101",
35293 => "000010011101111010110101",
35294 => "000010111110111010011010",
35295 => "000001111000011001110010",
35296 => "111110001001011111110011",
35297 => "111001111010111101001001",
35298 => "110111011001111000000100",
35299 => "110110100101011001000010",
35300 => "110101100101010011000011",
35301 => "110011110101000101101110",
35302 => "110011010110001111110110",
35303 => "110100100011001111101100",
35304 => "110110010111100110001010",
35305 => "111001110011110110110000",
35306 => "111111010010010000011011",
35307 => "000101000101011000111000",
35308 => "001010010110111101010011",
35309 => "001111000001111011010010",
35310 => "010010101011000101011010",
35311 => "010101001000000100000000",
35312 => "010110011110011110100100",
35313 => "010110001011001010010010",
35314 => "010010111010000111001100",
35315 => "001100010100011001110010",
35316 => "000011111110100100001111",
35317 => "111100000101111010000010",
35318 => "110101100100011101010011",
35319 => "101111011110001100111000",
35320 => "101001110000111100000110",
35321 => "100110110001101011011101",
35322 => "101000001110101011001000",
35323 => "101101010111000101011110",
35324 => "110100000001010110100101",
35325 => "111010100101011010001011",
35326 => "000000110001000100100000",
35327 => "000110110000110001101010",
35328 => "001100101011000011101000",
35329 => "010001110100100110100000",
35330 => "010100111101011001001000",
35331 => "010101111010110100011010",
35332 => "010101010011001000010110",
35333 => "010011001011011011001010",
35334 => "001111000010010100010100",
35335 => "001001001110010100101001",
35336 => "000011110101010100110111",
35337 => "000000000010000011111111",
35338 => "111101010001010001001010",
35339 => "111010100101000011010010",
35340 => "110110101110011010100100",
35341 => "110010110110110110111100",
35342 => "110001001101000001110000",
35343 => "110000101000111001111100",
35344 => "110000011000010101111110",
35345 => "110001110111000100000100",
35346 => "110100101100001101100000",
35347 => "110111111101100000101000",
35348 => "111011011111101001000001",
35349 => "111101011011100011101101",
35350 => "111100001001010100011110",
35351 => "111001001011110110110011",
35352 => "110110110000010011101000",
35353 => "110101000011010101100101",
35354 => "110011110011000011000010",
35355 => "110011001110100101000100",
35356 => "110011101001101001110100",
35357 => "110101100011011100000011",
35358 => "110111110111111010101010",
35359 => "111000100100000100011100",
35360 => "111001000010010100111100",
35361 => "111100000010001111011001",
35362 => "000000000011100010011011",
35363 => "000010010011011000110000",
35364 => "000010110010110111010110",
35365 => "000010100101101001110001",
35366 => "000010101011010000001010",
35367 => "000010111110110110110110",
35368 => "000010000110001110100110",
35369 => "000000111001110001110100",
35370 => "000001100110111010010010",
35371 => "000011100101101101111011",
35372 => "000101000010110110101101",
35373 => "000101010101110010110010",
35374 => "000101000001011010110001",
35375 => "000101011100101111001001",
35376 => "000110111100011011000101",
35377 => "001000001110010100110000",
35378 => "001000101101010001110100",
35379 => "001001101000111000011000",
35380 => "001011000111001101100001",
35381 => "001010111110100101111010",
35382 => "001000111111100010111100",
35383 => "000110110001101010101110",
35384 => "000100010110010000000001",
35385 => "000001011000010111000100",
35386 => "111110111101010101100011",
35387 => "111110011111010011100011",
35388 => "111111011011000010111010",
35389 => "111111101111010111111100",
35390 => "111111101101001100101010",
35391 => "000000011101000010100000",
35392 => "000000100111100010011011",
35393 => "111110101110101001011010",
35394 => "111011101110010010011110",
35395 => "111001011010001100001010",
35396 => "110111110001001001000110",
35397 => "110101110100011100001011",
35398 => "110100000001111100010001",
35399 => "110011001010110100011000",
35400 => "110011101110001010001010",
35401 => "110101110100000010101000",
35402 => "111000010000001111010011",
35403 => "111010000011001100100110",
35404 => "111010110111011110011000",
35405 => "111010100100100110001100",
35406 => "111001011011101111000101",
35407 => "110111001001001100101000",
35408 => "110011110011110001011010",
35409 => "110000100011000001100000",
35410 => "101110011010101000011100",
35411 => "101110101111001101000110",
35412 => "110001111001111000011100",
35413 => "110110101001000010111000",
35414 => "111011101101100110110110",
35415 => "000000101010101111011000",
35416 => "000101011000110001110011",
35417 => "001001000011001110111010",
35418 => "001011000000010111001001",
35419 => "001011111010011111010010",
35420 => "001100000110010110000010",
35421 => "001011011101110000010011",
35422 => "001010010100011011100110",
35423 => "001000111011111111010110",
35424 => "000111101110010111101001",
35425 => "000111000001110111110011",
35426 => "000111000100000111000011",
35427 => "000111101110110101010111",
35428 => "001000010010110100010010",
35429 => "001000011101011110011011",
35430 => "001000110100110010001010",
35431 => "001001111001100000010000",
35432 => "001010111000010011000010",
35433 => "001010101101110011011111",
35434 => "001010100010110111001000",
35435 => "001011101011010100110110",
35436 => "001101011111101111101000",
35437 => "001111001011000010000110",
35438 => "010000000011010011100100",
35439 => "001111111010010011101000",
35440 => "001111011000000111111110",
35441 => "001110011010011110110000",
35442 => "001100010100111010101000",
35443 => "001001100000011011100000",
35444 => "000111001000011000100111",
35445 => "000101000111110110000011",
35446 => "000010111000001100010110",
35447 => "000001000001111010011100",
35448 => "000000000101110100001110",
35449 => "111111011110011101100101",
35450 => "111101101101010110100011",
35451 => "111001111001111101101110",
35452 => "110101100011101000000000",
35453 => "110001110110011110011010",
35454 => "101110110101101101000110",
35455 => "101101100010001000001000",
35456 => "101110010110001011111110",
35457 => "110000100111110000010110",
35458 => "110011110101011101101100",
35459 => "111000001110011010010111",
35460 => "111110011000010100101001",
35461 => "000100101011100110110000",
35462 => "001001011000000101100011",
35463 => "001100110111000101010010",
35464 => "001111000000010010001000",
35465 => "010000000101100110001100",
35466 => "010000110101110110100110",
35467 => "010000001010001111110110",
35468 => "001101001001110011011100",
35469 => "001000011101000011101010",
35470 => "000011101101010110101100",
35471 => "000000010110100111000110",
35472 => "111110001100111000111100",
35473 => "111100001111000100011001",
35474 => "111001010011110001110110",
35475 => "110110001111011011010101",
35476 => "110101010011001011100010",
35477 => "110101110000101011001100",
35478 => "110110000011000111111111",
35479 => "110110001111101011000000",
35480 => "110110011010010010101101",
35481 => "111000000110111001100000",
35482 => "111101000001011011011011",
35483 => "000011101101101001100111",
35484 => "001010010101100101010011",
35485 => "010000101111111011000000",
35486 => "010110011001101101000100",
35487 => "011001111101100110111010",
35488 => "011011011000110000000111",
35489 => "011011011111000101100000",
35490 => "011010010001110101011100",
35491 => "010111000110011000000000",
35492 => "010001001010010001100010",
35493 => "001001101110111101000010",
35494 => "000011110000011101110011",
35495 => "111111111111111000100101",
35496 => "111101110001110100011100",
35497 => "111100100010110100000001",
35498 => "111011011110110010101010",
35499 => "111010100100100011110011",
35500 => "111010110001101001100010",
35501 => "111100110101101111001110",
35502 => "111110100100011111100010",
35503 => "111100100100101100010011",
35504 => "110111110110101010001101",
35505 => "110010001010101110000010",
35506 => "101011011101100001111100",
35507 => "100110011110010001101011",
35508 => "100101011100011100111111",
35509 => "100111000101010010111011",
35510 => "101010011011000100110110",
35511 => "101111010010010000010100",
35512 => "110100100110011101011111",
35513 => "111000000110100100010100",
35514 => "111000110011110111010010",
35515 => "111001001111010010010110",
35516 => "111011000100100001111101",
35517 => "111100001111111010001001",
35518 => "111011000100111010110000",
35519 => "111001001101110100100010",
35520 => "111001000101010000010010",
35521 => "111001111111001101010100",
35522 => "111001100110010101011010",
35523 => "111000100101101101001001",
35524 => "111001011100011000110111",
35525 => "111011100101001011100000",
35526 => "111100010100100000001111",
35527 => "111010010001111000100001",
35528 => "110110010001000110111111",
35529 => "110100001011100001101010",
35530 => "110110011110011101101011",
35531 => "111010001100110111111010",
35532 => "111110000011111011011110",
35533 => "000100010011100001011110",
35534 => "001101000000001101100010",
35535 => "010101110101001101111000",
35536 => "011011001110001111010001",
35537 => "011100001100011100010001",
35538 => "011011010000100011001001",
35539 => "010111100010000011000100",
35540 => "001111101011001000010000",
35541 => "000111001100000110111001",
35542 => "000001001001001001101100",
35543 => "111101101111111000111111",
35544 => "111011111100011110000010",
35545 => "111011010100001111110010",
35546 => "111101001100100000000000",
35547 => "000000110100110101001101",
35548 => "000011100000001101101011",
35549 => "000100110011111111101010",
35550 => "000101011101111001110001",
35551 => "000100110010010010111100",
35552 => "000001101011011000000100",
35553 => "111101000001110100111010",
35554 => "111001000111010101110001",
35555 => "110110101111000100101100",
35556 => "110101101110110110010111",
35557 => "110110011100110001011111",
35558 => "111000011111101010101000",
35559 => "111010011111000000111011",
35560 => "111011100010111110000101",
35561 => "111011000001100001000000",
35562 => "111000001011000010011000",
35563 => "110011110101001011111000",
35564 => "101111011011110010000000",
35565 => "101011100011010010101100",
35566 => "101001001001110000011100",
35567 => "101000100110001110011010",
35568 => "101001010101101010110010",
35569 => "101011100100000000100110",
35570 => "101111000100000001100010",
35571 => "110010111000001000100010",
35572 => "110101101101101110110101",
35573 => "110110101001011001101010",
35574 => "110110101111110010100010",
35575 => "110110111010110011100000",
35576 => "110110011100101010110100",
35577 => "110101000001100101010100",
35578 => "110011010010100101001110",
35579 => "110010100110010111110100",
35580 => "110011010101001011001100",
35581 => "110100100001000001111000",
35582 => "110110001101110111111101",
35583 => "111000100100011101110001",
35584 => "111011001001101101001000",
35585 => "111110001001001000110000",
35586 => "000001001111000001011101",
35587 => "000011110100100010011100",
35588 => "000110000000100000001100",
35589 => "001000011101001111101010",
35590 => "001011011001000110111111",
35591 => "001101101001110100000100",
35592 => "001111001001001001001010",
35593 => "010001001010010100101110",
35594 => "010010111001101001111000",
35595 => "010010101010110010001100",
35596 => "010000101111010111101010",
35597 => "001110100111001011110010",
35598 => "001101011101010000110100",
35599 => "001101000000110100101010",
35600 => "001100001011011001011110",
35601 => "001011000101100101101110",
35602 => "001011010001100010000100",
35603 => "001101000101101001010100",
35604 => "001110100110010001000010",
35605 => "001110100010110100111100",
35606 => "001110001010111111001000",
35607 => "001110110110001110010010",
35608 => "001111100101101101001000",
35609 => "001110101011010010001010",
35610 => "001100101000111101000110",
35611 => "001010110110000000011110",
35612 => "001001011100001101101010",
35613 => "001000010011011110000011",
35614 => "000111101010111111011000",
35615 => "001000001101111011100111",
35616 => "001001011100100110011110",
35617 => "001001110110000101010110",
35618 => "001001110010000001110011",
35619 => "001001000110011010011110",
35620 => "000110110010011011111111",
35621 => "000100100110000010111100",
35622 => "000011001101100010000010",
35623 => "000000110011000100000110",
35624 => "111100111101111001011101",
35625 => "111000011001110111010111",
35626 => "110100101000000010011100",
35627 => "110011001101010010111100",
35628 => "110011101010110111110000",
35629 => "110101000111001100111111",
35630 => "110111001011000011111000",
35631 => "111001101100111010001001",
35632 => "111100110010010100001100",
35633 => "111111011101110001010110",
35634 => "000000001000011101110011",
35635 => "111110101101001010001001",
35636 => "111100111101011001000110",
35637 => "111011101110001010101100",
35638 => "111010000000110000111101",
35639 => "111000100000011010001011",
35640 => "111000101011010011110011",
35641 => "111001011110001001010110",
35642 => "111001111100010010010010",
35643 => "111011100100000111011010",
35644 => "111111010000100100111000",
35645 => "000011000100101011111110",
35646 => "000100111001010101010000",
35647 => "000101001100110010101111",
35648 => "000101000110100001111011",
35649 => "000101001010010011010000",
35650 => "000101110110010000110001",
35651 => "000110011010101001101011",
35652 => "000101101000111001111010",
35653 => "000100001111101000110111",
35654 => "000100100100110111110000",
35655 => "000111011010111110101011",
35656 => "001010101011101110011111",
35657 => "001011011111010010110000",
35658 => "001000010110110001001010",
35659 => "000010101010101001101101",
35660 => "111100011110100001000000",
35661 => "110101100010101110001110",
35662 => "101111011011111011101000",
35663 => "101101010001101001110110",
35664 => "101101001011110110111010",
35665 => "101100100001101010110100",
35666 => "101101100011110111001110",
35667 => "110010001010100111011100",
35668 => "111000010110011011011111",
35669 => "111101110100110011001000",
35670 => "000010001010000110111001",
35671 => "000101011001110110010000",
35672 => "000111101100101001011110",
35673 => "001001001011100100101000",
35674 => "001001101000101110010000",
35675 => "001001101111101001001011",
35676 => "001001000110011010000000",
35677 => "000110000010100110011011",
35678 => "000011001111010100001011",
35679 => "000011100110101111001001",
35680 => "000011101111100000110001",
35681 => "000000110101100010111001",
35682 => "111100100000001010011100",
35683 => "111000000101111110010011",
35684 => "110100100101111101000000",
35685 => "110011000001100110001010",
35686 => "110010010010110101110110",
35687 => "110001111010100100011010",
35688 => "110100100111010001011110",
35689 => "111011001010011111110000",
35690 => "000001111110010111001100",
35691 => "000111000001110101001111",
35692 => "001011011110111110001010",
35693 => "001111100100110011000000",
35694 => "010001110001100110000100",
35695 => "010001001010101101111000",
35696 => "001111010011100100101010",
35697 => "001110001011101110101000",
35698 => "001101001000101001110000",
35699 => "001010100001001100011110",
35700 => "000110111001011010110011",
35701 => "000100010010011111001000",
35702 => "000011000011001100001000",
35703 => "000010010100011100001101",
35704 => "000010010110111101111100",
35705 => "000011000000011101111010",
35706 => "000011000110011101011010",
35707 => "000010010011101110110100",
35708 => "000001001010100010101100",
35709 => "000000100111100100100011",
35710 => "000000100001110111100111",
35711 => "111111110010100010001000",
35712 => "111110110110001000100111",
35713 => "111110100011100101100011",
35714 => "111110011100001011100011",
35715 => "111101010001100100101010",
35716 => "111010101110101110010101",
35717 => "111000101011111101100010",
35718 => "111000000011011000011111",
35719 => "110111100111000011100001",
35720 => "110111111000001001010010",
35721 => "111010010110001101011100",
35722 => "111110001111011101010000",
35723 => "000001000000001011001110",
35724 => "000001010010100111101100",
35725 => "000000001001001010010110",
35726 => "111101111011011100101100",
35727 => "111001110101010101001101",
35728 => "110100011100111100011011",
35729 => "101111010011101101110000",
35730 => "101011000010110111110100",
35731 => "100111000101001111110101",
35732 => "100011111100000100111111",
35733 => "100100000101111110110001",
35734 => "100111100000011111110101",
35735 => "101010111001100110110110",
35736 => "101101000001111101110010",
35737 => "101111011000110111001010",
35738 => "110001111101000100101000",
35739 => "110011101000010111010100",
35740 => "110101001011011001101110",
35741 => "110110110111010010110100",
35742 => "111000000100101010111000",
35743 => "111001110111100001111011",
35744 => "111100100000110110000001",
35745 => "111111000101000001011101",
35746 => "000001010010011101100100",
35747 => "000010011010000000101000",
35748 => "000010011100100111011100",
35749 => "000010010011000000011000",
35750 => "000001101101010101101110",
35751 => "000000000111000110001100",
35752 => "111101101000001000000011",
35753 => "111011100010110100101011",
35754 => "111011001100101011100110",
35755 => "111100100000000011011001",
35756 => "111110101110011111010101",
35757 => "000000111101100011100011",
35758 => "000011010010101101000110",
35759 => "000110001110000110001010",
35760 => "001000100111001000100010",
35761 => "001010010000100101011010",
35762 => "001100011010010111110000",
35763 => "001110110011111110001000",
35764 => "001111110011010001110100",
35765 => "001110100110000111101010",
35766 => "001101011001011111010110",
35767 => "001110011000101111011100",
35768 => "010000001000010001111010",
35769 => "010000111000101000011010",
35770 => "010000101011110010100010",
35771 => "010000100010011101100100",
35772 => "010001001111011110011010",
35773 => "010001011001011100101000",
35774 => "010000000110100011100100",
35775 => "001110111010010011100000",
35776 => "001110011101111101010010",
35777 => "001101110001110100110010",
35778 => "001100010110001110100110",
35779 => "001010111001001101000101",
35780 => "001010001000011111011110",
35781 => "001001101100011011000010",
35782 => "001001000010110100111001",
35783 => "001000010100011001001100",
35784 => "001000010111011110101100",
35785 => "001001100101011111111101",
35786 => "001010110100001011100111",
35787 => "001011010101001100111110",
35788 => "001011111110000000111110",
35789 => "001101000010100110000000",
35790 => "001101101011010010011100",
35791 => "001101011011101111111110",
35792 => "001100001101101110110100",
35793 => "001001010101100011100100",
35794 => "000101010010100101111011",
35795 => "000001010110000100001110",
35796 => "111100110101100001110100",
35797 => "110110010100001001101010",
35798 => "101101100100111001111110",
35799 => "100101011101101001100111",
35800 => "100001110111110011000001",
35801 => "100001100001101000010010",
35802 => "100010011101110101000111",
35803 => "100111000100011011001111",
35804 => "101110001000110000011110",
35805 => "110011110111110101100110",
35806 => "111001011001000111100101",
35807 => "000000000100100111100111",
35808 => "000110001101110100000010",
35809 => "001010110010001001100000",
35810 => "001101110000111111100010",
35811 => "001110101110111010100110",
35812 => "001100110101010111010010",
35813 => "000111111010100001000110",
35814 => "000001001001100100101111",
35815 => "111001101001001111111000",
35816 => "110001111100011011010010",
35817 => "101010111010111111100010",
35818 => "100101110010011110010011",
35819 => "100011110011101001000011",
35820 => "100100101011010011000111",
35821 => "100101100100010100000101",
35822 => "100101011111100110111000",
35823 => "100111000100111010111011",
35824 => "101011101000100101111100",
35825 => "110010001011001001100110",
35826 => "111001000011011000010101",
35827 => "111110111111111011010100",
35828 => "000101100011101010100111",
35829 => "001101110011100110010000",
35830 => "010101001001010010110110",
35831 => "011001101000010001001101",
35832 => "011011010111101010001000",
35833 => "011011011000011110010111",
35834 => "011010110110000000111011",
35835 => "011000110000000110001101",
35836 => "010011011010110100110110",
35837 => "001011000101100001001110",
35838 => "000010001001001011110010",
35839 => "111011011000001111011110",
35840 => "110110100011101110110011",
35841 => "110011000100100010101110",
35842 => "110010101100100010100100",
35843 => "110101100000100101101011",
35844 => "111001110101111110000100",
35845 => "111110011011100110001110",
35846 => "000001111100111001011111",
35847 => "000100011011001101001101",
35848 => "000110111110010010111110",
35849 => "001010000010001111111010",
35850 => "001101010011111011111000",
35851 => "010000010110101111001000",
35852 => "010011010010110010101100",
35853 => "010110000000111011101110",
35854 => "010111010011111001001010",
35855 => "010101100110010101001010",
35856 => "010000100001001111001000",
35857 => "001010000110011000010110",
35858 => "000011111011111101101010",
35859 => "111101010111010111001011",
35860 => "110110011011100110000000",
35861 => "110000100010110001101100",
35862 => "101100110011001111101010",
35863 => "101011100111001010100110",
35864 => "101100110111011101111110",
35865 => "110000001100110000110100",
35866 => "110100101010011000001100",
35867 => "111000111001011001001011",
35868 => "111011110000010001011101",
35869 => "111100110011000001010100",
35870 => "111100001010111111111010",
35871 => "111001010010010111110100",
35872 => "110100100000100000110101",
35873 => "110000010101001100100100",
35874 => "101110001100010011110110",
35875 => "101110100110100110110110",
35876 => "110001111101111010001000",
35877 => "110111001011000000100010",
35878 => "111101000101011110111110",
35879 => "000010111101100111010000",
35880 => "000111101001110101111100",
35881 => "001010000001011100000000",
35882 => "001001000010011000100110",
35883 => "000101010100110010111100",
35884 => "000000010000010000100111",
35885 => "111001111110000100001100",
35886 => "110011010110000101100100",
35887 => "101101101100101111111000",
35888 => "101001101111110001101110",
35889 => "101000000100000110001110",
35890 => "101000000100100110101010",
35891 => "101001101001111010001100",
35892 => "101101101001110011011100",
35893 => "110011000111011000000110",
35894 => "111000100101010111011000",
35895 => "111101100010010101000010",
35896 => "000001011101111110010100",
35897 => "000100010111111100111110",
35898 => "000110110000001011101001",
35899 => "001000111111111100101011",
35900 => "001010110101000011000010",
35901 => "001011011000010110000110",
35902 => "001010110100000000100100",
35903 => "001001110000100001001110",
35904 => "000111110011011111110000",
35905 => "000100111011000111100101",
35906 => "000010001100111101010100",
35907 => "111111111011000000011011",
35908 => "111101100001100011111000",
35909 => "111011001000011101010010",
35910 => "111000111011110100001101",
35911 => "110111010101111100011100",
35912 => "110111101111010000000001",
35913 => "111001111100100101001111",
35914 => "111011101100011001010110",
35915 => "111011111001101010011110",
35916 => "111011110101110000111101",
35917 => "111101000110010000110010",
35918 => "111111001110111001010010",
35919 => "000000111011011101111001",
35920 => "000010010001111101011000",
35921 => "000100000101010011100110",
35922 => "000111000111111000011010",
35923 => "001010110100001100001100",
35924 => "001101001110110111000010",
35925 => "001110100111001110101100",
35926 => "001111101110000111011010",
35927 => "001111001111000001000110",
35928 => "001100110000111101110110",
35929 => "001001011100111101111111",
35930 => "000110100010110001100001",
35931 => "000100110101000010011000",
35932 => "000011101010000000000011",
35933 => "000010001000001111101100",
35934 => "000000110001111101000101",
35935 => "000000111110011100001010",
35936 => "000010111101101011111000",
35937 => "000101111010011101110011",
35938 => "001001101010011000110001",
35939 => "001101101110101000110100",
35940 => "010001100000011001111100",
35941 => "010101010100011111000010",
35942 => "011000100011000001011011",
35943 => "011010100100010011000111",
35944 => "011011101010011111000000",
35945 => "011011101101001000100000",
35946 => "011011000000100010011011",
35947 => "011010000101110011101001",
35948 => "011001010110000010111001",
35949 => "011000110010110001101001",
35950 => "010111111001111110111110",
35951 => "010111010111100110110100",
35952 => "010110011000100100111110",
35953 => "010010001110100001110010",
35954 => "001011100010101010100110",
35955 => "000100100101010110100010",
35956 => "111101111011100000000111",
35957 => "110111100001110110010111",
35958 => "110001101110011111101000",
35959 => "101101101110111000111000",
35960 => "101011110011101000011000",
35961 => "101100001011011110100100",
35962 => "110000001110111111000110",
35963 => "110110110110110011110111",
35964 => "111101011011110011011110",
35965 => "000010111100010011011111",
35966 => "000111000110010100011011",
35967 => "001000100010001001000010",
35968 => "000101010001011010101101",
35969 => "111111001000101011100110",
35970 => "111000011111101100101100",
35971 => "101111100101100100100000",
35972 => "100110001111110111000001",
35973 => "100001101100100100101101",
35974 => "100001011111111111000000",
35975 => "100001110111111101011011",
35976 => "100001101101000111001101",
35977 => "100010001001101010111110",
35978 => "100011010010010101001110",
35979 => "100101010110011110101100",
35980 => "101001111000111010000010",
35981 => "101110111111000111111100",
35982 => "110001111100001100100010",
35983 => "110011101011010001101010",
35984 => "110101101001000000111100",
35985 => "111001101010110111011011",
35986 => "000000000000101110101010",
35987 => "000110001111101010011011",
35988 => "001100000100000101000100",
35989 => "010001001011010101101100",
35990 => "010011011000100010101010",
35991 => "010010001010101000100010",
35992 => "001110100101111011101110",
35993 => "001001010010101101101000",
35994 => "000010000111100101001101",
35995 => "111011001101011110010010",
35996 => "110111111001000011001100",
35997 => "110111010000101011011010",
35998 => "111000000001011110010100",
35999 => "111011000100001100010100",
36000 => "111111010111101001111101",
36001 => "000011101111011010101111",
36002 => "001000000001010111110110",
36003 => "001011110001110110001010",
36004 => "001111011101010110100000",
36005 => "010010111011000100111000",
36006 => "010100010000011100001110",
36007 => "010011010101111010110010",
36008 => "010011010010111010000000",
36009 => "010100111111111000111100",
36010 => "010101011100111111000110",
36011 => "010011110101000001010010",
36012 => "010001100011011110101000",
36013 => "001111010000111110011000",
36014 => "001101011111010110101100",
36015 => "001011000011010000010110",
36016 => "000101111101010101101111",
36017 => "111111000111000001110010",
36018 => "111001010100010011111001",
36019 => "110110100010010110001010",
36020 => "110110010000010101111110",
36021 => "110110111000110100010111",
36022 => "110111111001101011001111",
36023 => "111000111111001000110011",
36024 => "111001110001010101000101",
36025 => "111001101100011001101010",
36026 => "111000000100010111101000",
36027 => "110100111111111010111110",
36028 => "110000100010101100000010",
36029 => "101011100000000111000000",
36030 => "101000000111101101101010",
36031 => "100111010010001111111000",
36032 => "101000001101101010000100",
36033 => "101010010101011101111010",
36034 => "101101011101111000101100",
36035 => "110001011101111000101100",
36036 => "110101111001111000011001",
36037 => "111001111101111111010100",
36038 => "111100101110000001101101",
36039 => "111101001010000011011111",
36040 => "111010110001001110111100",
36041 => "110110101011101010010111",
36042 => "110010101011100110100010",
36043 => "101110111000101101011010",
36044 => "101010101110110010111100",
36045 => "100110111011000001011101",
36046 => "100101010010011001011101",
36047 => "100110010111011110101011",
36048 => "100111100100000001000000",
36049 => "101000011011101011001110",
36050 => "101100101000100110100110",
36051 => "110100001001111001010011",
36052 => "111100000000000101100100",
36053 => "000011110001101111110100",
36054 => "001011001110110100000111",
36055 => "010001011010010101000100",
36056 => "010101110001000000101110",
36057 => "010111010110110100111000",
36058 => "010110000011111000101010",
36059 => "010010110000000101110000",
36060 => "001110011000000110100000",
36061 => "001001110010100000110001",
36062 => "000101001001111111001000",
36063 => "000000100110110110011101",
36064 => "111101000011011100010110",
36065 => "111011011101000001011001",
36066 => "111100000011011000100010",
36067 => "111110010011011111000010",
36068 => "000000110111111010100010",
36069 => "000010011111000111010000",
36070 => "000011010101001101011110",
36071 => "000100000011010111011100",
36072 => "000100101101010101110001",
36073 => "000101011110001110110000",
36074 => "000101101110010111000000",
36075 => "000100111111110011000110",
36076 => "000100101110110000001011",
36077 => "000101100010011010111101",
36078 => "000110011101010110110101",
36079 => "000111010101010100100000",
36080 => "001000001000100100010111",
36081 => "001000010010101111110000",
36082 => "000111101101110001110101",
36083 => "000110001000100100100101",
36084 => "000010100111001100010101",
36085 => "111101101010101111110101",
36086 => "111001011101101000110011",
36087 => "110110100000101000100101",
36088 => "110011011101101001010010",
36089 => "110000010010001101011100",
36090 => "101110110001100010101000",
36091 => "101111111011111111111110",
36092 => "110010011110011100010000",
36093 => "110101000001111111011000",
36094 => "111000001111000101110010",
36095 => "111100101111101011110101",
36096 => "000001011100110010000011",
36097 => "000101001101110001111000",
36098 => "001000000000101100101011",
36099 => "001001110000011001111011",
36100 => "001010110010010111111100",
36101 => "001011111100111101000000",
36102 => "001101000110111101000010",
36103 => "001110001010100100011110",
36104 => "001111001100100101101110",
36105 => "001111110110111010100100",
36106 => "010001000001111001101110",
36107 => "010011000100000010011110",
36108 => "010100011111000011010110",
36109 => "010100110100111010111010",
36110 => "010101001100111000111010",
36111 => "010110000111101011000000",
36112 => "010101100001101111110110",
36113 => "010001111110110100100100",
36114 => "001101110100100110010010",
36115 => "001010010100100000011111",
36116 => "000110101101100010110001",
36117 => "000010111101101110111011",
36118 => "111110100110001011011001",
36119 => "111010101001011110101010",
36120 => "111001011111101100010000",
36121 => "111010101110110101111010",
36122 => "111100000110000001000110",
36123 => "111100011000011000111010",
36124 => "111100111110001011000101",
36125 => "111111001101101000100011",
36126 => "000001110011101111011101",
36127 => "000100000100011010101110",
36128 => "000110010110100011111000",
36129 => "001000010001110001000011",
36130 => "001001000100111010101000",
36131 => "000111111101011001010010",
36132 => "000110010101101000001101",
36133 => "000110000000001110101011",
36134 => "000101100000100100101011",
36135 => "000011011101110001110011",
36136 => "000000111110100010110001",
36137 => "111111001000000101000111",
36138 => "111100111110011001100100",
36139 => "111010000010000000011101",
36140 => "110111111111101111000101",
36141 => "110110110000100110010010",
36142 => "110101001110100010111000",
36143 => "110100000011100001000111",
36144 => "110010111001101010001010",
36145 => "110001110101110000110010",
36146 => "110001100100001111101010",
36147 => "110000110111110000101100",
36148 => "110000100011010100011110",
36149 => "110011100010001100011000",
36150 => "111001101001111101100010",
36151 => "111111111111100011000111",
36152 => "000101001000100011100000",
36153 => "001001110101111101011001",
36154 => "001101110000111100100110",
36155 => "010000000101011101000100",
36156 => "010000011100101101100110",
36157 => "001101011001100111101000",
36158 => "001000011011000110111000",
36159 => "000101011100000110000111",
36160 => "000100011101010111110011",
36161 => "000011111110110101000011",
36162 => "000011110100011111000101",
36163 => "000011100011010111101000",
36164 => "000011101000100111011001",
36165 => "000100100001011111101010",
36166 => "000100110100010110000010",
36167 => "000011101001110001010011",
36168 => "000010010111011101011000",
36169 => "000010011000010000100011",
36170 => "000011011011001100101101",
36171 => "000100011111000010001001",
36172 => "000101011010010111101000",
36173 => "000111010011000101111100",
36174 => "001010110111011110000100",
36175 => "001110111010111011111010",
36176 => "010001011011010011111110",
36177 => "010001100101100100001100",
36178 => "010000000001101000011110",
36179 => "001100011100100010111010",
36180 => "000101100100010100101010",
36181 => "111100110000110001111011",
36182 => "110101101011010101000011",
36183 => "110001111111111101011010",
36184 => "110000010110100111010100",
36185 => "101111001100001110011110",
36186 => "101111000000010010000100",
36187 => "110000001001001010110110",
36188 => "110010000001100101111000",
36189 => "110100011001010011110111",
36190 => "110101100101010010110010",
36191 => "110100010011000101010101",
36192 => "110010101010011111010110",
36193 => "110010011110100010011010",
36194 => "110010111010011010010000",
36195 => "110011010010011011001100",
36196 => "110100001101100111000101",
36197 => "110101110001100100110001",
36198 => "110111011010110101001101",
36199 => "111001001100011110011110",
36200 => "111001111110100011100101",
36201 => "110111111001100000110011",
36202 => "110011001110101101010010",
36203 => "101101011011000001000110",
36204 => "101000000110111111011010",
36205 => "100100101001100010011011",
36206 => "100011010110011111101111",
36207 => "100011101110011011111111",
36208 => "100100111001010101100111",
36209 => "101000000101101011001000",
36210 => "101111000001101100011010",
36211 => "110111111001011010000110",
36212 => "000000010001111100101110",
36213 => "000110100110000111011110",
36214 => "001001111011110111001001",
36215 => "001011010101101000110101",
36216 => "001010110110011010000000",
36217 => "001000001100100100101111",
36218 => "000100101001110100010000",
36219 => "000000101110111010000101",
36220 => "111101000011001100011100",
36221 => "111010100010111101100101",
36222 => "111001111100001100011010",
36223 => "111011111010101110000000",
36224 => "111111001000011100000001",
36225 => "000010010000010100110001",
36226 => "000101100010110110110110",
36227 => "001000101111000001000111",
36228 => "001011101101111010100011",
36229 => "001110001010011100101100",
36230 => "001111000101000000110110",
36231 => "001110100101110110100010",
36232 => "001101100100110101001110",
36233 => "001100100010001100110100",
36234 => "001011010011111101100000",
36235 => "001001101100110000010100",
36236 => "000111101110000000000110",
36237 => "000101011111011011011010",
36238 => "000011111001010101001000",
36239 => "000011010100010101101110",
36240 => "000011001011110000000010",
36241 => "000011010010001010100101",
36242 => "000011100111100111100001",
36243 => "000100001111101111101101",
36244 => "000100010001001011101101",
36245 => "000010110011101100110010",
36246 => "000000110111111011101110",
36247 => "111110110000001010010010",
36248 => "111100000010100100001100",
36249 => "111001010011001110100001",
36250 => "110110111101111110000111",
36251 => "110101110101000101110000",
36252 => "110101111110001100000100",
36253 => "110110010001000101110110",
36254 => "110110011110000100101110",
36255 => "110110111111000101111100",
36256 => "111000100101001111001010",
36257 => "111011011000010000000110",
36258 => "111110010100001010101001",
36259 => "000000111010110001101011",
36260 => "000010111100101010011100",
36261 => "000100101001100111111110",
36262 => "000110011101111100101100",
36263 => "000111011000010011101110",
36264 => "000111010011010001100001",
36265 => "000111100101001001111111",
36266 => "001000010010101110111010",
36267 => "001000011100101011101110",
36268 => "000111100100011010100000",
36269 => "000110001000001100000111",
36270 => "000100101101011101011101",
36271 => "000011101101110011110100",
36272 => "000010101011100001101111",
36273 => "000000010100001111011110",
36274 => "111101001011110001111110",
36275 => "111010010000110000101011",
36276 => "110110101000000011000000",
36277 => "110001010001001101010010",
36278 => "101010110100111011000010",
36279 => "100110100010101100111100",
36280 => "100110000010110111111001",
36281 => "100111100000011011111100",
36282 => "101100000110111011110100",
36283 => "110101011010000110010101",
36284 => "000000010011100101000011",
36285 => "001001111010110000000110",
36286 => "010001110000111111101100",
36287 => "011000001101100110011101",
36288 => "011100011100010111101000",
36289 => "011101000111010010111111",
36290 => "011011100011000110111101",
36291 => "011000001101000111010101",
36292 => "010010100001110000011100",
36293 => "001101000001000101001010",
36294 => "001000111110011111010100",
36295 => "000101101101011111110110",
36296 => "000100010100010100000100",
36297 => "000101010001111011010011",
36298 => "000110010000110100000001",
36299 => "000101001100111100001101",
36300 => "000011010111010011100110",
36301 => "000001110110000111111000",
36302 => "111111011110100010100111",
36303 => "111100101110101101110110",
36304 => "111010101001001001101101",
36305 => "111010010111000110111110",
36306 => "111110000001011011011111",
36307 => "000011101011010000010110",
36308 => "001000001100011000110100",
36309 => "001100110101110101100010",
36310 => "010001111110111001100000",
36311 => "010101010011010001111000",
36312 => "010101101110110011001010",
36313 => "010011101110010000111000",
36314 => "010000010100111110101100",
36315 => "001100101101010110110100",
36316 => "001001001011110000000011",
36317 => "000100101100011010111100",
36318 => "111110110010000100010011",
36319 => "111000101110011111010100",
36320 => "110011010001001001101010",
36321 => "101110111110010000110000",
36322 => "101100101001001111100110",
36323 => "101011111110010010100000",
36324 => "101101001010110001010000",
36325 => "101111100110110010100000",
36326 => "110000101000010100011110",
36327 => "110000111010010101010000",
36328 => "110100010110010100111010",
36329 => "111011100001110010100001",
36330 => "000010111001010000010101",
36331 => "001000000010000011100110",
36332 => "001100010010100110001110",
36333 => "010000011011111100101000",
36334 => "010010101001111110111100",
36335 => "010001111001111111010110",
36336 => "001101111111001000010000",
36337 => "000111100101000111000001",
36338 => "000001000110101011100100",
36339 => "111100001000111110010011",
36340 => "111000111101011111101100",
36341 => "110111000111001011101100",
36342 => "110101101100111011111001",
36343 => "110101000110100001100100",
36344 => "110101010100100110100101",
36345 => "110101011110011101000100",
36346 => "110101110111000001101000",
36347 => "110110011111000110001001",
36348 => "110110110101000011001100",
36349 => "110111001000100010001001",
36350 => "110111111000110000010110",
36351 => "111001011000000011100111",
36352 => "111011000110011111011101",
36353 => "111100110110100010000101",
36354 => "111110111100010011000110",
36355 => "000000101111101001100010",
36356 => "000010011001100001011010",
36357 => "000100100101100011011111",
36358 => "000110011110000001000100",
36359 => "000110100111110111111100",
36360 => "000100000111000111111111",
36361 => "000000000010111010000000",
36362 => "111100011100010101110100",
36363 => "111001001110001111001000",
36364 => "110101110111010111101110",
36365 => "110010011011110111000100",
36366 => "101111001000010101001010",
36367 => "101100110011111001010010",
36368 => "101100001001000010111100",
36369 => "101101101011001101011010",
36370 => "110001100100000101011000",
36371 => "110110111100101111101111",
36372 => "111100101000010001011101",
36373 => "000001010111111000110001",
36374 => "000101010101011010100010",
36375 => "001000011111000110010001",
36376 => "001000111110001010110010",
36377 => "000110111010110110100101",
36378 => "000100000010111010100000",
36379 => "000001000001100110000111",
36380 => "111110001100100100110110",
36381 => "111011010110111111011000",
36382 => "111001000001100100000000",
36383 => "111000101000110000110100",
36384 => "111010100111101001101110",
36385 => "111110010110111011110001",
36386 => "000010101000010010001110",
36387 => "000111000101010100110100",
36388 => "001011011001111000100101",
36389 => "001101111001000111100100",
36390 => "001110010110111110101000",
36391 => "001101010001001110110110",
36392 => "001010010000011111000110",
36393 => "000110011111011011000100",
36394 => "000011011110101110011101",
36395 => "000001100001011011101110",
36396 => "000000011111001101000100",
36397 => "000000011011100001110101",
36398 => "000001010110011111110011",
36399 => "000010110000100101110111",
36400 => "000101001010100111001110",
36401 => "001000101100000101100001",
36402 => "001011101100000010000000",
36403 => "001101100010010110010110",
36404 => "001101010110000111010000",
36405 => "001010000011001101100111",
36406 => "000101100110001010110000",
36407 => "000001111101101111110101",
36408 => "111110100110100101111000",
36409 => "111010101110110101100010",
36410 => "110111011011110110111010",
36411 => "110101111101101011101000",
36412 => "110101111101111001111111",
36413 => "110111111110100111010010",
36414 => "111011111010011101110110",
36415 => "111111101100010110010000",
36416 => "000011011001111011111010",
36417 => "000111011110100000100010",
36418 => "001010111011011110000110",
36419 => "001101100111111100001010",
36420 => "001110101011110010011100",
36421 => "001101011001100111011100",
36422 => "001010101001000001110110",
36423 => "000110111100011001101100",
36424 => "000010101110110101111111",
36425 => "111110111110101101011000",
36426 => "111100011101100001010111",
36427 => "111010100101101010101111",
36428 => "111001001011110000101111",
36429 => "111001101010110010001100",
36430 => "111011011111111011011111",
36431 => "111100110010000001000011",
36432 => "111011110000011011110001",
36433 => "110110100100101101001110",
36434 => "101110111110110010000110",
36435 => "101000011110000110000100",
36436 => "100100011101000111001001",
36437 => "100011010010011001100111",
36438 => "100011111011001010101011",
36439 => "100101000010100010000110",
36440 => "100101101101010110001110",
36441 => "100110110100101000011101",
36442 => "101100000000101100000000",
36443 => "110100011010001101001000",
36444 => "111011101100110000000010",
36445 => "000001001111100010101111",
36446 => "000101011001000010001100",
36447 => "001000111100001000110010",
36448 => "001100000111111000111010",
36449 => "001100100000111101001010",
36450 => "001010110110111110101111",
36451 => "001010001000001111111100",
36452 => "001010011000001010101001",
36453 => "001010011101111101011101",
36454 => "001001101000011001100000",
36455 => "001000100000000011110010",
36456 => "001000001111110000110111",
36457 => "000111110110000011100111",
36458 => "000101010100010010011011",
36459 => "000001100001000000111000",
36460 => "000000101101000010011101",
36461 => "000011111101110001000011",
36462 => "000111011001100101000100",
36463 => "001001011011110100111001",
36464 => "001010101101110100011000",
36465 => "001011010101000101111010",
36466 => "001100110111100010111000",
36467 => "001111110010000101110100",
36468 => "010001110010101111001010",
36469 => "010010101001001011110110",
36470 => "010100110110001101100000",
36471 => "011000100100001000000011",
36472 => "011010110101111000101101",
36473 => "011010010100000100111010",
36474 => "010111010111111010111100",
36475 => "010010011011000111010110",
36476 => "001100110001001110000010",
36477 => "000110101101010000101001",
36478 => "111111101100000011110101",
36479 => "111001100101100110101011",
36480 => "110110000111111100101101",
36481 => "110100001001110100011011",
36482 => "110010111101110100000010",
36483 => "110011110100110110011010",
36484 => "110111001100101001111100",
36485 => "111100000000001111000011",
36486 => "000000101101111101010101",
36487 => "000011011101001001000100",
36488 => "000011110001101110000001",
36489 => "000011000101000000011110",
36490 => "000001101111011101000000",
36491 => "111111101010000011111011",
36492 => "111101000101000011001100",
36493 => "111001001010111010101111",
36494 => "110100001111111110010010",
36495 => "110000111010001100011100",
36496 => "101111111111011100010010",
36497 => "110000010001010101110110",
36498 => "110001010110101000001110",
36499 => "110010010111011010000000",
36500 => "110010000000101100110100",
36501 => "110001100101111001001110",
36502 => "110010100111100110011100",
36503 => "110100001000100110011111",
36504 => "110101010111010011101010",
36505 => "110110101000011101111111",
36506 => "111000001100101001000111",
36507 => "111010001101000000111110",
36508 => "111100100111000011101011",
36509 => "111110110010010011110111",
36510 => "111111010100010010111100",
36511 => "111101100100100110100001",
36512 => "111010111011101111000101",
36513 => "111001001101010111010101",
36514 => "111000111000110101100110",
36515 => "111001000110101010001000",
36516 => "111001100100010100101100",
36517 => "111011001100001011001001",
36518 => "111110000101000010111111",
36519 => "000001101011000001010010",
36520 => "000101001110101110110001",
36521 => "000111010011011000110100",
36522 => "000111000111111010011001",
36523 => "000100111111011101101000",
36524 => "000001100111101101000000",
36525 => "111110010000101110101001",
36526 => "111011110000001110001100",
36527 => "111001111110001100101001",
36528 => "111000110101111000100000",
36529 => "111000110101010010110100",
36530 => "111010001010100000011111",
36531 => "111100100100111111001101",
36532 => "111111101100010001111111",
36533 => "000010011001000001001101",
36534 => "000011011011011010011001",
36535 => "000010100100111000011100",
36536 => "000000011101001000001000",
36537 => "111110010000110011100111",
36538 => "111100001100100001101000",
36539 => "111001110101011001100110",
36540 => "111000110000100111011110",
36541 => "111010010010101100000010",
36542 => "111101001000110101001010",
36543 => "000000000011010001100011",
36544 => "000011001111101010000110",
36545 => "000110100111101011100001",
36546 => "001000110100110101111110",
36547 => "001001010011110000010010",
36548 => "001000111101111111010010",
36549 => "000111111111001010111011",
36550 => "000101110000100101001111",
36551 => "000001011000111010010010",
36552 => "111011001101001110110010",
36553 => "110110100001110010111010",
36554 => "110100111101100011010010",
36555 => "110100001100010011011110",
36556 => "110011011101111001100010",
36557 => "110100011011010010100100",
36558 => "110111110100101111100110",
36559 => "111100111101010011010011",
36560 => "000010011001110111000111",
36561 => "000111100000110000101111",
36562 => "001100010001110100000010",
36563 => "001111101010011100101000",
36564 => "010000010100001101001110",
36565 => "001110000111100111100110",
36566 => "001010101011111010111111",
36567 => "000111111110110011100101",
36568 => "000101011111101000100111",
36569 => "000010001110000011100010",
36570 => "000000000010011110111011",
36571 => "000000011001111011100100",
36572 => "000010010110110011111001",
36573 => "000101000110111101101010",
36574 => "001000011001011000101001",
36575 => "001100011110111000101010",
36576 => "010001000000011011110100",
36577 => "010011101101101000100100",
36578 => "010100001011011011011000",
36579 => "010100000100101100010100",
36580 => "010011010110010101000100",
36581 => "010001010000100010000010",
36582 => "001110001000110010011000",
36583 => "001011000010100010001010",
36584 => "001000010011111101010110",
36585 => "000101000001011000111011",
36586 => "000001101001010001010111",
36587 => "111111010010110111000110",
36588 => "111100111100001001111000",
36589 => "111001101110010110010111",
36590 => "110110101000001001010110",
36591 => "110101000010001101100011",
36592 => "110101001000010011010010",
36593 => "110101101110011100001101",
36594 => "110110001010000100111101",
36595 => "110110000001010110000010",
36596 => "110100110011011011011001",
36597 => "110011010110101111101100",
36598 => "110010010001001010000100",
36599 => "110000111100010001100000",
36600 => "101111011010101011110000",
36601 => "101110100110101011110110",
36602 => "101111100101111011001010",
36603 => "110010011000100101111110",
36604 => "110101111000101001001001",
36605 => "111001100111001110001000",
36606 => "111101010010101101010000",
36607 => "000000110011111000011010",
36608 => "000100100000011111011011",
36609 => "000111000010010010011111",
36610 => "000110101001111110100000",
36611 => "000100011111010001000101",
36612 => "000010001011011010011100",
36613 => "111111100011000100001100",
36614 => "111100110110110010110010",
36615 => "111011011110101000000001",
36616 => "111100010000110001001110",
36617 => "111111000101101000101111",
36618 => "000010100101010101100000",
36619 => "000100111000101100000111",
36620 => "000110001101010011101100",
36621 => "000111100100001110100101",
36622 => "000111001000100111111100",
36623 => "000011100110010000110110",
36624 => "000000000101000010010110",
36625 => "111110111100110100100110",
36626 => "111111101000100000101101",
36627 => "000010011101100001010000",
36628 => "000110100110100111011010",
36629 => "001001101010011010110010",
36630 => "001100010101011011001010",
36631 => "001111111001110101110000",
36632 => "010010111010001101101110",
36633 => "010011111101111001101000",
36634 => "010010110111011000010010",
36635 => "001111110010111110100110",
36636 => "001011101001100001111000",
36637 => "000111010111101111100101",
36638 => "000011010011010100111000",
36639 => "000000100011101110001010",
36640 => "000000110010101101100111",
36641 => "000010111101110000000100",
36642 => "000100110010011010100100",
36643 => "000110001001111101010111",
36644 => "000110111110101111101100",
36645 => "000110010100111011000011",
36646 => "000100001100010110111000",
36647 => "000000111110000011000101",
36648 => "111101011001100001101111",
36649 => "111010110011011110001111",
36650 => "111001110110110111010111",
36651 => "111001111010100011111000",
36652 => "111010110001100100111110",
36653 => "111101110001000101011110",
36654 => "000010100001010000011011",
36655 => "000110100001100111101000",
36656 => "001000010100111001011000",
36657 => "000111100110110001100000",
36658 => "000101100010100100111011",
36659 => "000011100010000100010001",
36660 => "000000110110111111010110",
36661 => "111101110101001111100000",
36662 => "111011101110111011011001",
36663 => "111001011101010101111110",
36664 => "110110100000010101001110",
36665 => "110100110100011111000110",
36666 => "110101001000001110011000",
36667 => "110101011000011000000100",
36668 => "110011100001101110001110",
36669 => "101111111001000101100100",
36670 => "101100001111111011110110",
36671 => "101001111001010111011000",
36672 => "101001000001101101111000",
36673 => "101001101110010111000000",
36674 => "101100001000011100011110",
36675 => "101111100111100110110010",
36676 => "110100001111001000011110",
36677 => "111010011110110111001100",
36678 => "000001010010000111111001",
36679 => "000110111011110110011111",
36680 => "001010001001010110111010",
36681 => "001011000101101010101111",
36682 => "001010111100010001110101",
36683 => "001001010111100100101101",
36684 => "000101111100000000110100",
36685 => "000001010011000000010011",
36686 => "111100001011010110010000",
36687 => "110111011101001011110011",
36688 => "110011001101111001111100",
36689 => "101111111101001001000000",
36690 => "101110110000000010001010",
36691 => "101110110100001000001010",
36692 => "101111101110011000111000",
36693 => "110010001000010100100110",
36694 => "110101100111111100011010",
36695 => "111001011001101110010100",
36696 => "111100001110100010101001",
36697 => "111101101011101111110100",
36698 => "111111000110001111000101",
36699 => "000001011010111101111010",
36700 => "000100100110100000111011",
36701 => "000110111001010011001100",
36702 => "000110110101011001100100",
36703 => "000110010101111101011001",
36704 => "000110101000001010011000",
36705 => "000110001100100011010101",
36706 => "000101000000011110011111",
36707 => "000100011011001111101010",
36708 => "000100010001010001101110",
36709 => "000010110101110011110000",
36710 => "111111101000101101011000",
36711 => "111100001011001011110001",
36712 => "111001101001101100101000",
36713 => "111000010001100111010001",
36714 => "110111100001111101101111",
36715 => "110110011100001101110010",
36716 => "110101110110001011111001",
36717 => "110111101001100110101111",
36718 => "111011010011001010111101",
36719 => "111111001100011101000010",
36720 => "000011001110111010010111",
36721 => "000110111111001000010101",
36722 => "001001110001110000000000",
36723 => "001100100001100010101010",
36724 => "001111001101001110101000",
36725 => "010000001010110100001000",
36726 => "001111100001011101000100",
36727 => "001110010110111010111110",
36728 => "001100001000000010010100",
36729 => "001000000000101111001011",
36730 => "000010110111111110100010",
36731 => "111110100100101111011111",
36732 => "111100011000111011110111",
36733 => "111100100101001100110111",
36734 => "111110100101100010100000",
36735 => "000001011110111100000001",
36736 => "000100101111010001010010",
36737 => "001000001010001010101111",
36738 => "001011100111101111100100",
36739 => "001110011111100010001010",
36740 => "001111100001000111001100",
36741 => "001110101111101011010010",
36742 => "001101001111011101100000",
36743 => "001010100000101110110100",
36744 => "000101100111100100111111",
36745 => "111111100101110011001100",
36746 => "111010010100111110010101",
36747 => "110110101000100011000010",
36748 => "110101000000011111110011",
36749 => "110110010011001100101110",
36750 => "111010000000111100001010",
36751 => "111110111010011111011001",
36752 => "000100000110111111011100",
36753 => "000111101101001001010001",
36754 => "001000100000010110010010",
36755 => "000111001111000001010011",
36756 => "000011111101111010000001",
36757 => "111110100001101010100100",
36758 => "110111101010011110010100",
36759 => "110000010010011010110100",
36760 => "101001101000110011111000",
36761 => "100101001011111001000100",
36762 => "100100001010010001110111",
36763 => "100110011000011101110000",
36764 => "101010101100000000100010",
36765 => "110001100110100101111010",
36766 => "111010101000000111001010",
36767 => "000010011010111000011110",
36768 => "000111101101111110111100",
36769 => "001010110010110011011101",
36770 => "001010111101000011000100",
36771 => "001000110101111000000100",
36772 => "000101101011111100101010",
36773 => "000010011110111010001011",
36774 => "000000011100111110010011",
36775 => "111111000110011000110101",
36776 => "111101101111001011000101",
36777 => "111101001000111100111000",
36778 => "111101000010110011101011",
36779 => "111100001001001110110011",
36780 => "111010000010111111001010",
36781 => "110111100100100100011010",
36782 => "110101100100010100100001",
36783 => "110100010000111010010100",
36784 => "110100100000100100001010",
36785 => "110110010000001010001110",
36786 => "111000000110011011011011",
36787 => "111011010111010110010100",
36788 => "000000111101100101100001",
36789 => "000101101100000010110010",
36790 => "001000111000001110010110",
36791 => "001100101010010000000100",
36792 => "001111011011010111000010",
36793 => "001111000110011110001100",
36794 => "001100111000011110010010",
36795 => "001010010000001011110101",
36796 => "000111110111111111000011",
36797 => "000101101100100000010100",
36798 => "000010111111110111010000",
36799 => "000000100001100010101111",
36800 => "111111111111010001001000",
36801 => "000000110010001000110111",
36802 => "000000111100011110110101",
36803 => "000000101001101011010010",
36804 => "000000110010100101111110",
36805 => "000001000110011001101001",
36806 => "000010000100111001011011",
36807 => "000011101110100001010010",
36808 => "000100101111000010111010",
36809 => "000110001001100100000100",
36810 => "001001011010000000111110",
36811 => "001100110011101000000010",
36812 => "001111001000000000101110",
36813 => "010000111110101000011010",
36814 => "010010011011110110100110",
36815 => "010011000011001101111000",
36816 => "010010001110000001001000",
36817 => "001111110111101101110100",
36818 => "001100101110101101111110",
36819 => "001001000011100001001110",
36820 => "000101010110010010101100",
36821 => "000010101001101110111101",
36822 => "000001000011100111100101",
36823 => "000000001110111001001100",
36824 => "000000010101110000001100",
36825 => "000001011111111111001101",
36826 => "000011000010001000100101",
36827 => "000011101010011110001101",
36828 => "000011001000100100111110",
36829 => "000010001011100101111101",
36830 => "000001010000100110000000",
36831 => "000000100011011100101111",
36832 => "111111111000010100111010",
36833 => "111111011011011101010010",
36834 => "000000000010110011110100",
36835 => "000001010001110001001111",
36836 => "000010001101011000101011",
36837 => "000011000111000000110100",
36838 => "000100000110000000110111",
36839 => "000100111001111101100110",
36840 => "000101010001110001011011",
36841 => "000100101101110000110110",
36842 => "000011001011001001101111",
36843 => "000000000000010000101001",
36844 => "111001110001010010001000",
36845 => "110001010010000001100110",
36846 => "101001011100101000110110",
36847 => "100100001000010000000001",
36848 => "100001101010101110101111",
36849 => "100001100000100100001011",
36850 => "100010001011111110111101",
36851 => "100011010010101101001000",
36852 => "100110011011001011110110",
36853 => "101011110111000101000110",
36854 => "110001111000010110011010",
36855 => "110111111100010011100010",
36856 => "111101111111100100111101",
36857 => "000010111100000011010000",
36858 => "000110000000000010111101",
36859 => "000111001000000000011000",
36860 => "000110111000001000111011",
36861 => "000101011110011110001000",
36862 => "000010001101110000010011",
36863 => "111110011000111011001001",
36864 => "111100010011000100111011",
36865 => "111011011100100010011010",
36866 => "111010110000100111111111",
36867 => "111010000100110010111001",
36868 => "111001001110100100101000",
36869 => "111001010001000000100000",
36870 => "111010100000101100110000",
36871 => "111011100101111110100001",
36872 => "111100011101000010100100",
36873 => "111101010001000000000000",
36874 => "111101100111100100010010",
36875 => "111110010101000011000100",
36876 => "111111110101101011111101",
36877 => "000001111110001001011001",
36878 => "000101010000110001000001",
36879 => "001001010100110010101111",
36880 => "001101001010100010110000",
36881 => "010000110101110001111000",
36882 => "010100100110011100010010",
36883 => "011000001101111011011011",
36884 => "011010100111010100110101",
36885 => "011010000101000010010101",
36886 => "010110100001110001111000",
36887 => "010001100001010011011100",
36888 => "001011100011111000110001",
36889 => "000100101100100010001101",
36890 => "111110011111101011001000",
36891 => "111010010100110110000111",
36892 => "111000010111101010011111",
36893 => "111000111101111011100000",
36894 => "111011101100100010001000",
36895 => "111111010111111110011000",
36896 => "000011111111001101111000",
36897 => "001001011001111010000000",
36898 => "001110010010101011000010",
36899 => "010001010110010001110110",
36900 => "010001011011000000010100",
36901 => "001110001101010011100000",
36902 => "001000110010110100101101",
36903 => "000001111000010110111001",
36904 => "111001101111010111001001",
36905 => "110010010000001011100100",
36906 => "101110000010001011001100",
36907 => "101101001110011111001010",
36908 => "101110011000001000111110",
36909 => "110001101101010111010010",
36910 => "110111011000111110101011",
36911 => "111110000001110110010000",
36912 => "000100110000110110100110",
36913 => "001010000101010110000101",
36914 => "001011110100101011010010",
36915 => "001001111100110100100010",
36916 => "000101010000000010110011",
36917 => "111110110110011011101000",
36918 => "111000010011100101001000",
36919 => "110001000111101010011010",
36920 => "101001011011101100010100",
36921 => "100100011101000001001111",
36922 => "100100100000111011110011",
36923 => "101000111100100111001000",
36924 => "101111000110110011010110",
36925 => "110101011101010001000010",
36926 => "111100100110010001001110",
36927 => "000010111111000110110010",
36928 => "000110100011101100010111",
36929 => "001000011000011101000100",
36930 => "001001000100001001011000",
36931 => "001001000100101111001010",
36932 => "001001101011010001101000",
36933 => "001001000000001010110111",
36934 => "000101011110010110110011",
36935 => "000001011110101001101100",
36936 => "111110110001000000101111",
36937 => "111100011100101111111000",
36938 => "111001010100110011011110",
36939 => "110101111000010111011100",
36940 => "110011111110001001000010",
36941 => "110100010100101010100101",
36942 => "110110001111101111000100",
36943 => "111000000101010100100000",
36944 => "111000001110101010010111",
36945 => "110111011010101010000100",
36946 => "110111000010011010111110",
36947 => "110111110001010111100000",
36948 => "111010000110110011100011",
36949 => "111100010010110110000101",
36950 => "111100111110110011000000",
36951 => "111110011001101101110111",
36952 => "000001010001001100000101",
36953 => "000011011011011010111110",
36954 => "000100011000011101101111",
36955 => "000101000111100110100011",
36956 => "000101111101011000111110",
36957 => "000110000111010011000110",
36958 => "000100000110011101001000",
36959 => "111111100111101101001101",
36960 => "111010100100111100000110",
36961 => "110110110101010011101110",
36962 => "110100000110000000101000",
36963 => "110010001011010110111010",
36964 => "110010011110110010000000",
36965 => "110101010010000100001100",
36966 => "111001100011011011101000",
36967 => "111101111011000110101110",
36968 => "000000101001111001101000",
36969 => "000010010110001101101010",
36970 => "000100101110111110000000",
36971 => "000110110010011111000101",
36972 => "000111011101001000000100",
36973 => "000111101110110101100100",
36974 => "001000100010010110011110",
36975 => "001010000000001001111001",
36976 => "001011010101100000111100",
36977 => "001011111001001110110100",
36978 => "001100000000011010111100",
36979 => "001011101001001111111010",
36980 => "001010110000010011110010",
36981 => "001001010100101110110110",
36982 => "000111000110101111111000",
36983 => "000100111110001010111010",
36984 => "000011100011101010100001",
36985 => "000010011101000010111111",
36986 => "000010000101010101100111",
36987 => "000010110010001101000001",
36988 => "000100000100001010111110",
36989 => "000101101010100011100110",
36990 => "000111011010100010000111",
36991 => "001001000111001101010111",
36992 => "001010000000100101010010",
36993 => "001001001110000010100111",
36994 => "000111010010111100011110",
36995 => "000101001000001110101011",
36996 => "000011001111000011110011",
36997 => "000010011010100010101000",
36998 => "000010101000100000100010",
36999 => "000011010000001111010011",
37000 => "000011111101011111110001",
37001 => "000100001011110000100010",
37002 => "000011010111000100010001",
37003 => "000001001010001011100010",
37004 => "111101110000110011111111",
37005 => "111010001011000010110100",
37006 => "110110110000101101000001",
37007 => "110011100001101000111110",
37008 => "110001010001000000010010",
37009 => "110000001100100111110010",
37010 => "110000000000000100100100",
37011 => "110001010010110010010000",
37012 => "110100100101001101111110",
37013 => "111001000010000110011111",
37014 => "111101010110100110010010",
37015 => "000000110100001001001000",
37016 => "000010101010110111010011",
37017 => "000010001010011110001111",
37018 => "000000000101110010111011",
37019 => "111101011110111001010000",
37020 => "111001100000110001011100",
37021 => "110011111100010111111100",
37022 => "101110111000101111001000",
37023 => "101100010011110011011010",
37024 => "101100001111101110001000",
37025 => "101101101000010001000010",
37026 => "110000000000111010011010",
37027 => "110011101000001110001100",
37028 => "110111110010110111011100",
37029 => "111011110010010010111110",
37030 => "000000011111000011011010",
37031 => "000110010001111010000110",
37032 => "001011010101010010010010",
37033 => "001110010011011001010010",
37034 => "010000011000011011111110",
37035 => "010010110011101111100000",
37036 => "010100010101110110101000",
37037 => "010011010100011000000000",
37038 => "010000110010000001000000",
37039 => "001110110111110100101000",
37040 => "001101111000011011101000",
37041 => "001101010001100011000000",
37042 => "001100110100100001100010",
37043 => "001100000100111101010100",
37044 => "001011001101000010110111",
37045 => "001010101001001110011111",
37046 => "001010000101111010010000",
37047 => "001001110100001101001000",
37048 => "001010011001111000110000",
37049 => "001011010100011010101001",
37050 => "001011110110001101000011",
37051 => "001011110101110101111010",
37052 => "001011110011001101110010",
37053 => "001100100100010101110110",
37054 => "001110000001100111111010",
37055 => "001111011100010010110010",
37056 => "010000011001001011110000",
37057 => "010000110011000110100000",
37058 => "010000110010110101001010",
37059 => "001111100010000001001100",
37060 => "001100000000000111100110",
37061 => "000110110000101010000100",
37062 => "000000010000111011110010",
37063 => "111001000001001110111001",
37064 => "110010111111101000011110",
37065 => "101111101110100001100000",
37066 => "101111001111101001011100",
37067 => "110000100101110110001110",
37068 => "110011011110111100100010",
37069 => "111000111011001010010100",
37070 => "111111100011011100000110",
37071 => "000100111001011111010100",
37072 => "001001100011101110101010",
37073 => "001101011101101101101010",
37074 => "001110011010110111001100",
37075 => "001011101111000111011010",
37076 => "000110001101100010000010",
37077 => "111111000000111010001001",
37078 => "110101101100010111101010",
37079 => "101010010010011101110110",
37080 => "100010010100001110001101",
37081 => "100000111100111010110001",
37082 => "100001100100000011000001",
37083 => "100001011010011001111010",
37084 => "100001111111001010011001",
37085 => "100101001000000101001111",
37086 => "101100011110001011111010",
37087 => "110101101011101011001001",
37088 => "111101010111110100000001",
37089 => "000100100000101000110101",
37090 => "001011010010000111100010",
37091 => "010000000111111100000110",
37092 => "010010110011000000100000",
37093 => "010010010001010111100000",
37094 => "001110000111101110110000",
37095 => "000111110010111111000001",
37096 => "000000110000010001000110",
37097 => "111010111000111010101000",
37098 => "110110111010111111001101",
37099 => "110100000110101100010000",
37100 => "110010100011001100100110",
37101 => "110010010010011111111110",
37102 => "110100000100101100100001",
37103 => "111000001110011000000110",
37104 => "111011010110001010101001",
37105 => "111100000101011101011010",
37106 => "111101001001110110011101",
37107 => "111110101001111110010101",
37108 => "111111011110100110011011",
37109 => "000000000110100100001000",
37110 => "000000101000110010111110",
37111 => "000001110110010001001000",
37112 => "000011101111100011010111",
37113 => "000100010010111001010101",
37114 => "000011101110011111111001",
37115 => "000011110000110101110111",
37116 => "000011111001100111001111",
37117 => "000011000000011110000110",
37118 => "000000101000001100101101",
37119 => "111100011111101010001011",
37120 => "110111110001000111011100",
37121 => "110101000000101111111010",
37122 => "110100111010100111001101",
37123 => "110101010111000101111000",
37124 => "110101100001100010101111",
37125 => "110110111101010001000010",
37126 => "111010001001001011011100",
37127 => "111101110000010011101010",
37128 => "111111100100000101001010",
37129 => "111110011010010111101111",
37130 => "111100101100010001110111",
37131 => "111100110101101000001110",
37132 => "111101100111100001101001",
37133 => "111101100111100110011011",
37134 => "111101110010110111011010",
37135 => "111111010101001101010100",
37136 => "000001111111000100100010",
37137 => "000100100111110001101111",
37138 => "000110011100011110100100",
37139 => "000111010011011100101100",
37140 => "000111011100100111101111",
37141 => "000110101000101100110010",
37142 => "000011111111011110010100",
37143 => "000000011000100010100010",
37144 => "111101110000101000110011",
37145 => "111100000001000101101001",
37146 => "111010100010000101101010",
37147 => "111001101111111101011010",
37148 => "111001111110010010001110",
37149 => "111011001100010010000000",
37150 => "111100101010111110100111",
37151 => "111101011101001111100100",
37152 => "111101010101001001100010",
37153 => "111100000110010010101111",
37154 => "111010100010001101100000",
37155 => "111010001111011000101101",
37156 => "111011010011000000001110",
37157 => "111101000100101111010111",
37158 => "111111010110010011010011",
37159 => "000010001111100011110100",
37160 => "000110000001100010101010",
37161 => "001001001010011001100011",
37162 => "001001101010010110011111",
37163 => "001000000010011110111000",
37164 => "000101100000110101001110",
37165 => "000010011001001101001111",
37166 => "111110100000100011000100",
37167 => "111001101000110101001011",
37168 => "110100101101100101110001",
37169 => "110001000010100011111100",
37170 => "101111001101101111110000",
37171 => "101111100101000001100110",
37172 => "110001110001110110000000",
37173 => "110101010010011000011000",
37174 => "111001100001100011011001",
37175 => "111101000000100010000100",
37176 => "111111010010100010101111",
37177 => "000001011001111011010000",
37178 => "000011101100100111111100",
37179 => "000101100001100001001000",
37180 => "000110000100010100101000",
37181 => "000101110001000111101000",
37182 => "000101111001010111100001",
37183 => "000110010010010010101110",
37184 => "000110100010010100101111",
37185 => "000111000110101011101110",
37186 => "001000000010010011010011",
37187 => "001000111101110001000010",
37188 => "001001000010011000100110",
37189 => "001000010101000011101010",
37190 => "001000110000101011101000",
37191 => "001010001111100101010011",
37192 => "001010001111101100000110",
37193 => "001000010101111011101100",
37194 => "000111000010101010110000",
37195 => "000111111011000101000000",
37196 => "001000010110000000001100",
37197 => "000101001110111110000100",
37198 => "000000110100011100111101",
37199 => "111111001110111011101101",
37200 => "000001001000000111001100",
37201 => "000100001101101010001111",
37202 => "000110001010010111101010",
37203 => "000111011101110111100011",
37204 => "001010000001000110001000",
37205 => "001101001001111100101110",
37206 => "001110111110100110111000",
37207 => "001111101110100101001100",
37208 => "010001010110101111111110",
37209 => "010011111101110101100100",
37210 => "010100111011001010110010",
37211 => "010011000011011011111000",
37212 => "001111101000011001101100",
37213 => "001011100001100110011000",
37214 => "000110111010100100111001",
37215 => "000001101001111010000011",
37216 => "111100011100010001110000",
37217 => "111001001000000100011110",
37218 => "110111010000001011101101",
37219 => "110100101110001001001011",
37220 => "110001011010001010110110",
37221 => "101110011101111000110010",
37222 => "101101001001110100011100",
37223 => "101110010010111111111000",
37224 => "110001100100100000011110",
37225 => "110110001111110111000100",
37226 => "111011011101001110011001",
37227 => "000000001101110110110101",
37228 => "000100000000110101000101",
37229 => "000111011010011011111001",
37230 => "001011011111000100101111",
37231 => "001110111100010100100000",
37232 => "001111011101000100100010",
37233 => "001101110110101010010010",
37234 => "001100000011110010001010",
37235 => "001001110010101100110111",
37236 => "000101010010110101101110",
37237 => "111101111001000101101011",
37238 => "110110000110000010100110",
37239 => "110000001101111100111010",
37240 => "101011110001001001001110",
37241 => "101000001010101000011010",
37242 => "100101001010100101011001",
37243 => "100011101110001101000110",
37244 => "100101111011000010110101",
37245 => "101010111111101101100110",
37246 => "110001110110001000000010",
37247 => "111011000111010010000110",
37248 => "000101100000000110101111",
37249 => "001111100010011101011010",
37250 => "011000000010111011101001",
37251 => "011100101101100000010011",
37252 => "011101100001101001100001",
37253 => "011010111011010100111111",
37254 => "010100000011001000100110",
37255 => "001010110010110101011110",
37256 => "000010010000100110111001",
37257 => "111011111101001110011101",
37258 => "111000000010010010110101",
37259 => "110101010101011100110100",
37260 => "110011110101001011111000",
37261 => "110011110101111110101000",
37262 => "110100010100111111000100",
37263 => "110101110011011001100000",
37264 => "111000101001010000001100",
37265 => "111011000001111101111101",
37266 => "111100001010101111000000",
37267 => "111100000100010111110110",
37268 => "111011010001101110111100",
37269 => "111011111101101111011000",
37270 => "111110101011110011001111",
37271 => "000001111001001010101011",
37272 => "000101011010010100111101",
37273 => "001001111010000001100101",
37274 => "001110010010001000111000",
37275 => "010000011011010010111010",
37276 => "001111110010001110011100",
37277 => "001101001111101110010100",
37278 => "001001101101100111010110",
37279 => "000101101101011001000100",
37280 => "000000111001000111000010",
37281 => "111011111110000001110110",
37282 => "111001100111000100001011",
37283 => "111001111100011011100000",
37284 => "111010011000011101001100",
37285 => "111010011001010111011100",
37286 => "111010101101010001010001",
37287 => "111011000010110000110000",
37288 => "111011001100011111001000",
37289 => "111010101110001010111011",
37290 => "111001001010010010101100",
37291 => "111000001100011110000010",
37292 => "111001110111011011111100",
37293 => "111101010100011010110000",
37294 => "000001000110010011000110",
37295 => "000101010010110100010101",
37296 => "001001101000011000001100",
37297 => "001101100110010111100110",
37298 => "010000011000110111010110",
37299 => "001111111111011010001110",
37300 => "001100010000100111011110",
37301 => "000110100110101011101000",
37302 => "111110111011011111010100",
37303 => "110110010111111011110011",
37304 => "101111110000011000011100",
37305 => "101100000001000001110100",
37306 => "101010111000110011001000",
37307 => "101011101110011101001110",
37308 => "101101010100111010000110",
37309 => "101111100011101000110010",
37310 => "110010110100110000111110",
37311 => "110110010011010101000000",
37312 => "111000101011110110110100",
37313 => "111001101011111010010010",
37314 => "111001110010100010111100",
37315 => "111001100100100010101000",
37316 => "111001110101110110001000",
37317 => "111010101010111111001000",
37318 => "111011011011000111110111",
37319 => "111100011111001000011110",
37320 => "111101100101111100100001",
37321 => "111101001111100110011111",
37322 => "111011101101000000101110",
37323 => "111001110110101100110010",
37324 => "110111100000000100010100",
37325 => "110100111100111011111001",
37326 => "110010100010000100001110",
37327 => "101111110110100001110010",
37328 => "101101000011111110100110",
37329 => "101011010111001001001000",
37330 => "101011110010001111101100",
37331 => "101101110110000010110110",
37332 => "110001000000100001011000",
37333 => "110101101101011010000000",
37334 => "111011010111011111100011",
37335 => "000000010101101110110000",
37336 => "000011100000011101010111",
37337 => "000101011010001011000110",
37338 => "000111100010001101100000",
37339 => "001001011011101101000001",
37340 => "001010010100111000001001",
37341 => "001011001111101010001001",
37342 => "001011111001011101000010",
37343 => "001011100101101101110100",
37344 => "001011011000100011011000",
37345 => "001011011010100111100001",
37346 => "001011000100011001000110",
37347 => "001010100001100110110000",
37348 => "001010011011111000100001",
37349 => "001011100000111001011000",
37350 => "001100111111100100000000",
37351 => "001101110111010000000000",
37352 => "001110101010100101011010",
37353 => "001111101010100111000110",
37354 => "010000110001010000011110",
37355 => "010001110111111110000110",
37356 => "010010110001000000011110",
37357 => "010100000011010100100000",
37358 => "010101100011000111010010",
37359 => "010110011111001010010110",
37360 => "010111000101010001000110",
37361 => "010111000101101001001010",
37362 => "010110101111100101110000",
37363 => "010110100110011101010010",
37364 => "010101111001001010111010",
37365 => "010101001001110000010000",
37366 => "010100111100111010000100",
37367 => "010011101010000100110110",
37368 => "010000100110010100100010",
37369 => "001100001101110100111100",
37370 => "000111000100100100010010",
37371 => "000001111011110001110000",
37372 => "111100100000011010000010",
37373 => "110110111001111100101000",
37374 => "110001101101011001110110",
37375 => "101100110111010001111110",
37376 => "101001011001100000111110",
37377 => "101000000101010010001100",
37378 => "101000100010010000010010",
37379 => "101001111100011000000010",
37380 => "101010010111111001011000",
37381 => "101010010101110101000100",
37382 => "101100101001011001011110",
37383 => "110001001110110101100010",
37384 => "110111000110101110000010",
37385 => "111101011000111001000110",
37386 => "000010000010111111010110",
37387 => "000100101111110011010001",
37388 => "000110010001100001100010",
37389 => "000110110111010010000111",
37390 => "000110010010000110110010",
37391 => "000011010110000110101111",
37392 => "111110011110001001000011",
37393 => "111001010011100010000110",
37394 => "110100110111111011011100",
37395 => "110010111111000110000010",
37396 => "110010101111100100100110",
37397 => "110001000010111000110110",
37398 => "101111001011001110110110",
37399 => "101111101110101000011010",
37400 => "110010001110101010100100",
37401 => "110100011111000110001011",
37402 => "110100011100011000000000",
37403 => "110011100111100110001010",
37404 => "110100101101100100100000",
37405 => "110111001010100001110000",
37406 => "111010100010111010001100",
37407 => "111111110000100101011100",
37408 => "000111001010100011011011",
37409 => "001111100100000000111010",
37410 => "010101100011111010111010",
37411 => "011000101001000100101001",
37412 => "011011000000011111111111",
37413 => "011010101101001001111001",
37414 => "010101110000010000011100",
37415 => "001110100011111010101010",
37416 => "000111001001011100100010",
37417 => "000000100010101011001110",
37418 => "111100001000010111100100",
37419 => "111010001110111111010101",
37420 => "111010010110111100011101",
37421 => "111011111010000100101000",
37422 => "111110000000000101100110",
37423 => "111111011100101011000111",
37424 => "000000101010010000000101",
37425 => "000011001111100100111000",
37426 => "000101010011101100011100",
37427 => "000100000110111000110001",
37428 => "000001000001001101001110",
37429 => "111101110001100011100111",
37430 => "111011011001100101111101",
37431 => "111011000011101100110010",
37432 => "111011010101001011000000",
37433 => "111100000010000001100101",
37434 => "111111001100001110110000",
37435 => "000010011000000110011111",
37436 => "000001111101010111010001",
37437 => "111111010010000110111110",
37438 => "111100101111001100010001",
37439 => "111010110110110011100010",
37440 => "111001110000011000000100",
37441 => "111001000001010010110011",
37442 => "111000011000101111010010",
37443 => "111000111000110111111100",
37444 => "111010110011100000001101",
37445 => "111100010001001011111110",
37446 => "111100001110010001011010",
37447 => "111011101011111100000110",
37448 => "111011000110110100100000",
37449 => "111010000101110011101010",
37450 => "111000100001010010110000",
37451 => "110110010111011111111001",
37452 => "110100110110110011110010",
37453 => "110101110111111011010110",
37454 => "111001001101111010110100",
37455 => "111101110011011101001011",
37456 => "000011011110001001110111",
37457 => "001001010011101101100000",
37458 => "001101110110100001100000",
37459 => "010000100101011101110110",
37460 => "010000110111011101111100",
37461 => "001110001111000110001110",
37462 => "001001100111010111000001",
37463 => "000011101110011111001011",
37464 => "111101001101101000000110",
37465 => "110111110011101100100110",
37466 => "110100010010111111001010",
37467 => "110010100100011000011010",
37468 => "110011000100101101010100",
37469 => "110101000100100000001000",
37470 => "110111010100011101100100",
37471 => "111010000110100101111011",
37472 => "111101011000011100000100",
37473 => "000000001010011001110001",
37474 => "000001110010010101001000",
37475 => "000001111101001000011100",
37476 => "000001001001001010011111",
37477 => "000000011101111000111100",
37478 => "000000001001011111111001",
37479 => "111111010000010011011010",
37480 => "111101100010111110011000",
37481 => "111100010000000101110101",
37482 => "111011101001000100111010",
37483 => "111010011100011010000011",
37484 => "111000011001100010011010",
37485 => "110110010000001000001110",
37486 => "110100011000101011011111",
37487 => "110010100111100110000100",
37488 => "110000001011010010100110",
37489 => "101101001011011110100110",
37490 => "101011000100110000010010",
37491 => "101010101101010100000110",
37492 => "101100001010100101111100",
37493 => "101111010000101111101110",
37494 => "110011000111010110111000",
37495 => "110110111010010100011100",
37496 => "111010110011110111111011",
37497 => "111111001000100100100111",
37498 => "000011000100101001101111",
37499 => "000101100111110111100101",
37500 => "000111000111110011100110",
37501 => "001000000011101000110011",
37502 => "001000011000111101010010",
37503 => "001000010001001100001100",
37504 => "000111100001100010001000",
37505 => "000110100001010101101010",
37506 => "000110011011110111000100",
37507 => "000111001001110010011101",
37508 => "001000001110000011010101",
37509 => "001001111011000001111000",
37510 => "001011110001111011100000",
37511 => "001101101000110111001110",
37512 => "010000001000010101001110",
37513 => "010010110100011100111100",
37514 => "010100101110001110011000",
37515 => "010101011100111000100110",
37516 => "010110011001000111111100",
37517 => "011001101000110111110000",
37518 => "011101001100111000011100",
37519 => "011101101110000111011001",
37520 => "011100110010000101011100",
37521 => "011100011101010101011001",
37522 => "011011111001000010111011",
37523 => "011011000101110011011011",
37524 => "011001010011111110001110",
37525 => "010100110001010000111110",
37526 => "001111100010010010110010",
37527 => "001100011100110110101000",
37528 => "001010010010111111001010",
37529 => "000111000011111101011010",
37530 => "000011011100000011100000",
37531 => "000001110100010000101111",
37532 => "000010000111011101111011",
37533 => "000001100000001001010010",
37534 => "000000010110111010101100",
37535 => "000000111000001011011101",
37536 => "000001100101000000000110",
37537 => "000000101000101010011001",
37538 => "111110010010000010011100",
37539 => "111011011110101111001001",
37540 => "111001100101101000001010",
37541 => "110111110111001101010000",
37542 => "110101101011000110100100",
37543 => "110101000101000000000001",
37544 => "110101100011111101110000",
37545 => "110101001111001000011111",
37546 => "110101001001000110111110",
37547 => "110101010101001100101011",
37548 => "110100101011010100111100",
37549 => "110011100111101010111110",
37550 => "110010011100001000101010",
37551 => "110000111110101001011110",
37552 => "101111001110111000001000",
37553 => "101101111000111000111110",
37554 => "101110011011001110000010",
37555 => "110000100111110010110110",
37556 => "110011100001000100011110",
37557 => "110111001100000110010101",
37558 => "111010110110111111000111",
37559 => "111101111110001101000011",
37560 => "000000110110110001101010",
37561 => "000010010010101000011000",
37562 => "000000111000100001110110",
37563 => "111101000110001111000010",
37564 => "111000110000000001101111",
37565 => "110101101111100101011011",
37566 => "110100011100101011111100",
37567 => "110100101001111011111000",
37568 => "110110101001100111011100",
37569 => "111010011100101110010010",
37570 => "111111111001001010011110",
37571 => "000101100011010000011011",
37572 => "001001011000111100110011",
37573 => "001011100000000110010111",
37574 => "001100010000010100100110",
37575 => "001011011110110101000011",
37576 => "001010010100000111000001",
37577 => "001001001111011000011110",
37578 => "000111010110011010000100",
37579 => "000101000100111100100101",
37580 => "000100100010000011010010",
37581 => "000110000110101100001011",
37582 => "000111011111100010001111",
37583 => "001000001000001000001010",
37584 => "001001000110010001110100",
37585 => "001001010011110100101110",
37586 => "000111111000010000010110",
37587 => "000101011001001011111100",
37588 => "000010000000100000000010",
37589 => "111110110011001110000001",
37590 => "111100111000001110000100",
37591 => "111011011111101010011000",
37592 => "111010001000001111111100",
37593 => "111001100100000101010010",
37594 => "111010010101100011101011",
37595 => "111011100110010101101010",
37596 => "111100001000010001010101",
37597 => "111011100110010000110001",
37598 => "111010010101001001001100",
37599 => "111001011111100010101000",
37600 => "111001111011101000011111",
37601 => "111010110000010111000101",
37602 => "111011010000111000010111",
37603 => "111011101110110111111001",
37604 => "111100010111011101111000",
37605 => "111101011010101100110110",
37606 => "111110001101010101011100",
37607 => "111100111101000111111001",
37608 => "111001011110100001101001",
37609 => "110101101010100011100000",
37610 => "110010011010111010101110",
37611 => "101110110010000011101110",
37612 => "101010011111000000100100",
37613 => "100111010010111010101000",
37614 => "100111010111100110101001",
37615 => "101010110111001101011100",
37616 => "110000010101010110010000",
37617 => "110111001100010110000011",
37618 => "111111001001000101011000",
37619 => "000110110000001100010011",
37620 => "001100100110111100111110",
37621 => "001111110000011100010000",
37622 => "001111111001100111000010",
37623 => "001101110010011101101010",
37624 => "001010001010111100111000",
37625 => "000101100101010010110110",
37626 => "000000101001001110011011",
37627 => "111100000000010010010000",
37628 => "111000110110011111000001",
37629 => "111000001010101110110111",
37630 => "111001011101111100100000",
37631 => "111011011111010100100011",
37632 => "111101110000011000011111",
37633 => "000000101001100011011100",
37634 => "000011111101011101100111",
37635 => "000110011110101100010010",
37636 => "000111001100010011101110",
37637 => "000110001010100010011000",
37638 => "000100000110101101100100",
37639 => "000001011111001000110110",
37640 => "111110011000100011000010",
37641 => "111010110011010100101010",
37642 => "110111101100110100011011",
37643 => "110110100001000010001000",
37644 => "110110110100010101100100",
37645 => "110111100101011000111101",
37646 => "111001000001000001001100",
37647 => "111010110100100011111000",
37648 => "111100001111100111011101",
37649 => "111100110101010000011100",
37650 => "111100010101101111000010",
37651 => "111011000101110001101011",
37652 => "111001000000110000100101",
37653 => "110110001001010100000011",
37654 => "110011100111111011001100",
37655 => "110010011100110111000010",
37656 => "110010110111001000101000",
37657 => "110011110100101100101010",
37658 => "110100101100011000000100",
37659 => "110110100010010000110111",
37660 => "111000111011101111100000",
37661 => "111010011101100011100010",
37662 => "111011010000111011111110",
37663 => "111011111010010000011010",
37664 => "111100101110010011110111",
37665 => "111101000101010001111111",
37666 => "111100100011001100100100",
37667 => "111100100100010111001101",
37668 => "111101101011001101110011",
37669 => "111111011001000111010111",
37670 => "000001111000110101111110",
37671 => "000100101100111111100001",
37672 => "000111011101100000110010",
37673 => "001010000011100100111001",
37674 => "001011110111001101111100",
37675 => "001101000001000011110010",
37676 => "001110001010010110010000",
37677 => "001111010100110100000000",
37678 => "001111110101010011111110",
37679 => "001111101011101110110100",
37680 => "010000010101110000111110",
37681 => "010001010110100001000100",
37682 => "010000011111010011110100",
37683 => "001110100000100101011100",
37684 => "001101100001011001011000",
37685 => "001101101001001010010100",
37686 => "001110010100001111111010",
37687 => "001110110001000011000010",
37688 => "001110110110110101111010",
37689 => "001111100000110010101100",
37690 => "001111101101111111101100",
37691 => "001110010101110110011110",
37692 => "001101010000101101000110",
37693 => "001101011011110001101010",
37694 => "001101100000110100000100",
37695 => "001100110000101011100010",
37696 => "001011011100000111010100",
37697 => "001010001001000100101111",
37698 => "001000001001010011111100",
37699 => "000100010000011101111000",
37700 => "111111100101101000111110",
37701 => "111100000101111010000001",
37702 => "111011000001000101100001",
37703 => "111011111011000001001100",
37704 => "111101010110001000011000",
37705 => "111111110001001001011111",
37706 => "000010101011100001010110",
37707 => "000100010101010110011010",
37708 => "000101110000011011100010",
37709 => "000111101010101110000101",
37710 => "001001100011101011001001",
37711 => "001010100000101101100011",
37712 => "001000110111010011011010",
37713 => "000110011100011101110000",
37714 => "000101011011010001100101",
37715 => "000100101111000010100110",
37716 => "000100100011100110111001",
37717 => "000101000110010110111110",
37718 => "000110111011010000010010",
37719 => "001011001110011100110000",
37720 => "001101111110111100001110",
37721 => "001011011000111011100101",
37722 => "000101111101110011000100",
37723 => "000000111001011000100011",
37724 => "111100100010010111011011",
37725 => "110111010100101101001000",
37726 => "110001001011111111001000",
37727 => "101100010101111101100010",
37728 => "101001011011010101101110",
37729 => "101000110011111001110110",
37730 => "101011011010111010001000",
37731 => "110000010110111000001100",
37732 => "110110011101010101111111",
37733 => "111100100101001101100011",
37734 => "000001100000010000000101",
37735 => "000101101000000000100011",
37736 => "001001101111000100100011",
37737 => "001101101111011110100100",
37738 => "010000111011011001001100",
37739 => "010010011101100101001010",
37740 => "010010000010011001101000",
37741 => "001111111100001110001100",
37742 => "001101101000010110010110",
37743 => "001100000110101010011000",
37744 => "001001011110011100000100",
37745 => "000011111100100000100101",
37746 => "111100100000001011011101",
37747 => "110101000101101111001000",
37748 => "101111011110000001000000",
37749 => "101011111110010111000000",
37750 => "101000110011110011101100",
37751 => "100101110011000010100011",
37752 => "100101101000000110110010",
37753 => "101001100000111001000100",
37754 => "101111100001110000101000",
37755 => "110101000100001011011001",
37756 => "111001011111111010111010",
37757 => "111110001011101110000100",
37758 => "000011110000000011110101",
37759 => "001001010000010101000000",
37760 => "001101001010100010110000",
37761 => "001110101000000010110110",
37762 => "001110011010010011011110",
37763 => "001100111111101010100100",
37764 => "001010000000000110011100",
37765 => "000101011100111001010111",
37766 => "111111011010110011010001",
37767 => "111001001010111110001101",
37768 => "110011111001100010010110",
37769 => "101110110110010011011010",
37770 => "101010001110101110100100",
37771 => "100110101111101011111011",
37772 => "100100011111100001011011",
37773 => "100100011111100100001001",
37774 => "100110111010011100101010",
37775 => "101011010111001100101010",
37776 => "110010000011010001101110",
37777 => "111010011101111000110110",
37778 => "000011011011111111010111",
37779 => "001010110011111111000100",
37780 => "001111101100100011000110",
37781 => "010011100001111111011110",
37782 => "010101111001011101000010",
37783 => "010101010000000010001100",
37784 => "010001000110100000111110",
37785 => "001001111100001011101101",
37786 => "000010001001100111110000",
37787 => "111010111011000111100111",
37788 => "110011111011111111010010",
37789 => "101110011010001100001110",
37790 => "101011000100110111110100",
37791 => "101010010000010011111000",
37792 => "101100100100011000011100",
37793 => "110001001001000110010010",
37794 => "110110111111110111100001",
37795 => "111101000001000010101011",
37796 => "000001100001110011110101",
37797 => "000100011100101001011101",
37798 => "000110000110011110000101",
37799 => "000110000101100000001000",
37800 => "000100011110010001111100",
37801 => "000001011000100000000101",
37802 => "111101000100000001010010",
37803 => "111001000011111011000100",
37804 => "110111001010111101111010",
37805 => "110111100001111000101100",
37806 => "111001001001111011000000",
37807 => "111011010100001110111010",
37808 => "111101101010000111010101",
37809 => "000000000000111010011101",
37810 => "000001111010011010000101",
37811 => "000010011001011010011100",
37812 => "000000110001100011100011",
37813 => "111101011001000111010001",
37814 => "111001010111101001011001",
37815 => "110101011110010011010010",
37816 => "110010011100011111011100",
37817 => "110000101110110001001000",
37818 => "101111011101101101111010",
37819 => "101110101101111011100110",
37820 => "101111101010001001001110",
37821 => "110001111110011110100100",
37822 => "110101000011100110001100",
37823 => "111000110100000011011001",
37824 => "111100111000111110001001",
37825 => "000000100100100111001011",
37826 => "000010101111010010111000",
37827 => "000011101110111010011010",
37828 => "000101000111001101111011",
37829 => "000110101111011101110010",
37830 => "000111101100110000000011",
37831 => "001000001001011111110110",
37832 => "001000100100011100010010",
37833 => "001000010000001011111100",
37834 => "000110001011001111010100",
37835 => "000011101000001100110111",
37836 => "000010010110101000100000",
37837 => "000010000000110100011101",
37838 => "000001111011001001010111",
37839 => "000001101010011001001011",
37840 => "000001000010011000100101",
37841 => "000000011110100100000010",
37842 => "000000001110111001011100",
37843 => "000000100100011011000101",
37844 => "000001011111110101111000",
37845 => "000010101110000110000100",
37846 => "000100110010111010010010",
37847 => "000111111010110011000000",
37848 => "001010110011111101111110",
37849 => "001100001111000111010000",
37850 => "001100011000110101111110",
37851 => "001100010010101110101110",
37852 => "001011110100010010100101",
37853 => "001010001111000001011011",
37854 => "001000000010011111101110",
37855 => "000110000010010000010010",
37856 => "000100010000101001001101",
37857 => "000001110011010011110001",
37858 => "111101101011101100010011",
37859 => "111000110111011011001110",
37860 => "110101001110000010011000",
37861 => "110011011000101100111110",
37862 => "110011100000101000011000",
37863 => "110101110100010100000010",
37864 => "111010000001101100011000",
37865 => "111110111100110101001100",
37866 => "000011001011000110001010",
37867 => "000110111000110001010100",
37868 => "001011001010111000010100",
37869 => "001111101000001011000100",
37870 => "010010111000101110100000",
37871 => "010100000000001110110000",
37872 => "010011011101010110001000",
37873 => "010010111111000000001000",
37874 => "010010101101001101011100",
37875 => "010001010001101010111010",
37876 => "001111001000001001000010",
37877 => "001101101111110101101010",
37878 => "001101101011111100100110",
37879 => "001110100010111011110100",
37880 => "001111001101100010110100",
37881 => "001110111100011011111000",
37882 => "001101011010100000001000",
37883 => "001001101001010100001111",
37884 => "000011101111100001100110",
37885 => "111110010111101011100110",
37886 => "111011011111001001010110",
37887 => "111001101010011100100000",
37888 => "110111010111000000010001",
37889 => "110101101101000010110010",
37890 => "110110100101001111000100",
37891 => "111010000111011100100001",
37892 => "111101101010100010001110",
37893 => "111111110101101111100111",
37894 => "000011010111000100010100",
37895 => "001000011001001001000001",
37896 => "001011110100110101110010",
37897 => "001101101011100010101010",
37898 => "001110011010101111110010",
37899 => "001101001010000101110010",
37900 => "001010100011100101101100",
37901 => "000110111111001011110101",
37902 => "000010101011111101111010",
37903 => "111110010101110010000010",
37904 => "111001010100000001001000",
37905 => "110011011111101001101100",
37906 => "101101110010111011001100",
37907 => "101000111010011010001000",
37908 => "100101110001100000001111",
37909 => "100101000000111000011011",
37910 => "100110101001101111101011",
37911 => "101001010001011001001110",
37912 => "101011001101110000111000",
37913 => "101101110001011011010100",
37914 => "110010000100010111000110",
37915 => "110111000001110111101110",
37916 => "111100001111110011011100",
37917 => "000000110100100110110100",
37918 => "000100100010101111011000",
37919 => "001001110011000001010110",
37920 => "001111110101000011001010",
37921 => "010010001011101011011110",
37922 => "001111100111111101010100",
37923 => "001011011000000001100011",
37924 => "001000010111110011011001",
37925 => "000101011110001110010100",
37926 => "000000000100000100010100",
37927 => "111001000010110111111100",
37928 => "110011101011010000001110",
37929 => "110001011100101101110110",
37930 => "110000110011011111111100",
37931 => "110000010011111001011000",
37932 => "110001010100011001000010",
37933 => "110100101000000010011111",
37934 => "111001011110010001010111",
37935 => "111111011100110101101101",
37936 => "000101000000000100010001",
37937 => "001001001101011011001101",
37938 => "001101000010111100111010",
37939 => "001111111101001011000010",
37940 => "010001010101010110111100",
37941 => "010010010001011001011100",
37942 => "010011011110100111100110",
37943 => "010100110101010000101110",
37944 => "010101000101000011100110",
37945 => "010010111100011111001010",
37946 => "001110111100111100011000",
37947 => "001010010011001000001100",
37948 => "000101011110110001111001",
37949 => "000000000000100001010110",
37950 => "111010001010010100100111",
37951 => "110101101011110111111110",
37952 => "110011011101011011011000",
37953 => "110011101110111011100010",
37954 => "110110001100000111001100",
37955 => "111001011000101010010000",
37956 => "111101000000101110111100",
37957 => "000001000101010111100001",
37958 => "000100100110101100101111",
37959 => "000110110001101010011001",
37960 => "000110100000001100010100",
37961 => "000011011011011011100100",
37962 => "111111000100001010001001",
37963 => "111010101010100001011100",
37964 => "110110100000010000010100",
37965 => "110011000110010101101000",
37966 => "110001011000110111110110",
37967 => "110001010110001111111000",
37968 => "110010011000001110000000",
37969 => "110100111010001001110100",
37970 => "111000011001101011111000",
37971 => "111011001001111101011110",
37972 => "111100011101011011010101",
37973 => "111011001101111001000001",
37974 => "110110110011110011011111",
37975 => "110001011011100010100000",
37976 => "101101011000101011001100",
37977 => "101010101001110100101000",
37978 => "101000010100111110101010",
37979 => "100110110100011000010011",
37980 => "100111100110010000010001",
37981 => "101010111010100110001000",
37982 => "101111110101011110111000",
37983 => "110101111000111011111011",
37984 => "111100101100111010001101",
37985 => "000010111111101111010000",
37986 => "000111011001000011110011",
37987 => "001001110001111001011011",
37988 => "001011001111011000101111",
37989 => "001100001111110100110110",
37990 => "001011100010010011011011",
37991 => "001000110000110010111100",
37992 => "000101111111001100000011",
37993 => "000100001010110010001111",
37994 => "000010011100000001010101",
37995 => "000000001001110010110101",
37996 => "111101011101010100011000",
37997 => "111100001111100010011011",
37998 => "111101111000110010101011",
37999 => "000000111000010111100010",
38000 => "000011101000010100100110",
38001 => "000101111001100110011111",
38002 => "001000010100001011101100",
38003 => "001011010101010111011100",
38004 => "001110000000111001001000",
38005 => "001111111001011001110100",
38006 => "010001010010010000111000",
38007 => "010001111000000000111100",
38008 => "010001001001001110110010",
38009 => "001110010001100110111110",
38010 => "001001101000000011100001",
38011 => "000101000010100011100100",
38012 => "000001011001010011111100",
38013 => "111110100011111100001100",
38014 => "111100000110000110111001",
38015 => "111010001100001111001100",
38016 => "111001100110010000101101",
38017 => "111001011000010001001011",
38018 => "111000000010111110111111",
38019 => "110101010110101100101110",
38020 => "110010001000111100011110",
38021 => "101111110101010000000110",
38022 => "101110110001011101111110",
38023 => "101111011001001000111110",
38024 => "110010101100111011101000",
38025 => "110110111101000111001101",
38026 => "111001101010010101010000",
38027 => "111011101011101001100111",
38028 => "111111001010001101000111",
38029 => "000011110110010000001100",
38030 => "000111011100011111101100",
38031 => "001000111011110011100010",
38032 => "001001001010010111110010",
38033 => "001000110111100111100110",
38034 => "001000011101000010111001",
38035 => "000111110011010000011101",
38036 => "000110011010101000011001",
38037 => "000101010110100011010101",
38038 => "000110101110001101111011",
38039 => "001010000110000010011000",
38040 => "001100110100101111111110",
38041 => "001101111110000101001010",
38042 => "001110001101111101011110",
38043 => "001110000011011000000010",
38044 => "001100110110101011101010",
38045 => "001001001000101100110001",
38046 => "000100010000111101000100",
38047 => "000001011101100101011010",
38048 => "000000100100110101111100",
38049 => "111111100101011010110100",
38050 => "111101101100111011101111",
38051 => "111011101101000000000001",
38052 => "111010111011111001110100",
38053 => "111011101111111110001110",
38054 => "111110000110101011011101",
38055 => "000001001010000010101001",
38056 => "000100001110010011011111",
38057 => "001000001110001101000110",
38058 => "001100000010101010111100",
38059 => "001101111011110000010100",
38060 => "001110010111010001100000",
38061 => "001101011100111100111000",
38062 => "001011110110011110111011",
38063 => "001001101010110010011001",
38064 => "000101100100011000011010",
38065 => "000000101001111111111100",
38066 => "111100001101000001000100",
38067 => "111000001010110001001000",
38068 => "110101010100000111111000",
38069 => "110011110111001011000100",
38070 => "110011101000011110111010",
38071 => "110011111100010011111110",
38072 => "110100101010000000011001",
38073 => "110111000101111000110000",
38074 => "111001011111001011111111",
38075 => "111001001001110110100001",
38076 => "110111001100110111101100",
38077 => "110101101010000001001100",
38078 => "110110000110001001110010",
38079 => "111000011101110010101100",
38080 => "111010001111011000100010",
38081 => "111010011101011011110001",
38082 => "111010110001010001001111",
38083 => "111100010011100000011011",
38084 => "111110001001001011011110",
38085 => "111111001001110000000001",
38086 => "111111001001100100111001",
38087 => "111101101111100011111001",
38088 => "111011100000000000011110",
38089 => "111001001011010101010001",
38090 => "110110100000100011010000",
38091 => "110101010100101000000011",
38092 => "110111001000001000001010",
38093 => "111010001010101011100100",
38094 => "111101110000011101011100",
38095 => "000010011011001100011010",
38096 => "000111000000010000010100",
38097 => "001001111101011101000000",
38098 => "001010011111000100101010",
38099 => "001000010101010011111001",
38100 => "000100111000111111110010",
38101 => "000010111110101101111011",
38102 => "000011001110001000111010",
38103 => "000011100001110011111001",
38104 => "000011100100010001010100",
38105 => "000100111010001100101000",
38106 => "000111110011110110101010",
38107 => "001011000011011110001100",
38108 => "001101000010101111000100",
38109 => "001100101101010000011100",
38110 => "001010011101000000100000",
38111 => "000111110011110100110101",
38112 => "000101110000001011100000",
38113 => "000100001010101000110011",
38114 => "000010101100101110011110",
38115 => "000001000110010000001011",
38116 => "111111111011000001011010",
38117 => "000000000001000111000100",
38118 => "000000110101100100100011",
38119 => "000001100101110011010100",
38120 => "000001110101000100101101",
38121 => "000000100101011000011011",
38122 => "111101011110111001011000",
38123 => "111001010011110011000010",
38124 => "110101001000100001110100",
38125 => "110001100001001011011110",
38126 => "101110101110010001101100",
38127 => "101101001111101111100110",
38128 => "101101100001111101110110",
38129 => "110000010100001011101100",
38130 => "110101010110111001100010",
38131 => "111010010101111000011000",
38132 => "111101101011111001110000",
38133 => "111111000110100011100011",
38134 => "111110101110010010011110",
38135 => "111101010001101000011001",
38136 => "111010011110110000000010",
38137 => "110101111111101110101001",
38138 => "110000100101000110011000",
38139 => "101010111100011110100010",
38140 => "100110100110001110110011",
38141 => "100100111110010100011101",
38142 => "100110000001011101111101",
38143 => "101001000110101010111000",
38144 => "101101001000110011001000",
38145 => "110001100110000110001100",
38146 => "110110110010101100111110",
38147 => "111100101010110011010000",
38148 => "000010101000110111110001",
38149 => "000111100101001000101001",
38150 => "001011000111100011000101",
38151 => "001101110011111010001100",
38152 => "001111011001111011111100",
38153 => "001111100000100101010000",
38154 => "001110100110100101011100",
38155 => "001101101110110100011010",
38156 => "001101010110000111010100",
38157 => "001100110110111101111110",
38158 => "001100010001010110110110",
38159 => "001011110111111010101100",
38160 => "001100000110010100011110",
38161 => "001101101011101010000010",
38162 => "001111011010010011000000",
38163 => "001111110111100110000010",
38164 => "001111111001001111000100",
38165 => "010000110001111010111000",
38166 => "010010101111000001110010",
38167 => "010011111101110111010010",
38168 => "010011000111101100010110",
38169 => "010001011101100101001010",
38170 => "001111110010111000010000",
38171 => "001101110011011010010110",
38172 => "001011000001101100110011",
38173 => "000111110100101010010110",
38174 => "000110001000001000100111",
38175 => "000101100010100000001011",
38176 => "000100001001110000010101",
38177 => "000010001101001000010011",
38178 => "111111011111101010101100",
38179 => "111011111000101101000001",
38180 => "111000011110010001111001",
38181 => "110110000010111011101100",
38182 => "110101101001111001101100",
38183 => "110110011010110010000110",
38184 => "110110011111000110100101",
38185 => "110110110111010010001111",
38186 => "111000001011010100010110",
38187 => "111001101100001010011110",
38188 => "111011100001001111000000",
38189 => "111101111000111111111011",
38190 => "000000111000101100101101",
38191 => "000010110010000110000000",
38192 => "000001100111100011110001",
38193 => "111111011111101001000110",
38194 => "111110111011001100100011",
38195 => "111111000011100100011101",
38196 => "111110000100110010110101",
38197 => "111011101110011001100110",
38198 => "111001110011011001111100",
38199 => "111001100111101101010010",
38200 => "111010111101010101010110",
38201 => "111101001001011001111101",
38202 => "111110011000011111011001",
38203 => "111110010011101101011010",
38204 => "111110110110110000101111",
38205 => "000000000110011111110010",
38206 => "000001110110100110100110",
38207 => "000100101011011000101101",
38208 => "000110001010111011111110",
38209 => "000100010101000110000011",
38210 => "000001011000000101000111",
38211 => "111111001000111011011101",
38212 => "111100010111101110101011",
38213 => "110111111111100100100110",
38214 => "110010111011110000110000",
38215 => "101111100100000111111010",
38216 => "110000101001110010101010",
38217 => "110101100100000111111110",
38218 => "111010011001101010000100",
38219 => "111110110111010110000010",
38220 => "000100010010110111010001",
38221 => "001000001100111100100110",
38222 => "001010000001000011110001",
38223 => "001100010000001111010100",
38224 => "001110100011011000000000",
38225 => "001111001100100100000000",
38226 => "001101011110010110010000",
38227 => "001001101000111101110010",
38228 => "000101101000101110110000",
38229 => "000011101011001110110011",
38230 => "000100011101000101010000",
38231 => "000101110001010000100001",
38232 => "000101000001101111011001",
38233 => "000011000011100011111001",
38234 => "000000100001101011100111",
38235 => "111101010001100010110000",
38236 => "111010101001001110110000",
38237 => "110111110011010111100010",
38238 => "110100001000110111010000",
38239 => "110010110010010010111010",
38240 => "110101001010100011000000",
38241 => "111010001111000100000101",
38242 => "000000100101111111001000",
38243 => "000101111101111110111001",
38244 => "001010001000001011110001",
38245 => "001110011010000011110100",
38246 => "010001111011101010100100",
38247 => "010010111001101110000100",
38248 => "010001001010100110001100",
38249 => "001101110001110101001000",
38250 => "001000111111100100111011",
38251 => "000010101001010001101110",
38252 => "111011111000100100001111",
38253 => "110110011100000110010100",
38254 => "110100001010111010111100",
38255 => "110101010001000110001101",
38256 => "110110100110100000011011",
38257 => "110110001000000101101111",
38258 => "110100101101100011011110",
38259 => "110011110000000010010000",
38260 => "110100100010111111111100",
38261 => "110110000110110001001000",
38262 => "110110110000001000110001",
38263 => "111000001001110111001111",
38264 => "111011100101100100110110",
38265 => "111111110010011011101110",
38266 => "000011100110010010010011",
38267 => "000110101001110100100110",
38268 => "001001111011101010111101",
38269 => "001101110110001100001110",
38270 => "010000100100011011101000",
38271 => "010000101110000011010000",
38272 => "001110101101001011000110",
38273 => "001011110011111100010100",
38274 => "000111101111101000110111",
38275 => "000001010101000000011011",
38276 => "111010110011100111010101",
38277 => "110110101001110011010000",
38278 => "110100001100010110101011",
38279 => "110010110001110010011100",
38280 => "110001111110111110110010",
38281 => "110001101110100101100100",
38282 => "110010010011011010111110",
38283 => "110010110010100111010010",
38284 => "110011010001011001111010",
38285 => "110100001111100011000111",
38286 => "110100111100100010110100",
38287 => "110101100011111010010010",
38288 => "110110101011101010111000",
38289 => "111000110011111001101110",
38290 => "111011111001000110110111",
38291 => "111110011000000011000110",
38292 => "000000000011010101101100",
38293 => "000001100000101101101110",
38294 => "000010010100001011010001",
38295 => "000010100010101100011110",
38296 => "000001100001010000111000",
38297 => "111110001111101110110100",
38298 => "111001011001000010001110",
38299 => "110011100111111001111110",
38300 => "101101101110010101010000",
38301 => "101001001010001100001110",
38302 => "100110100110101000110010",
38303 => "100101111111110110000101",
38304 => "100111010010110010000111",
38305 => "101010110010000010110010",
38306 => "110000100000111100000110",
38307 => "110111011011000011101100",
38308 => "111110001010100101010100",
38309 => "000100010101011100001111",
38310 => "001010000110101001010111",
38311 => "001110101111101010001010",
38312 => "010000110011001100100000",
38313 => "010000001100000001101110",
38314 => "001110011011000110100000",
38315 => "001100110011100001001010",
38316 => "001011011101001010110011",
38317 => "001010000110100010110001",
38318 => "001000110001000011111100",
38319 => "000111100011011100010101",
38320 => "000110100100010001000111",
38321 => "000101101100101100000100",
38322 => "000101011000011000010000",
38323 => "000110101010111111001010",
38324 => "001001001111011100101001",
38325 => "001100000101101010110010",
38326 => "001110100001010011100110",
38327 => "001111011010010111100110",
38328 => "001110111010100001101110",
38329 => "001110000110000101001010",
38330 => "001101000011001010000110",
38331 => "001011100111011111101111",
38332 => "001001011111011111111011",
38333 => "000111000000100110110000",
38334 => "000101000011011001100001",
38335 => "000011100001110101100010",
38336 => "000010000110101000101001",
38337 => "111111101101000101011101",
38338 => "111011110110110000110111",
38339 => "111001001001001010000010",
38340 => "111000110100010100100010",
38341 => "111001010001111101000000",
38342 => "111010001110101101100010",
38343 => "111011110101001001010010",
38344 => "111100111001110000010110",
38345 => "111100101111100001101100",
38346 => "111100000001100010100000",
38347 => "111011100100111101011110",
38348 => "111011101101011001001110",
38349 => "111100000101000001101010",
38350 => "111011101000010011001001",
38351 => "111010110001101111001111",
38352 => "111011001111101100110011",
38353 => "111100100100101101001100",
38354 => "111101111001000000000100",
38355 => "111111111110101011001011",
38356 => "000010100000111010000011",
38357 => "000100010011011000011111",
38358 => "000101010010011111110100",
38359 => "000101100011001111110010",
38360 => "000100100001010011000000",
38361 => "000010010100001110001011",
38362 => "111111111111001000000100",
38363 => "111101111001110101100001",
38364 => "111100010000001001111001",
38365 => "111011111000011100110111",
38366 => "111101000100010011100110",
38367 => "111111001011111000000000",
38368 => "000001110001000111000111",
38369 => "000101000010111100001100",
38370 => "000111101100011000011111",
38371 => "000110110001101101010000",
38372 => "000010110100010101110011",
38373 => "111110101000100111010111",
38374 => "111010111010010101101110",
38375 => "110111011111011011010101",
38376 => "110100011011101000111110",
38377 => "110010011101101010001110",
38378 => "110010010001111101000110",
38379 => "110011010111110011001010",
38380 => "110110000101100101110010",
38381 => "111010010011111010011011",
38382 => "111111001101011111100011",
38383 => "000100110100110101000011",
38384 => "001000101010010001110101",
38385 => "001001000100001110101001",
38386 => "001000100001001011110100",
38387 => "000111110101111001101011",
38388 => "000111000011111000101110",
38389 => "000110110000110000010111",
38390 => "000101100000111000111011",
38391 => "000011010111000110110100",
38392 => "000010011010000101000101",
38393 => "000011000100110111110100",
38394 => "000011110100110101111011",
38395 => "000011011000111100100110",
38396 => "000010010010000011111001",
38397 => "000000110101101010010000",
38398 => "111111110001011011001001",
38399 => "000000110100100000110010",
38400 => "000010011101111111110010",
38401 => "000010111011010100010011",
38402 => "000011110111010011011111",
38403 => "000101010111010010111110",
38404 => "000110100110010101011110",
38405 => "001000100001111100111110",
38406 => "001010100000011011110110",
38407 => "001011110010010110110010",
38408 => "001101101000001110100010",
38409 => "001111001010110111000110",
38410 => "001110011100110010010100",
38411 => "001100101010011101001000",
38412 => "001011000101110101000111",
38413 => "001001000101111000101010",
38414 => "000111010111110000011100",
38415 => "000110011011111010111001",
38416 => "000100011010000101010001",
38417 => "000001010000001001111110",
38418 => "111111100101111100101011",
38419 => "111111011110110100111101",
38420 => "111110110100100000110011",
38421 => "111101111100011001001010",
38422 => "111101110011111011001110",
38423 => "111101101000111011000000",
38424 => "111101010101110000100111",
38425 => "111101011010011001000010",
38426 => "111101111101110010000100",
38427 => "111111010100100111100100",
38428 => "000001000001011110100110",
38429 => "000010011110000001000110",
38430 => "000100001010110010101001",
38431 => "000111000000001010010100",
38432 => "001010110011110011111110",
38433 => "001101000011001101000110",
38434 => "001011010101010000100000",
38435 => "000101111011100101110001",
38436 => "111110011100011111010011",
38437 => "110111001000000111110010",
38438 => "110001001001001011111100",
38439 => "101100000011110101100000",
38440 => "101000001011111001101000",
38441 => "100101111001010011111010",
38442 => "100101011001101100101111",
38443 => "100111000110000101111000",
38444 => "101010100111001001110010",
38445 => "101111011100010001101110",
38446 => "110100011101110100001011",
38447 => "111001001110011111011110",
38448 => "111110011001100010001101",
38449 => "000010011101101011010101",
38450 => "000100000100000001001010",
38451 => "000011100100010011011101",
38452 => "000000111010101101001111",
38453 => "111101100111001111100100",
38454 => "111011001100011101111010",
38455 => "111001100010000011101010",
38456 => "111000101001011110010100",
38457 => "110111001111101010011000",
38458 => "110100100011111100101111",
38459 => "110001111001101010011100",
38460 => "101111101101010111001010",
38461 => "101110011001010100010110",
38462 => "101110000101110101000000",
38463 => "101101111001001001110110",
38464 => "101101110111011101011100",
38465 => "101110110111101100110010",
38466 => "110010010000100101011010",
38467 => "111000000010110111111001",
38468 => "111110001100011011001000",
38469 => "000100001011010111101000",
38470 => "001010001100100000101000",
38471 => "001111101010001010000110",
38472 => "010100001001010000010000",
38473 => "010110110001001100111100",
38474 => "010111001111101110011110",
38475 => "010101101100110110111000",
38476 => "010010001001101100111100",
38477 => "001110010000001101011010",
38478 => "001010111001011010100011",
38479 => "000111010111101001001001",
38480 => "000100001000101000000110",
38481 => "000001101101000101101111",
38482 => "000000010100011001101110",
38483 => "000001000101010001000000",
38484 => "000011111010100010011000",
38485 => "000110111000111000101110",
38486 => "001001001011110100001011",
38487 => "001011111001000011101110",
38488 => "001110100100010000011100",
38489 => "001111010010000000111110",
38490 => "001110001101001110000000",
38491 => "001100001011001010100000",
38492 => "001000111000010010100000",
38493 => "000100100100101100000100",
38494 => "111111101000101000000100",
38495 => "111010010011000010001000",
38496 => "110101010101010011010000",
38497 => "110000011101101010010000",
38498 => "101011011110110100011010",
38499 => "101001000101011100001100",
38500 => "101011010110100101110010",
38501 => "110000010000100010010000",
38502 => "110101011110100110111110",
38503 => "111010011100011101010011",
38504 => "111110011111110100110000",
38505 => "000001011001001011011010",
38506 => "000011001000001011011010",
38507 => "000011001101010001110011",
38508 => "000001100111011111100110",
38509 => "111110010011100101001110",
38510 => "111001101110111011101001",
38511 => "110110000001010010010111",
38512 => "110100011010010011111010",
38513 => "110100000111010011110010",
38514 => "110100110110010010000000",
38515 => "110111011110101100111000",
38516 => "111100000000001110111011",
38517 => "000001001100011100011000",
38518 => "000101111101000011010110",
38519 => "001001000110111100001110",
38520 => "001001111010111010101100",
38521 => "001001011111110111000010",
38522 => "001000011111010010011011",
38523 => "000110000111011011000011",
38524 => "000011110000001011110100",
38525 => "000011101101111110010010",
38526 => "000100111000001010111100",
38527 => "000101001001100100010110",
38528 => "000101000011111001010111",
38529 => "000101101000111000101010",
38530 => "000110110010100000011001",
38531 => "000111111000000001100000",
38532 => "001000101110011100010000",
38533 => "001010001011001000000100",
38534 => "001011011100110100001110",
38535 => "001010010111010111000011",
38536 => "000111001000000101111010",
38537 => "000011000111100010011100",
38538 => "111110110000101110100001",
38539 => "111001111001101011110010",
38540 => "110100011101110110110110",
38541 => "110000000010000010110000",
38542 => "101101110010110011111010",
38543 => "101101011010010100111110",
38544 => "101111010010000000110100",
38545 => "110010111111110110111010",
38546 => "111000000010110111110001",
38547 => "111110001111110101011001",
38548 => "000010111111110000110111",
38549 => "000101100100101110001100",
38550 => "000111000111001100110001",
38551 => "000110011011101010100000",
38552 => "000100010011111100001010",
38553 => "000001110010010000111011",
38554 => "111101010001011100001101",
38555 => "111000000001100111011011",
38556 => "110100111110011001100001",
38557 => "110101001010011011010100",
38558 => "110111101100111111001100",
38559 => "111010010011000000001100",
38560 => "111100001010010001101001",
38561 => "111101011101000111100101",
38562 => "111110000011110001000011",
38563 => "111101111001011011100111",
38564 => "111011110110111001110110",
38565 => "111001000100101110000100",
38566 => "110111111101110110111110",
38567 => "110111110101011101111001",
38568 => "111000100101100001010111",
38569 => "111010011011000111111000",
38570 => "111100001011010000001111",
38571 => "111111011110010100110100",
38572 => "000101010000001011001111",
38573 => "001010100010111100001011",
38574 => "001101100110100101010100",
38575 => "001110110011010110101110",
38576 => "001110100000101100101010",
38577 => "001101010110001110010010",
38578 => "001011101001000001001110",
38579 => "001000110010001001110000",
38580 => "000101100111101011100101",
38581 => "000100111100101101110011",
38582 => "000110100100111011110100",
38583 => "000111011111011101011011",
38584 => "000111001101111010001010",
38585 => "000110111100001000000010",
38586 => "000111000000010110001000",
38587 => "000111000111101100011111",
38588 => "000110010101100101110100",
38589 => "000101010000101000101001",
38590 => "000110011001101101100101",
38591 => "001001101100010111110100",
38592 => "001100010111110101100010",
38593 => "001110000110101011101000",
38594 => "010000011111110010110000",
38595 => "010010111110000010010100",
38596 => "010100001010011111110100",
38597 => "010011011011011101100000",
38598 => "001111110001000001100100",
38599 => "001010000000101001011000",
38600 => "000100110000110110101101",
38601 => "000000111100111001111100",
38602 => "111110001001011001100011",
38603 => "111011111000110001110011",
38604 => "111001111110011010010100",
38605 => "111001000111100011011010",
38606 => "111001100111101011011000",
38607 => "111010100010011010010110",
38608 => "111011110000110011011000",
38609 => "111101101011101100010100",
38610 => "111110001110111110100000",
38611 => "111011010000100010100000",
38612 => "110110010011010010010110",
38613 => "110001100100001000110110",
38614 => "101101100100010100000100",
38615 => "101011001001001011000110",
38616 => "101010111111001111101110",
38617 => "101100100010111101101100",
38618 => "101110111010110000111010",
38619 => "110001110010101000100000",
38620 => "110101110000110000010100",
38621 => "111011000110110001000100",
38622 => "000000011001000111100000",
38623 => "000011110000010010101111",
38624 => "000101001000111110110010",
38625 => "000101100001011001010000",
38626 => "000100111101100101110011",
38627 => "000011010111110010001100",
38628 => "000000101011111011111001",
38629 => "111101000010101001011110",
38630 => "111010011111010000010101",
38631 => "111010011110110001101101",
38632 => "111011101011111001111000",
38633 => "111101101010011111101000",
38634 => "000001011101110011011110",
38635 => "000101111111011000000001",
38636 => "001001000011100111010001",
38637 => "001011000100011011010010",
38638 => "001101001100101111100010",
38639 => "001110110010100111111100",
38640 => "001111001110000010010100",
38641 => "001110000100100011011110",
38642 => "001100000110010001101010",
38643 => "001100011011011000111100",
38644 => "001110111000101101100000",
38645 => "001111111100110110111100",
38646 => "001111000011010001110100",
38647 => "001100101011100100110000",
38648 => "001000110110100000010110",
38649 => "000101011010010111111101",
38650 => "000011110011111111111010",
38651 => "000010110011011100110010",
38652 => "000000010110001000101010",
38653 => "111100011001101010111011",
38654 => "110111100111111101100110",
38655 => "110010011010001100010000",
38656 => "101110111000100011100110",
38657 => "101101010110001100111000",
38658 => "101100000110000100010100",
38659 => "101100110100001001111110",
38660 => "110000101011101000011010",
38661 => "110101110011111010010010",
38662 => "111010110110001101111101",
38663 => "111110100110100001111111",
38664 => "000001001110110001100011",
38665 => "000011111110000010000110",
38666 => "000110000000001110110110",
38667 => "000101111111110011101110",
38668 => "000011001011100001100001",
38669 => "111101100110001010111001",
38670 => "110110110101110111011000",
38671 => "110000111011100101001000",
38672 => "101101011001101011011100",
38673 => "101011110111000100000010",
38674 => "101011101010100110000010",
38675 => "101110000100011000000100",
38676 => "110010001111010010011100",
38677 => "110110001000101110101010",
38678 => "111010111011001010000010",
38679 => "000001101001111110011111",
38680 => "001000000101000011101010",
38681 => "001011010000011010000010",
38682 => "001011011011101101101110",
38683 => "001011010001010010100001",
38684 => "001011001001111110111111",
38685 => "001001111000001000001010",
38686 => "000111110010011101110011",
38687 => "000101110010100000111111",
38688 => "000100010100110101111011",
38689 => "000011110000101011101011",
38690 => "000100100110001010111001",
38691 => "000110101110011011000000",
38692 => "001000110010101101000100",
38693 => "001010011001001110100110",
38694 => "001100101010010111000110",
38695 => "001111101110011011001010",
38696 => "010010011000010000000100",
38697 => "010011010011011110111110",
38698 => "010001100001111111001100",
38699 => "001100101110100111100010",
38700 => "000101100010100000011010",
38701 => "111101101101100001101010",
38702 => "110110110100101010000110",
38703 => "110000100101001011110010",
38704 => "101010011000001101101100",
38705 => "100101111100011010101110",
38706 => "100101100001000000001001",
38707 => "101001000001011010000000",
38708 => "101111001100110011101110",
38709 => "110110111011011000000111",
38710 => "111110101110110110110001",
38711 => "000100110010001100000000",
38712 => "001000000111111101101111",
38713 => "001000111100101101011101",
38714 => "000110111001000101011000",
38715 => "000010010001100001000010",
38716 => "111101100101001000101111",
38717 => "111001101111110111100110",
38718 => "110101111101111010011000",
38719 => "110010110000000110011110",
38720 => "110000110010000001011100",
38721 => "110000001110100001110100",
38722 => "110000100110111000111010",
38723 => "110000101100001010000110",
38724 => "110000010110110000001010",
38725 => "101111110011100000001100",
38726 => "101110111101100011001000",
38727 => "101110010010101011100110",
38728 => "101101100010000100001010",
38729 => "101100011011011101111110",
38730 => "101011101000010110011010",
38731 => "101011111101011000010000",
38732 => "101110101100000010110010",
38733 => "110011101111101001010110",
38734 => "111001010011010000110011",
38735 => "111110110001111110011110",
38736 => "000100011111110100011001",
38737 => "001001100101110111100100",
38738 => "001100100000011011100110",
38739 => "001100100011000111010100",
38740 => "001010101100110000011010",
38741 => "001000100001101101101110",
38742 => "000110010111000100110110",
38743 => "000011010100000101111000",
38744 => "111111100000001000011110",
38745 => "111100101011000101110000",
38746 => "111011111001011101011110",
38747 => "111100100111011000100101",
38748 => "111101111001111110111001",
38749 => "111111110111011000010011",
38750 => "000011010100011111101111",
38751 => "000111110110100100111010",
38752 => "001011110100110110000101",
38753 => "001110010000101101110100",
38754 => "001111101110001011111100",
38755 => "010001010100000111000000",
38756 => "010010111110010100000110",
38757 => "010100010110110011000100",
38758 => "010101011100100101100010",
38759 => "010101101011011100111010",
38760 => "010101010100000000000010",
38761 => "010100100111010111010110",
38762 => "010010011100111010011000",
38763 => "001110110001010101100110",
38764 => "001010110000010110111000",
38765 => "000111010100010111101001",
38766 => "000100111000110011011011",
38767 => "000011000110001100000010",
38768 => "000001101001011110110111",
38769 => "000000011010111010111101",
38770 => "111111011001111110000111",
38771 => "111110111111011111110111",
38772 => "111110110000100001100110",
38773 => "111110010000101000010000",
38774 => "111101101011000011101101",
38775 => "111100110100110101001111",
38776 => "111011101110111010000100",
38777 => "111010100011100111110100",
38778 => "111010001011011110001101",
38779 => "111011101100011010011111",
38780 => "111110001001011001010101",
38781 => "000000010100110100011001",
38782 => "000001101110111000001110",
38783 => "000010001110010111010010",
38784 => "000011000100001000100000",
38785 => "000100000001100111100011",
38786 => "000011010110010010010111",
38787 => "000001011000111010100000",
38788 => "111110101111010010010100",
38789 => "111010011011101011111100",
38790 => "110011110101100111001110",
38791 => "101101000001001011011110",
38792 => "101001100111011100101010",
38793 => "101001111101000001100100",
38794 => "101100011001001101001000",
38795 => "110000101111110001111110",
38796 => "110110001011001110000101",
38797 => "111011100100110001011011",
38798 => "000000101011010010000101",
38799 => "000101101011100100100100",
38800 => "001011011011111011100010",
38801 => "010000101000101110000000",
38802 => "010011000110111011010000",
38803 => "010100001001101011001000",
38804 => "010101000111001111100000",
38805 => "010100010101110100000000",
38806 => "010000010111011110111110",
38807 => "001010011100101001111000",
38808 => "000101010011001101011101",
38809 => "000001001111010000011111",
38810 => "111100100011110110100100",
38811 => "110111111110110111101110",
38812 => "110101000000100111110011",
38813 => "110010011010100101111100",
38814 => "101111010011111010100110",
38815 => "101101101010010010010000",
38816 => "101111001000010101011100",
38817 => "110010101010101010001100",
38818 => "110110001101101111000101",
38819 => "111001011111010010100010",
38820 => "111101111111110001000000",
38821 => "000100001000111011010100",
38822 => "001001110101101111000001",
38823 => "001101001000011111000000",
38824 => "001111000111100100110100",
38825 => "010001100010000100000000",
38826 => "010010010101000011111110",
38827 => "001111010100010001010110",
38828 => "001011001000101000001100",
38829 => "001000100100110011100000",
38830 => "000110000101101111011001",
38831 => "000001001010111110000110",
38832 => "111011000010000001000111",
38833 => "110111110100111001001001",
38834 => "111000001101010011010000",
38835 => "111000010100011010100000",
38836 => "110110100100111001101001",
38837 => "110101100101010110000100",
38838 => "110111111101100011111100",
38839 => "111100101000000100110011",
38840 => "000000011011000011001101",
38841 => "000011111011111100101100",
38842 => "001001101110110111001101",
38843 => "010000010111001010011110",
38844 => "010100101101000010100100",
38845 => "010110001111011011001110",
38846 => "010101111100111101001110",
38847 => "010011110110000111100100",
38848 => "001111011100011001100000",
38849 => "001001111110100100001101",
38850 => "000101011001101111001011",
38851 => "000010001011010010001000",
38852 => "111111110101000011001100",
38853 => "111110011101000001110001",
38854 => "111111000100101101010001",
38855 => "000001101111010110010010",
38856 => "000100100110111010110010",
38857 => "000111000110111010010111",
38858 => "001010011000011010000111",
38859 => "001101100110000001010000",
38860 => "001110101101010101010110",
38861 => "001101110010000111111100",
38862 => "001011101010000011100000",
38863 => "001000010101000111011100",
38864 => "000100000010101000011101",
38865 => "111111001100100101001001",
38866 => "111010011011100001001110",
38867 => "110110011011101010011000",
38868 => "110010101011011000110000",
38869 => "101111000010110110110110",
38870 => "101100110010010001110010",
38871 => "101100010111110010101100",
38872 => "101100110010001110011110",
38873 => "101100111011010100010110",
38874 => "101110000100011000100110",
38875 => "110010010001101111001000",
38876 => "110111111010111100010110",
38877 => "111100000110001110000010",
38878 => "111110011010101100010001",
38879 => "111111100101110001010101",
38880 => "111111101100010101100010",
38881 => "111110000000001100110010",
38882 => "111011001000101110100011",
38883 => "111000101100100001110001",
38884 => "110110101001110101001100",
38885 => "110101010001000001011100",
38886 => "110100111000000110110010",
38887 => "110100111100001010010100",
38888 => "110101101110100101100000",
38889 => "110101110001110010100010",
38890 => "110100000001100000001111",
38891 => "110011001100110011011010",
38892 => "110011011100011011010010",
38893 => "110010010110011100101000",
38894 => "110000001000111101011110",
38895 => "101101101100000111001110",
38896 => "101100010101000010101110",
38897 => "101101110001101000011010",
38898 => "110001101000011101101100",
38899 => "110110111101000101110000",
38900 => "111101101010110100110111",
38901 => "000100111010101111100111",
38902 => "001010000101110000101001",
38903 => "001011100101101110111000",
38904 => "001011000010011011000001",
38905 => "001001101001010001110011",
38906 => "000110101000000010000001",
38907 => "000001100010111110100100",
38908 => "111011001011101001001000",
38909 => "110110010000100011001010",
38910 => "110100110101000001000000",
38911 => "110101011111010110011101",
38912 => "110111001001011011001110",
38913 => "111010001011011101010100",
38914 => "111101110100001000100111",
38915 => "000001001011101100110010",
38916 => "000011111000110011110010",
38917 => "000100110001011111101111",
38918 => "000011100110111111100011",
38919 => "000010100001100101100101",
38920 => "000011000000000000000100",
38921 => "000100010001000101011111",
38922 => "000101111111110111011010",
38923 => "001000010100111000110001",
38924 => "001010100101001100000000",
38925 => "001100011101001101001000",
38926 => "001101100001110001010000",
38927 => "001101010100101111111000",
38928 => "001100011000101010001000",
38929 => "001010101010010011001100",
38930 => "001000000100000101101010",
38931 => "000101110000111011000101",
38932 => "000100000010110001010100",
38933 => "000010100000011110100110",
38934 => "000001110011100101010100",
38935 => "000010010100011000000101",
38936 => "000011001110111000000011",
38937 => "000011101110111001110100",
38938 => "000100000110100110110011",
38939 => "000100100000001101000011",
38940 => "000011101111010110100000",
38941 => "000001100000101100000111",
38942 => "111111001000001010010111",
38943 => "111101100111111111000000",
38944 => "111101011111000101011000",
38945 => "111101111110011101001100",
38946 => "111110010010000111011100",
38947 => "111111101110100100110001",
38948 => "000010101011011000010111",
38949 => "000101100101000010100111",
38950 => "001000000110101111010010",
38951 => "001010010111100001011010",
38952 => "001011111101001111000010",
38953 => "001100000111101011001100",
38954 => "001001111010101011100000",
38955 => "000110001110101111100011",
38956 => "000010100001111101001010",
38957 => "111111001000000101110110",
38958 => "111100011000010110000011",
38959 => "111010100100101001111000",
38960 => "111010101010110101111011",
38961 => "111101001001110010010100",
38962 => "111111100011100011000111",
38963 => "000000010101011010000100",
38964 => "000000100000011011101110",
38965 => "000000110101000111011100",
38966 => "000001001111111010011100",
38967 => "000000000001000010001000",
38968 => "111100000000101010011010",
38969 => "110111010010000000000101",
38970 => "110011011000101010100010",
38971 => "110000100101000001111010",
38972 => "101111000111101000101100",
38973 => "101101111100000011000110",
38974 => "101100001101011110010100",
38975 => "101011011001100010011100",
38976 => "101101101000010010010100",
38977 => "110010110000111101010110",
38978 => "111000101000110011110001",
38979 => "111110010010110011110010",
38980 => "000011101100100110000111",
38981 => "001000010100000110111010",
38982 => "001011110101010001010010",
38983 => "001101100100101101001100",
38984 => "001101010100010000001100",
38985 => "001011100100110100101000",
38986 => "000111110000001110010111",
38987 => "000010011011110011000010",
38988 => "111110011001000101001111",
38989 => "111100100100110110010110",
38990 => "111011101111110010100001",
38991 => "111011011000000100110111",
38992 => "111011111101001001110011",
38993 => "111110000011111000000101",
38994 => "000001100010111101111010",
38995 => "000100011111000001010010",
38996 => "000101000111100101010011",
38997 => "000100110010111100110110",
38998 => "000101001011000000100111",
38999 => "000101111011001111011011",
39000 => "000111001000100001101100",
39001 => "001001000100010110101100",
39002 => "001011100001110110101100",
39003 => "001110001011001101010010",
39004 => "001111101101010100011000",
39005 => "001111111111110000110010",
39006 => "010000100010011110101110",
39007 => "010000110110010001010100",
39008 => "001110101100000010111100",
39009 => "001001101000100010011111",
39010 => "000100100100111000111100",
39011 => "000010000010111101101011",
39012 => "000000011111100010111011",
39013 => "111110010101101111100001",
39014 => "111100101101001101111001",
39015 => "111100010011110010011110",
39016 => "111101001101001000101110",
39017 => "111111010110101100010101",
39018 => "000010001101101111010011",
39019 => "000101100010001100011010",
39020 => "001000011011101101111000",
39021 => "001001011011111001101011",
39022 => "001000111110100010011101",
39023 => "001000110111100101011001",
39024 => "001000111101011110011010",
39025 => "000111011101111010110101",
39026 => "000100110010011010001000",
39027 => "000010001011010010011000",
39028 => "111110001110010011001001",
39029 => "110111111000100001010100",
39030 => "110000010001101110011110",
39031 => "101000100000111001010100",
39032 => "100010111000010000011110",
39033 => "100001011111110011111101",
39034 => "100010010010110111001011",
39035 => "100010111000000111111101",
39036 => "100101011101001000100110",
39037 => "101100010100000011100010",
39038 => "110101011100110100001110",
39039 => "111110010101001001110101",
39040 => "000101110111111101101010",
39041 => "001010010111000111001011",
39042 => "001011100000110111100100",
39043 => "001011000000010000010111",
39044 => "001000100111011111010100",
39045 => "000011111110101101011111",
39046 => "111111000011010100100101",
39047 => "111011010010110101110001",
39048 => "111001000000000100110000",
39049 => "111000100110000111101110",
39050 => "111010010000110010110010",
39051 => "111101100000010110100011",
39052 => "000000111101100110100011",
39053 => "000011000101000010100101",
39054 => "000010110110110101111010",
39055 => "000000101100110111100001",
39056 => "111110100111011100111110",
39057 => "111101000111110001010100",
39058 => "111011000100010101110011",
39059 => "111000110001010101010100",
39060 => "110111000010010111111100",
39061 => "110111000001011010011100",
39062 => "111010000111010110100100",
39063 => "111110101111000101001110",
39064 => "000011011000101000010100",
39065 => "001001010100110000101010",
39066 => "001111100000101001000100",
39067 => "010011000010110101000110",
39068 => "010011111100001110010110",
39069 => "010011000111001110011110",
39070 => "001111110001111100010100",
39071 => "001010010001101010100001",
39072 => "000100100101001010111011",
39073 => "111110110010100100101001",
39074 => "111000110000110111110000",
39075 => "110100011101100111101000",
39076 => "110010011011011100000100",
39077 => "110010010000010101011110",
39078 => "110100001010011101010010",
39079 => "110110101011110110100000",
39080 => "111001000110100111111000",
39081 => "111011110111111000010000",
39082 => "111101011010000111011101",
39083 => "111101100100101011011011",
39084 => "111110101011010110011110",
39085 => "000000110101111000010011",
39086 => "000010011000001100000011",
39087 => "000011000111000111001101",
39088 => "000100001110111110110110",
39089 => "000101101011101011010110",
39090 => "000111000001001101110101",
39091 => "001000101101001101111000",
39092 => "001001001010010001100100",
39093 => "000111000110101100001001",
39094 => "000100011000011000101101",
39095 => "000001010101010011000011",
39096 => "111101101100011110010111",
39097 => "111010111100001111011110",
39098 => "111000011110001010101101",
39099 => "110100111101000010010010",
39100 => "110001011101100000001010",
39101 => "101111111111011110001010",
39102 => "110001101010011110001010",
39103 => "110101000001001110110100",
39104 => "110111101101110111010011",
39105 => "111001110110111011001001",
39106 => "111100111011100000101010",
39107 => "000001011001101110010011",
39108 => "000110000000000111010001",
39109 => "001001111100001101101000",
39110 => "001110001011011100110000",
39111 => "010010000111011001000010",
39112 => "010100011000101110010000",
39113 => "010101110000101110010100",
39114 => "010110100000101001101100",
39115 => "010101101010001001011000",
39116 => "010010101101011010100000",
39117 => "001101111000000101100110",
39118 => "001000101110000110001000",
39119 => "000100000111110110011001",
39120 => "111111000101001000010010",
39121 => "111001111010011011010000",
39122 => "110110000111000000110101",
39123 => "110100011000110010111100",
39124 => "110101011010101110010111",
39125 => "111001000001101111000001",
39126 => "111101110101010100000001",
39127 => "000010101101101001010101",
39128 => "000110001100010111000011",
39129 => "000111000101101011010000",
39130 => "000110111111010000100101",
39131 => "000111100101000110001010",
39132 => "000110111010011001001000",
39133 => "000010110010011010011000",
39134 => "111100100101011001100011",
39135 => "110111010001001000000000",
39136 => "110100101010110011010001",
39137 => "110100100001010001010110",
39138 => "110101011110001100000010",
39139 => "110111100100001001110011",
39140 => "111011000010111011111000",
39141 => "111110000011110111100000",
39142 => "111111011011011000100011",
39143 => "000000011110010001010101",
39144 => "000001100001010101001111",
39145 => "000000100100101111110011",
39146 => "111100100101000101110100",
39147 => "110111000100011000010100",
39148 => "110010100111101010011000",
39149 => "110000101100110100011010",
39150 => "110000101111111000111000",
39151 => "110010000000101111101110",
39152 => "110101000001011101111010",
39153 => "111001111110110110111101",
39154 => "111111110110111010010010",
39155 => "000101011100011100100010",
39156 => "001010010001010110011000",
39157 => "001110001110001111110110",
39158 => "010000010011100111000000",
39159 => "010000011011001010111110",
39160 => "010000100010110000001000",
39161 => "010000110111010101100100",
39162 => "001111101110111110011100",
39163 => "001100111100110111010110",
39164 => "001001000110001001010000",
39165 => "000101001001000000100101",
39166 => "000001111101100110110001",
39167 => "111110111101100111010100",
39168 => "111011111110011000011111",
39169 => "111001100011111010010011",
39170 => "110111111011111100101011",
39171 => "111000000010000000000110",
39172 => "111010001101001011000101",
39173 => "111101001111001010010010",
39174 => "111111110101000111011001",
39175 => "000001011110110101101011",
39176 => "000011001101010100010111",
39177 => "000101111010111101011010",
39178 => "001000100111100000011101",
39179 => "001010011110111011011110",
39180 => "001011011101110101000111",
39181 => "001011000101000111110001",
39182 => "001001010000101000000111",
39183 => "000111010011100110001101",
39184 => "000110111001100101111010",
39185 => "000111010010111000001010",
39186 => "000101111110111100000100",
39187 => "000010101011100101010101",
39188 => "111110100010111101100110",
39189 => "111010000010001010001101",
39190 => "110101101101000011101000",
39191 => "110001111011100000000100",
39192 => "101110110100111110100110",
39193 => "101100111011000110100110",
39194 => "101100010110100001001100",
39195 => "101100101010010010000010",
39196 => "101110000011110110101010",
39197 => "110001010111011110001110",
39198 => "110101011011100010101111",
39199 => "110111101010110101101111",
39200 => "111000010100100011101101",
39201 => "111001100011100010101100",
39202 => "111011111001000010100110",
39203 => "111110000010100101010100",
39204 => "111110010110110101001000",
39205 => "111101010111111100010101",
39206 => "111100110110000111111000",
39207 => "111100011101000010111010",
39208 => "111011101001100100000010",
39209 => "111010110001000001000001",
39210 => "111010000111110111111100",
39211 => "111010110110011000111010",
39212 => "111100110111001010011000",
39213 => "111110100110001011100100",
39214 => "111111111011111011000010",
39215 => "000001011011010010001001",
39216 => "000011001111111000011111",
39217 => "000101000100001011000000",
39218 => "000101111011111001111000",
39219 => "000101100100110010011100",
39220 => "000011111001000001111011",
39221 => "000001011100100100001011",
39222 => "111111011011110101111111",
39223 => "111101001010001001011100",
39224 => "111010001111000111101111",
39225 => "111000001011100110000010",
39226 => "111000001001100010110001",
39227 => "111011001100110001011101",
39228 => "000000010011011101011110",
39229 => "000100110010010100110100",
39230 => "001001011100001001001010",
39231 => "001111001101000110010100",
39232 => "010011010111001010111100",
39233 => "010011011111101111010110",
39234 => "001111010110000111111000",
39235 => "001000101101101111100011",
39236 => "000010001000111101101010",
39237 => "111011111000110101010110",
39238 => "110101010111000010011001",
39239 => "101111101100101010001000",
39240 => "101100111010110101000010",
39241 => "101101100111000011110100",
39242 => "110000011011110110000100",
39243 => "110100010111011111110110",
39244 => "111000111111010001000001",
39245 => "111101100011111111111101",
39246 => "000001001110010011000000",
39247 => "000010001100101001110110",
39248 => "000000001010000011101010",
39249 => "111110001011110010110111",
39250 => "111110000100101110111101",
39251 => "111110100111110110000101",
39252 => "111110110000100100011000",
39253 => "111110100110011010111100",
39254 => "111111010110111110000101",
39255 => "000001011011111000111011",
39256 => "000011000001000100011001",
39257 => "000010110100010000001011",
39258 => "000001101010010001110011",
39259 => "000000010011110101111010",
39260 => "111101110010011101011100",
39261 => "111001101001000110110011",
39262 => "110101111101011001101011",
39263 => "110100000101011000010000",
39264 => "110011011001001000101100",
39265 => "110100001101100110010101",
39266 => "110111000011101000110100",
39267 => "111011001010011001101101",
39268 => "111111011110111000011110",
39269 => "000011011010010100111101",
39270 => "000111011010011111101010",
39271 => "001011100000101101011110",
39272 => "001110001100101111010000",
39273 => "001111010001001011101110",
39274 => "001111110100010011010100",
39275 => "001111101110011100111110",
39276 => "001110101110100101100100",
39277 => "001101100001110110111000",
39278 => "001100101001101101111010",
39279 => "001011111110000100010010",
39280 => "001011000111110110101001",
39281 => "001001111101000111001010",
39282 => "001000101011000111011011",
39283 => "000111011000001000100101",
39284 => "000101101000010000000111",
39285 => "000011001001001101010011",
39286 => "000000100100111110110100",
39287 => "111110101000010010110011",
39288 => "111101011001001101000110",
39289 => "111101010111010010111111",
39290 => "111111000010111111000111",
39291 => "000001101111100000001101",
39292 => "000100010010001000110001",
39293 => "000101011000110110011100",
39294 => "000011111000100001111101",
39295 => "000001000001110001110011",
39296 => "111111011111101010101010",
39297 => "111111011100010101001110",
39298 => "111111101101010010010011",
39299 => "000000000111110000011101",
39300 => "000000101110100000111001",
39301 => "000001111110001100011001",
39302 => "000011110101011110111111",
39303 => "000101010110000110100000",
39304 => "000111000010000010111111",
39305 => "001001010000100111111101",
39306 => "001010000010011100000110",
39307 => "001000100101000100011101",
39308 => "000110011010100001010000",
39309 => "000100101111011000100101",
39310 => "000011100111101101010001",
39311 => "000010101101110100100001",
39312 => "000010011111011111000110",
39313 => "000011101110100000011110",
39314 => "000101110001001000100110",
39315 => "000111100001000001011011",
39316 => "001001011010010010011000",
39317 => "001011111101101100010010",
39318 => "001101001110111101100100",
39319 => "001011111100001100100111",
39320 => "001010101011010001101110",
39321 => "001011000110001111010110",
39322 => "001011101010010011101010",
39323 => "001010100001101010100011",
39324 => "000101011001000001110111",
39325 => "111100010101000111100010",
39326 => "110011101010011110111010",
39327 => "101110001001110001111000",
39328 => "101011111001101001001110",
39329 => "101100010100011010111110",
39330 => "101101011111111111000000",
39331 => "101111010011011011011010",
39332 => "110011001010101010000110",
39333 => "111000011001101101000111",
39334 => "111110010100011010110100",
39335 => "000100111001111001000101",
39336 => "001010100101001000101011",
39337 => "001101111010000011000100",
39338 => "001111010010110000110010",
39339 => "001111101010001001100010",
39340 => "001110100111010100001100",
39341 => "001010110010111011011101",
39342 => "000011111110001010101000",
39343 => "111100001010000000010100",
39344 => "110110101111100111111000",
39345 => "110100110110101111110100",
39346 => "110011111110001111001010",
39347 => "110010011100101011000100",
39348 => "110000111011110110010100",
39349 => "110000001100011010011110",
39350 => "110001001110000001110110",
39351 => "110100000001000111110101",
39352 => "110110110111001110101011",
39353 => "111001000010010010010010",
39354 => "111011100100101011011000",
39355 => "111111100010110000010111",
39356 => "000100111011100010010000",
39357 => "001010110010111111101100",
39358 => "001111100110010000011110",
39359 => "010001000011010100010110",
39360 => "001110000101100000011010",
39361 => "001000011101100110011110",
39362 => "000010011101111111010011",
39363 => "111100100110110110000000",
39364 => "110101111111110111001000",
39365 => "101110011000010010001100",
39366 => "100111100100010011010110",
39367 => "100100011111000110111101",
39368 => "100110011110101000100101",
39369 => "101011011100100010001010",
39370 => "110000110100101111110000",
39371 => "110110101111111101011110",
39372 => "111100110100110100010001",
39373 => "000001110000011111011000",
39374 => "000110010010000100100001",
39375 => "001010010011110101100101",
39376 => "001100011111010100001000",
39377 => "001101000011010100000100",
39378 => "001100010100000101111100",
39379 => "001010101101010000111000",
39380 => "001001011001110110010000",
39381 => "001000000100011000100110",
39382 => "000101011011000000001011",
39383 => "000001010101110110110101",
39384 => "111100110110011100010000",
39385 => "111000011111101100000100",
39386 => "110100010001011111101010",
39387 => "110001011011110100100000",
39388 => "110000001100111011100110",
39389 => "101111001010111011101100",
39390 => "101111010110000010000110",
39391 => "110001110001010111001000",
39392 => "110101011000010010111010",
39393 => "111001110000000001110101",
39394 => "111101100100001101100000",
39395 => "111111111001110011110111",
39396 => "000010110111001010111011",
39397 => "000110001011011000110010",
39398 => "000111000010001101001010",
39399 => "000101010100000110101011",
39400 => "000010000010110011000101",
39401 => "111101110100001101010111",
39402 => "111001111000010111001001",
39403 => "110110111010001110110101",
39404 => "110100110010010000000010",
39405 => "110100001110010100110100",
39406 => "110110001100010110101110",
39407 => "111001011011100010110001",
39408 => "111011100110100111100101",
39409 => "111100111011001100101011",
39410 => "111110100100010111010010",
39411 => "111111110101110011011110",
39412 => "111111100110001010100100",
39413 => "111101011110000110110011",
39414 => "111010011110001001010111",
39415 => "111000100101001001111000",
39416 => "111000000111111111010110",
39417 => "111000010010010101101001",
39418 => "111001010100101111100001",
39419 => "111011100100100011101100",
39420 => "111110111001101011110000",
39421 => "000011001011010000110110",
39422 => "000111010011100000101101",
39423 => "001001101011011011010010",
39424 => "001001111100110001111100",
39425 => "001000111111010110010001",
39426 => "000111011110000110010010",
39427 => "000101010110100000000000",
39428 => "000010110111011101111000",
39429 => "000001000111000010110000",
39430 => "000000110010010100110101",
39431 => "000001001011101000100110",
39432 => "000001011011101110011011",
39433 => "000010000110000110111001",
39434 => "000011110110110110001101",
39435 => "000101100100110000010010",
39436 => "000110001000110000101001",
39437 => "000110010100001101101100",
39438 => "000110010100111000111000",
39439 => "000101011010001000001110",
39440 => "000100000110100001011011",
39441 => "000011000110010010111010",
39442 => "000010100011100111011111",
39443 => "000011000001100010011010",
39444 => "000011110101101100001000",
39445 => "000011111010011010011011",
39446 => "000011111101101010011010",
39447 => "000100010110000100000000",
39448 => "000011111100111000101100",
39449 => "000010001011011001011010",
39450 => "111111010010000110101111",
39451 => "111011110111011001001000",
39452 => "111000010101111011111010",
39453 => "110100100110001101110011",
39454 => "110000110000011010000000",
39455 => "101101110110010110011100",
39456 => "101101000010111011010110",
39457 => "101110010111100001110110",
39458 => "110001010011111001100000",
39459 => "110101011100111100111001",
39460 => "111001001011011010110111",
39461 => "111011100001111011110001",
39462 => "111110000110001110100101",
39463 => "000001011111000010010000",
39464 => "000100000101111110100011",
39465 => "000101000110001001101100",
39466 => "000101010011000100111000",
39467 => "000110001000100100110101",
39468 => "000111111001000101000011",
39469 => "001001011000101010110010",
39470 => "001010000011111000010011",
39471 => "001010011010011101111100",
39472 => "001011000111010100110100",
39473 => "001100001110010111111100",
39474 => "001100101101111011000010",
39475 => "001100000110001100111110",
39476 => "001011000001101010110001",
39477 => "001010000110100100011110",
39478 => "001001100110000010111110",
39479 => "001001000011101011001011",
39480 => "001000001010001111011000",
39481 => "001000000100111010010110",
39482 => "001001101001110100100001",
39483 => "001011111011110110010001",
39484 => "001101101010010101010110",
39485 => "001110100000011110111000",
39486 => "001110100010111010010100",
39487 => "001101011110010100001000",
39488 => "001011100000100001001100",
39489 => "001001011100011001000010",
39490 => "000111011101011100001111",
39491 => "000110010110100101101001",
39492 => "000111010111001001100000",
39493 => "001001011010110101110110",
39494 => "001010011010110101011101",
39495 => "001010001110010111011010",
39496 => "001001111100010001100100",
39497 => "001001101101100000111110",
39498 => "001000101001101000010000",
39499 => "000110011110011010010001",
39500 => "000011010111101010000000",
39501 => "111110110110010001100010",
39502 => "111000101101001011111111",
39503 => "110010010001000011111110",
39504 => "101101111000011001100100",
39505 => "101100111110100110111100",
39506 => "101110110000110101010010",
39507 => "110001100111000110000010",
39508 => "110100010111110111100110",
39509 => "110110011110101010010100",
39510 => "111000011011101110111011",
39511 => "111011001100110001010010",
39512 => "111110110001001001010111",
39513 => "000010001001100011110101",
39514 => "000101000001001010110010",
39515 => "001000010110100111010100",
39516 => "001100000111111000111110",
39517 => "001110111100000010101100",
39518 => "001111111111010000011100",
39519 => "001110011011100100110100",
39520 => "001010010100111110001100",
39521 => "000110000010101101011100",
39522 => "000010111100101100110100",
39523 => "000000011111010011000001",
39524 => "111110010111010010011110",
39525 => "111100000110010010001110",
39526 => "111001000101110101101000",
39527 => "110101110000000000010101",
39528 => "110011001101101011010000",
39529 => "110010010101000110011110",
39530 => "110010110011011111100110",
39531 => "110011101111010111001100",
39532 => "110100011111101100110110",
39533 => "110101110010111101000011",
39534 => "111001110011010011001001",
39535 => "000000001111011010001101",
39536 => "000110010110010111100000",
39537 => "001011011001111111101110",
39538 => "001111100001000000001010",
39539 => "010010001101010110011100",
39540 => "010100000111011011100000",
39541 => "010100100100011110100010",
39542 => "010001110001101001101000",
39543 => "001100011110010010000110",
39544 => "000110010111011111011110",
39545 => "000000000101100110001100",
39546 => "111010000111100001100100",
39547 => "110101000100101101111110",
39548 => "110001011111100100111010",
39549 => "101111001111101000100110",
39550 => "101101100100101100110000",
39551 => "101100010010110011111110",
39552 => "101100011010011100100010",
39553 => "101111001000101011001110",
39554 => "110011000010111100000110",
39555 => "110101001111010101000000",
39556 => "110110000110111100001010",
39557 => "110111001111000011100110",
39558 => "110111111101100101101110",
39559 => "111000011100010110000111",
39560 => "111001011110100101011000",
39561 => "111010011010000111110101",
39562 => "111011100000111000110000",
39563 => "111101011000001010111111",
39564 => "111110101110011011100011",
39565 => "111110100101010101000101",
39566 => "111101000110010001111010",
39567 => "111010110010010100110110",
39568 => "111001000010011111000011",
39569 => "111000101111011100101000",
39570 => "111000101001010101100101",
39571 => "110111001011011010011110",
39572 => "110101001001011001000100",
39573 => "110100110001010000111111",
39574 => "110110001001100110000111",
39575 => "110111011110001110001011",
39576 => "111000000110010001000011",
39577 => "111001000001111101101100",
39578 => "111011001111011101001011",
39579 => "111101100011110100111010",
39580 => "111110000001110011100001",
39581 => "111110110000001111010110",
39582 => "000011000001100111101011",
39583 => "001000101111111110100110",
39584 => "001100100110111010111110",
39585 => "001111010011010110101110",
39586 => "010010000110000001001100",
39587 => "010100001000001101101100",
39588 => "010011111100100110001010",
39589 => "010001100110001100000100",
39590 => "001110110110110101101110",
39591 => "001100100010010111111000",
39592 => "001001111000100010111011",
39593 => "000110101111011010010111",
39594 => "000011110010100111110010",
39595 => "000001100000000001000010",
39596 => "111111100100000110011100",
39597 => "111110000111100111100010",
39598 => "111110100101001111011001",
39599 => "000001000001110000001100",
39600 => "000011110100110101101001",
39601 => "000110001000111011111101",
39602 => "000111101010001110100010",
39603 => "001000010010100000101010",
39604 => "000111111001010101011011",
39605 => "000101110010101000111100",
39606 => "000011001010111111100111",
39607 => "000001111101000010101000",
39608 => "000000101011011011110101",
39609 => "111101101000111101000110",
39610 => "111010101001110000010111",
39611 => "111001100100110110101010",
39612 => "111000110100111000000100",
39613 => "110101111111001110011010",
39614 => "110010000000010101000100",
39615 => "101110011001111100000000",
39616 => "101001110000010100001110",
39617 => "100100101110011011000000",
39618 => "100010101111011011011111",
39619 => "100011010111101000011011",
39620 => "100100001110011110111100",
39621 => "100101000100111001000101",
39622 => "100110010100100111101101",
39623 => "101001100101110010001100",
39624 => "101111110111001000111110",
39625 => "110110001110100001011111",
39626 => "111010100001001110011100",
39627 => "111101101100111011000011",
39628 => "000000010100101110111111",
39629 => "000010001000110010100000",
39630 => "000010011111101101011000",
39631 => "000001011000001010000011",
39632 => "000001000000111110111110",
39633 => "000010010100000100000101",
39634 => "000011010011110100101011",
39635 => "000011001100010101110110",
39636 => "000010110100101110110101",
39637 => "000010101110110100010110",
39638 => "000010100000010000000010",
39639 => "000001100101001101100011",
39640 => "000000111111011100110000",
39641 => "000001101010010110111010",
39642 => "000010110100111010111110",
39643 => "000100100101101010010100",
39644 => "000111011110101001000011",
39645 => "001010101001010110110110",
39646 => "001101011001100011100100",
39647 => "001111101001110010111100",
39648 => "010001100100110010111000",
39649 => "010011010001111000001010",
39650 => "010100001110101000101100",
39651 => "010100111000000000011100",
39652 => "010110010001111010110000",
39653 => "010111101111000000010110",
39654 => "011000000110000001101100",
39655 => "010111000010011101010010",
39656 => "010100101100011010000010",
39657 => "010001110100001101010000",
39658 => "001110110111111011010010",
39659 => "001100001000000011010100",
39660 => "001010000011000011011100",
39661 => "000111111111101011011000",
39662 => "000101000100100000101111",
39663 => "000001110101100001000010",
39664 => "111111100111111101000101",
39665 => "111111000011011001100000",
39666 => "111111000100010111111000",
39667 => "111110110110100100111111",
39668 => "111111011000011101000110",
39669 => "000000110110101000000010",
39670 => "000010010011100101110000",
39671 => "000011010110101010100001",
39672 => "000011111000001101110111",
39673 => "000100100000010010100010",
39674 => "000101011101000101010111",
39675 => "000101000101100100110101",
39676 => "000011100010111000100100",
39677 => "000011000100101110110000",
39678 => "000011001111110011001001",
39679 => "000001100010011000100111",
39680 => "111101001110011111101011",
39681 => "111000010000111101001001",
39682 => "110101000111100011101000",
39683 => "110011111011100011100000",
39684 => "110011010010101110100000",
39685 => "110010100100100111111010",
39686 => "110001110100100011100010",
39687 => "110010000000110001110110",
39688 => "110100101011100011111010",
39689 => "111001110011001111111100",
39690 => "000000000110100000110000",
39691 => "000110010111111111101011",
39692 => "001011000111110011000110",
39693 => "001101000111111101010010",
39694 => "001100100101001010100010",
39695 => "001010001111001010110001",
39696 => "000110000010111010111101",
39697 => "111111111110111101011001",
39698 => "111001000001011010110010",
39699 => "110010010111111000001000",
39700 => "101101110101100010101010",
39701 => "101101010110110110101000",
39702 => "110000000010001000101100",
39703 => "110011011011000110101000",
39704 => "110110111100100011110100",
39705 => "111010011000000010101111",
39706 => "111101011001111101001000",
39707 => "000000110010010001011110",
39708 => "000011100101010111100011",
39709 => "000011110010110010001111",
39710 => "000010100101010001100101",
39711 => "000010000000000111110110",
39712 => "000001011000111110110100",
39713 => "000000010010101100100000",
39714 => "111111111001000111001010",
39715 => "000000000011000111011011",
39716 => "000000001001010111001110",
39717 => "000000111110011100011111",
39718 => "000001101101011010011010",
39719 => "000000010001101100100001",
39720 => "111101011110001000001000",
39721 => "111010100111011111010111",
39722 => "110111011100111000011001",
39723 => "110100110001000111100010",
39724 => "110010100011101010010110",
39725 => "101111101101001111111110",
39726 => "101110101000111010100000",
39727 => "110001101111000111000000",
39728 => "110110110010110101000000",
39729 => "111100010111101110011100",
39730 => "000011001100101010001000",
39731 => "001001110011111010100110",
39732 => "001110010001010100011010",
39733 => "010000011001011101000000",
39734 => "001111111000101010101010",
39735 => "001100111100001001010100",
39736 => "001000111111100000001100",
39737 => "000100001010001000010010",
39738 => "111110000010010000001000",
39739 => "111000101011011110010000",
39740 => "110110000100110001011100",
39741 => "110101010010110111000010",
39742 => "110101001000001011101111",
39743 => "110101100011100001011010",
39744 => "110110111100010001110000",
39745 => "111010001111111001010111",
39746 => "111111011000001101011101",
39747 => "000100101100101111010000",
39748 => "001001111011101000110010",
39749 => "001111101111100111000100",
39750 => "010101101011110011100100",
39751 => "011010011001010011100101",
39752 => "011100001111000100000101",
39753 => "011011100111000001100001",
39754 => "011010100101101101011010",
39755 => "011000011100111100100111",
39756 => "010100000000010100000100",
39757 => "001111010010110110011110",
39758 => "001011010000001100001000",
39759 => "000111000011001010000000",
39760 => "000100000001010001111110",
39761 => "000011010110011111010010",
39762 => "000100000111001100001010",
39763 => "000101011111001111101100",
39764 => "000110101111010000001010",
39765 => "000111001000001000100110",
39766 => "000111000011111101111001",
39767 => "000110101011110101000000",
39768 => "000101000000100111000000",
39769 => "000010000001001001100110",
39770 => "111110110110011101001111",
39771 => "111011001011111011111100",
39772 => "110110000011100010010001",
39773 => "110000100110010111111000",
39774 => "101011100100001111001110",
39775 => "100110000011101101101000",
39776 => "100010001011000101110011",
39777 => "100011010011011111100101",
39778 => "100111111110000101101101",
39779 => "101100100000011000011010",
39780 => "101111100101001010110100",
39781 => "110001010010100010100010",
39782 => "110010100010000001000010",
39783 => "110011110010011111111000",
39784 => "110100000000110111000100",
39785 => "110010110110100011100110",
39786 => "110000100110111010110100",
39787 => "101101010011101111110100",
39788 => "101010101110101110100000",
39789 => "101010101001110100000010",
39790 => "101011111101101010100100",
39791 => "101101101011101111001000",
39792 => "110000101100010010110110",
39793 => "110100110010110001110100",
39794 => "111000000100111010110110",
39795 => "111001011000101001111001",
39796 => "111001001011000010100111",
39797 => "110111110111011000110001",
39798 => "110101111101110000111010",
39799 => "110101011101100001101011",
39800 => "110111010101101100100111",
39801 => "111010010001110011000101",
39802 => "111101111101010111000101",
39803 => "000010010111001101010100",
39804 => "000101110001111110101110",
39805 => "000111111100000001101010",
39806 => "001010001011011010100000",
39807 => "001100001111011011010100",
39808 => "001100110110010100100000",
39809 => "001011100011110011011000",
39810 => "001001011001011000110110",
39811 => "000111110110000101011100",
39812 => "000110101111000110000010",
39813 => "000101100110100000001110",
39814 => "000101010000110101000010",
39815 => "000101111101001111011111",
39816 => "000111100011100010011100",
39817 => "001010100111010010010001",
39818 => "001110110111111000111000",
39819 => "010010110000110110111000",
39820 => "010100001101101111101000",
39821 => "010010101010011101100110",
39822 => "010000010100101100010100",
39823 => "001110101100100101100010",
39824 => "001101000111110110101000",
39825 => "001011110010000110000010",
39826 => "001010111010011110100100",
39827 => "001001101100011110101100",
39828 => "001000010110000001011100",
39829 => "000111001111011101011110",
39830 => "000101101111110010001000",
39831 => "000011110111000011111101",
39832 => "000010010100001010010101",
39833 => "000001100110110101100100",
39834 => "000001110101101001001111",
39835 => "000010110110010001111000",
39836 => "000100100110010010111000",
39837 => "000110110100010010000111",
39838 => "001001000000100000101100",
39839 => "001011000000100111011100",
39840 => "001100001011010000011110",
39841 => "001011100111011110110110",
39842 => "001001011101111001101000",
39843 => "000110001010111011111110",
39844 => "000010000100011001101001",
39845 => "111101111001001100100101",
39846 => "111010011000010101010000",
39847 => "111000010111110110001001",
39848 => "111000100010100011100001",
39849 => "111010001010110100000000",
39850 => "111011111100110000111010",
39851 => "111101101011111111010110",
39852 => "111111110110011111100110",
39853 => "000010000111111111101011",
39854 => "000011110001110001110110",
39855 => "000100101100101011110001",
39856 => "000100010011110101110101",
39857 => "000001100001001000101001",
39858 => "111101001010100110000010",
39859 => "111001000010110100100000",
39860 => "110101000101011110010010",
39861 => "110000111110111001100000",
39862 => "101101100111101011001000",
39863 => "101011000110110001111110",
39864 => "101000111001001011011110",
39865 => "100111101110110011111101",
39866 => "101000110110110100011000",
39867 => "101100001101100101100110",
39868 => "110000111111100100000100",
39869 => "110110100011000110010001",
39870 => "111100001010011111011001",
39871 => "000001011110001101111111",
39872 => "000110001101010110011101",
39873 => "001000110111000100011111",
39874 => "001000000110110111101010",
39875 => "000100111100001001100111",
39876 => "000001010011111010011110",
39877 => "111110011111110000100001",
39878 => "111100100000001101000100",
39879 => "111001110101011000000010",
39880 => "110110000001010010010110",
39881 => "110011010111110011110010",
39882 => "110011100111010111100010",
39883 => "110101101001011001111001",
39884 => "111000001101101011011000",
39885 => "111011000111001001100111",
39886 => "111101100110010110110100",
39887 => "111111010001101100000011",
39888 => "000000111011111011110010",
39889 => "000010010111001011111101",
39890 => "000010110001000110001110",
39891 => "000010101011000010000111",
39892 => "000010000111011110010111",
39893 => "000001000011100000011000",
39894 => "000001010110000101011110",
39895 => "000011101011110011001110",
39896 => "000110100110110110101000",
39897 => "001001100010101001101000",
39898 => "001011110001100101111100",
39899 => "001011101011111001110101",
39900 => "001001011111011111001100",
39901 => "000110101110110101110010",
39902 => "000011111011101110001111",
39903 => "000000111010110110001010",
39904 => "111101111101111101011110",
39905 => "111100001110111110111100",
39906 => "111101000010001111111101",
39907 => "000000011101100010000101",
39908 => "000100110000101100100101",
39909 => "001000000001100100101110",
39910 => "001010111001100110011111",
39911 => "001110101101001011000000",
39912 => "010001100110010011010110",
39913 => "010000111110001000101100",
39914 => "001101001110110000110110",
39915 => "001000111100000110110100",
39916 => "000110010111111011011100",
39917 => "000101000101101001010101",
39918 => "000011001010111101101101",
39919 => "000001101001000100010111",
39920 => "000010100111001110000110",
39921 => "000101001001110011000100",
39922 => "000111010010111011010111",
39923 => "001000011111000010110010",
39924 => "001001011001111010101110",
39925 => "001010101111000010000010",
39926 => "001010111111010110110000",
39927 => "001000100100001010100010",
39928 => "000101001101111010010101",
39929 => "000010110011000001111111",
39930 => "111111111000001110101001",
39931 => "111011000000111100001110",
39932 => "110101011111101010101000",
39933 => "110001000000011001001110",
39934 => "101101010010011111111100",
39935 => "101001111111010011111000",
39936 => "101000101100101101110010",
39937 => "101010101010110111101100",
39938 => "101110010011100111000100",
39939 => "110001000011101110100010",
39940 => "110010111101010011110110",
39941 => "110110001010011000001010",
39942 => "111010101001000010111010",
39943 => "111101111110001001100101",
39944 => "111111101010000100001111",
39945 => "000000110110000001100010",
39946 => "000001001001101010110100",
39947 => "111111101001011001000110",
39948 => "111100100111111110111111",
39949 => "111001001011100001010010",
39950 => "110110010001001001101100",
39951 => "110100001110111100000001",
39952 => "110011011111110111110010",
39953 => "110100010101101100100100",
39954 => "110101110100110111000110",
39955 => "110111010100010110110101",
39956 => "111001010001101001111001",
39957 => "111011010101101101110111",
39958 => "111100100111110010000011",
39959 => "111101010101101001110010",
39960 => "111110000111111011010001",
39961 => "111111000101011110111010",
39962 => "111111111101001010111100",
39963 => "000000011000101111110010",
39964 => "000000010111000001001101",
39965 => "000000011011101100000000",
39966 => "000001001110011001111100",
39967 => "000010100010010011101111",
39968 => "000011100111001100011100",
39969 => "000100001100010110101001",
39970 => "000100100111100010100000",
39971 => "000101011110010010010111",
39972 => "000110110001110010110000",
39973 => "000111011010110111111110",
39974 => "000111000101100011010011",
39975 => "000110111110010110110000",
39976 => "000111001111100011001001",
39977 => "000111010010011100100000",
39978 => "000111011110001011101000",
39979 => "000111010111001100110111",
39980 => "000101111000010101000100",
39981 => "000100000000110100101000",
39982 => "000011010101110101111100",
39983 => "000011101111010010100101",
39984 => "000100110101111010101001",
39985 => "000110100111110010101011",
39986 => "001000010111000111111001",
39987 => "001001011011111100010000",
39988 => "001001101010111001010001",
39989 => "001000110011001111000101",
39990 => "000111100001111111111011",
39991 => "000110111111000011101110",
39992 => "000110011011011110110010",
39993 => "000101001011000001011110",
39994 => "000100111010011100010110",
39995 => "000110100001111110011100",
39996 => "001000010011010011010100",
39997 => "001001001000010010011100",
39998 => "001001001011011111101010",
39999 => "000111111001110100111011",
40000 => "000101000101111110101011",
40001 => "000010001010100101100111",
40002 => "000000011101011011010110",
40003 => "000000000111010110010110",
40004 => "000000101000101110001101",
40005 => "000001000101000000111111",
40006 => "000000111101011010000011",
40007 => "000001010001110110110100",
40008 => "000010110001010110011010",
40009 => "000100101011111101011100",
40010 => "000110011011011100010001",
40011 => "000111110111110010111000",
40012 => "001000100010100000010000",
40013 => "001000001111101011010110",
40014 => "000111011010000101100110",
40015 => "000110100111011101000101",
40016 => "000110000000110010001101",
40017 => "000100111010100101101010",
40018 => "000011011010100000100011",
40019 => "000010101111100011011111",
40020 => "000010110001100011100100",
40021 => "000010000111110111111110",
40022 => "000000100101110111001101",
40023 => "111111011000000110001110",
40024 => "111111101100111101101000",
40025 => "000001100000110101011100",
40026 => "000011011110010101101100",
40027 => "000100000111101111110100",
40028 => "000010011100010101100001",
40029 => "111110101111011010001100",
40030 => "111010011000000011110001",
40031 => "110101110100100110100100",
40032 => "110000110111100110011110",
40033 => "101011001110000011011110",
40034 => "100101001001110001100100",
40035 => "100001011001000111110101",
40036 => "100001010111110011111001",
40037 => "100010100100110001101101",
40038 => "100101001100100011000111",
40039 => "101011010001011111111000",
40040 => "110001111000111111110000",
40041 => "110111010101101010111010",
40042 => "111110110000001001000101",
40043 => "000111101001111001100011",
40044 => "001101111001100010011000",
40045 => "010000000111111110101010",
40046 => "001111100110000001011100",
40047 => "001101110111011110111100",
40048 => "001011011000101110010011",
40049 => "000111111011010011110011",
40050 => "000100000111011001010000",
40051 => "111111111111001110001101",
40052 => "111011001111110010000110",
40053 => "110111000111100111111000",
40054 => "110100100101101000110110",
40055 => "110011111000001001101010",
40056 => "110100110010101111011110",
40057 => "110101110000010101101010",
40058 => "110110001101111100111110",
40059 => "110111010101011011110010",
40060 => "111001010100010100111110",
40061 => "111100010010111100000111",
40062 => "000000011010100010001011",
40063 => "000101001100010011110000",
40064 => "001011011010000011110101",
40065 => "010010100110100001010010",
40066 => "010111011100111000110100",
40067 => "011000111101010100111001",
40068 => "011000111100111101000011",
40069 => "010111110100111100100110",
40070 => "010100110000010111000000",
40071 => "010000000010001111000010",
40072 => "001011011010001011110100",
40073 => "000111011001111111111010",
40074 => "000010010000011110010101",
40075 => "111100010011011101101011",
40076 => "111000101011001101110100",
40077 => "111000000010101001100111",
40078 => "111000000001000000101100",
40079 => "110111010011010110011011",
40080 => "110111101001000100010000",
40081 => "111010100100101101100011",
40082 => "111110000111111000011010",
40083 => "000000110100100100100001",
40084 => "000100001010110011100000",
40085 => "000111111010001000001111",
40086 => "001010011001001111110100",
40087 => "001011110110101001110000",
40088 => "001100100111100001110010",
40089 => "001100011101000010011000",
40090 => "001010001011110010011101",
40091 => "000100000001100000110011",
40092 => "111011100001100110010000",
40093 => "110011000010101100100110",
40094 => "101010001110111010111010",
40095 => "100011010100000101111010",
40096 => "100001010100110101000001",
40097 => "100001101010100010001111",
40098 => "100001110001010110010001",
40099 => "100011011101101101111101",
40100 => "100111111100000001001101",
40101 => "101110111110001111101100",
40102 => "111000000011011111010100",
40103 => "000000011001110000001001",
40104 => "000101000110000101111111",
40105 => "000110101111110111000010",
40106 => "000111001111000011000011",
40107 => "000110000111100011000011",
40108 => "000010101101110110101000",
40109 => "111111000000110001000010",
40110 => "111101000001101010111010",
40111 => "111100100011011010111100",
40112 => "111101010001110100111111",
40113 => "111111001100110101001100",
40114 => "000001010101000000110100",
40115 => "000010101001100111010100",
40116 => "000010110100110111011111",
40117 => "000001100110110110000100",
40118 => "111111001010111101011110",
40119 => "111100011110100001000110",
40120 => "111010100010101101001100",
40121 => "111001110100110111110001",
40122 => "111010010101100111010001",
40123 => "111011100101000010100101",
40124 => "111100101001111010100001",
40125 => "111101010111110110111101",
40126 => "111110011001111101100101",
40127 => "111111111010110110000011",
40128 => "000001001011111110101011",
40129 => "000001110000110111101000",
40130 => "000010100011101000101110",
40131 => "000100110010100110011000",
40132 => "000111100110000100110101",
40133 => "001000110010000110011011",
40134 => "000111111101001001001010",
40135 => "000110011000100110110001",
40136 => "000100110011000100110001",
40137 => "000011000110100000111010",
40138 => "000001010001011111010101",
40139 => "111111010000100010011000",
40140 => "111100011011011010011010",
40141 => "111000101101111110110011",
40142 => "110101101110110000111110",
40143 => "110100111101100001001111",
40144 => "110110000100110100100000",
40145 => "110111110001111111010100",
40146 => "111001010101101010111110",
40147 => "111010110011000000110110",
40148 => "111011100101110101011101",
40149 => "111010101110001110001010",
40150 => "111001000110101111011110",
40151 => "111000011110011001011000",
40152 => "111001000101011100010111",
40153 => "111011000011111101101101",
40154 => "111110011010001011101110",
40155 => "000001111000001010111110",
40156 => "000100111001111011011000",
40157 => "000111101010110101000001",
40158 => "001001001100010110111100",
40159 => "001000110111010010101111",
40160 => "000111101100010010001001",
40161 => "000110011001011111100000",
40162 => "000100100010001011001011",
40163 => "000001110010101010110010",
40164 => "111110100110001001100001",
40165 => "111011011110001010111010",
40166 => "111001001010010000101111",
40167 => "111000100110110011101100",
40168 => "111001110000111101101100",
40169 => "111100001011000110001101",
40170 => "000000000001001101010110",
40171 => "000100110100011010111111",
40172 => "001001010010100001010010",
40173 => "001100101001001001110100",
40174 => "001110100100100000100000",
40175 => "001111101110011001111010",
40176 => "010001001110001100110100",
40177 => "010010100000001101000010",
40178 => "010010101010100111101010",
40179 => "010010011100100111000110",
40180 => "010010001100100100111100",
40181 => "010001000111011111010100",
40182 => "001111011000110011000110",
40183 => "001101111110111011000100",
40184 => "001100110100011010011000",
40185 => "001011001001010011010011",
40186 => "001001001110111000000101",
40187 => "001000000101011100100010",
40188 => "000111110000000100011110",
40189 => "000111100010110000000001",
40190 => "000111100101110000001101",
40191 => "001000011010001001110010",
40192 => "001001101011000111011000",
40193 => "001010110010110101100011",
40194 => "001011001000110110101100",
40195 => "001001011101010010010000",
40196 => "000101101001101000000110",
40197 => "000001011100011110010001",
40198 => "111101011011000010101011",
40199 => "111001000111011111001011",
40200 => "110101100000100011110010",
40201 => "110011010101110111110110",
40202 => "110010010100110100010100",
40203 => "110011010100001010111100",
40204 => "110110110011001100101000",
40205 => "111011001100011001100110",
40206 => "111111010001000101111001",
40207 => "000010111100011111101010",
40208 => "000101100110110111111011",
40209 => "000101111011010111111000",
40210 => "000011000011101010100001",
40211 => "111101111011011011000010",
40212 => "111000111011111100010100",
40213 => "110101001010101111010110",
40214 => "110001100011101100000100",
40215 => "101110001101000011010010",
40216 => "101101100011011001010010",
40217 => "110000011111100000000000",
40218 => "110101001001001111001001",
40219 => "111010011000011011000010",
40220 => "111111111110000111110101",
40221 => "000100100011001101000110",
40222 => "000111011000001101001111",
40223 => "001001000011100111100101",
40224 => "001001000101010100110011",
40225 => "000110010011100001011111",
40226 => "000001100000100000100000",
40227 => "111100110101111010100101",
40228 => "111001100010000110100000",
40229 => "111000000011001000010111",
40230 => "111001000010010101111010",
40231 => "111100010101101100010100",
40232 => "000001000110101010100010",
40233 => "000110101001001011001010",
40234 => "001010111101101101101000",
40235 => "001011111100001111101100",
40236 => "001010110110101011010111",
40237 => "001010001001110110110010",
40238 => "001001100111100011001100",
40239 => "000111101011010110000111",
40240 => "000100001000111111100010",
40241 => "000001010010100010101011",
40242 => "000001011111101011111100",
40243 => "000011000011011101001001",
40244 => "000010110011100010101000",
40245 => "000001100110000001111110",
40246 => "000001011010110111100101",
40247 => "000000111011111010101100",
40248 => "111110101000101101101110",
40249 => "111100001011101001001110",
40250 => "111011010111101000011101",
40251 => "111011001101001111010000",
40252 => "111001111010010000000100",
40253 => "110111011001010000100011",
40254 => "110100101101101110011100",
40255 => "110010100111011110001010",
40256 => "110001100110111101001110",
40257 => "110010101000001101001000",
40258 => "110101101111111111101110",
40259 => "111000110111010101011000",
40260 => "111010010101100000011100",
40261 => "111011010010110100000100",
40262 => "111101001010010101111000",
40263 => "111111011010100001100110",
40264 => "000000100100111110011000",
40265 => "000000000101110110110110",
40266 => "111110111101101111010000",
40267 => "111110000111001111011111",
40268 => "111100111111010111101001",
40269 => "111010101010110001001011",
40270 => "110111010101000011001010",
40271 => "110100101001110000001000",
40272 => "110011111001101000110110",
40273 => "110100001101111101110110",
40274 => "110100111110010110110110",
40275 => "110110101100011000010011",
40276 => "111000111011000000001100",
40277 => "111011001110010001110001",
40278 => "111110000110110000011010",
40279 => "000001100100101100000110",
40280 => "000101011110101101111101",
40281 => "001001011011010100100010",
40282 => "001100001100100110101010",
40283 => "001101000000010111011110",
40284 => "001011100101010111110011",
40285 => "000111111111101010001100",
40286 => "000010111110000001100011",
40287 => "111101011001010100010000",
40288 => "111000111001000001101110",
40289 => "110110111010101100100100",
40290 => "110110111000101101001100",
40291 => "111000010010001110000011",
40292 => "111011010010100010011010",
40293 => "111110011111000001110101",
40294 => "000000100011011010111101",
40295 => "000001101111011011110100",
40296 => "000010001110100111000100",
40297 => "000010000001111110111010",
40298 => "000000111010010000010111",
40299 => "111110010111001100001000",
40300 => "111010111001011010001000",
40301 => "110111010101100111101100",
40302 => "110100001100111111111110",
40303 => "110010101000110011011010",
40304 => "110011011001110110111100",
40305 => "110101101100111001011110",
40306 => "111000011111011101010011",
40307 => "111011101001010000000001",
40308 => "111110011110010111111001",
40309 => "111111000010001001101000",
40310 => "111101001101100110000100",
40311 => "111011010101011011111011",
40312 => "111010000101001100101000",
40313 => "111000011111011110101110",
40314 => "110110111001000111001010",
40315 => "110110000010000010010100",
40316 => "110110001110101010110101",
40317 => "110111100000110100000000",
40318 => "111000111111100101111010",
40319 => "111010011111010010001001",
40320 => "111100111000101110001101",
40321 => "111111101001011001000101",
40322 => "000001010111000011101111",
40323 => "000001100001011001111001",
40324 => "000000010011101011001011",
40325 => "111110011110001000101101",
40326 => "111100111101111100101010",
40327 => "111100001000001111100110",
40328 => "111011110111101111110001",
40329 => "111100100010011111111000",
40330 => "111110011110001011001001",
40331 => "000000101001001111010000",
40332 => "000001111000111101000110",
40333 => "000010101101110011100100",
40334 => "000011101101100000110111",
40335 => "000100100010101100011100",
40336 => "000101000110111001000100",
40337 => "000101100001011100000010",
40338 => "000110000000100001011101",
40339 => "000110111011100000001001",
40340 => "001000001101110101010110",
40341 => "001001011110110011111001",
40342 => "001010000010111001101011",
40343 => "001001100110000011010111",
40344 => "001001000011101001111100",
40345 => "001001001010001000111111",
40346 => "001001101110010010101101",
40347 => "001010011011110111011111",
40348 => "001010110001101001001001",
40349 => "001010101101011001011000",
40350 => "001010111010011001100011",
40351 => "001011101111011100010011",
40352 => "001100110110011100100110",
40353 => "001101001111010011001010",
40354 => "001100110101111001110100",
40355 => "001101001110001001011100",
40356 => "001110010001111000000000",
40357 => "001110001110100011111110",
40358 => "001101011001101101100000",
40359 => "001101000011010110001110",
40360 => "001100110111100000111010",
40361 => "001100001100011111011100",
40362 => "001010101010000110111000",
40363 => "001000010010010101001000",
40364 => "000101011001001001010100",
40365 => "000001111111101110000100",
40366 => "111110101000111001010000",
40367 => "111011101001001010001000",
40368 => "111000101001001110010110",
40369 => "110110011000000011000000",
40370 => "110101100001011110100101",
40371 => "110101110001000111011010",
40372 => "110111010100011111001000",
40373 => "111001111010010000000010",
40374 => "111100100000100100000001",
40375 => "111111010000111011101010",
40376 => "000010011100100001101000",
40377 => "000101010011100111100101",
40378 => "000111011001001011101010",
40379 => "001000101011101101000100",
40380 => "001000111101010111101110",
40381 => "000111111001110111101001",
40382 => "000101011110100100001111",
40383 => "000001110101110010010100",
40384 => "111101101110001100000011",
40385 => "111011010101010100100100",
40386 => "111010110011101100010101",
40387 => "111000101100001110000011",
40388 => "110100101100110000110001",
40389 => "110001110111110110101100",
40390 => "110001011111110101010000",
40391 => "110100000001101100101110",
40392 => "110111110011001111100010",
40393 => "111001100100110101101100",
40394 => "111010001110111111110100",
40395 => "111100001000001001100101",
40396 => "111111000100111010110010",
40397 => "000011010001000011101111",
40398 => "001000101111110100000000",
40399 => "001110011100111001101100",
40400 => "010100010101101110001010",
40401 => "011001100001110101010001",
40402 => "011011111011110010110100",
40403 => "011010111101100011010010",
40404 => "010110011010001110011110",
40405 => "001110111001101010010010",
40406 => "000110110001010100110100",
40407 => "111111001011101110000001",
40408 => "111000010101010111001100",
40409 => "110011001110100000001000",
40410 => "110000110001011101010110",
40411 => "110000010011000011101000",
40412 => "101111110001111101100100",
40413 => "101111001101110000110100",
40414 => "110000100000011000111000",
40415 => "110010111110010100001100",
40416 => "110100011011101111111010",
40417 => "110101100100100100110100",
40418 => "111000111100110110111010",
40419 => "111110111111001110001111",
40420 => "000100111111111000110000",
40421 => "001000101010111111110101",
40422 => "001011011000100110011110",
40423 => "001111000111110100000010",
40424 => "010010100011011010101010",
40425 => "010100000111010100001010",
40426 => "010011110110101011001110",
40427 => "010001001011111001110000",
40428 => "001011110010100110001100",
40429 => "000100111100000111001111",
40430 => "111110010010001110100001",
40431 => "111000100000011011010101",
40432 => "110100000011010010000000",
40433 => "110010001100110000000010",
40434 => "110011000111111011101100",
40435 => "110101101000111010001011",
40436 => "111000111100000111001110",
40437 => "111100101111011000011001",
40438 => "000001000101010011100110",
40439 => "000101000000001101100010",
40440 => "000111101101110101001000",
40441 => "001010010100101000101010",
40442 => "001100100001100001010110",
40443 => "001100110001000100110100",
40444 => "001011010011001010111000",
40445 => "001000101111001110011001",
40446 => "000101000010110101011111",
40447 => "000001000110010010000110",
40448 => "111110001101000101011100",
40449 => "111011001000001000000010",
40450 => "110101110100100111111110",
40451 => "110000100010110011111000",
40452 => "101110101101110110101000",
40453 => "101111011000011101100100",
40454 => "110000001000100000010000",
40455 => "110001000100100110110010",
40456 => "110011001000000100001000",
40457 => "110101101010110100001101",
40458 => "110111110110011101101110",
40459 => "111010010000010011011111",
40460 => "111100101111101101100110",
40461 => "111101011010100100011110",
40462 => "111011110001100010010000",
40463 => "111001100011110000010000",
40464 => "111000001011011000110000",
40465 => "110111100011001101001010",
40466 => "110110101111001110001001",
40467 => "110110000011001110011000",
40468 => "110110101001110101010011",
40469 => "110111101101111010100110",
40470 => "111000000100010110100011",
40471 => "110111110000111001000110",
40472 => "110110100001111010100100",
40473 => "110100111110000011110011",
40474 => "110100110000101101101011",
40475 => "110101111110111001111001",
40476 => "110111011101111101011010",
40477 => "111000111100000111100110",
40478 => "111010011000111010011001",
40479 => "111011010010100100011010",
40480 => "111100010001110010001001",
40481 => "111110010100000100101100",
40482 => "000000100011001011110001",
40483 => "000001111100010001000110",
40484 => "000010011110111000110011",
40485 => "000010011100110101110101",
40486 => "000001111100100010111010",
40487 => "000001010001101000010110",
40488 => "000001011010001100101000",
40489 => "000010100100001110010010",
40490 => "000011100010101101010001",
40491 => "000011001101111100111101",
40492 => "000010010100010000110100",
40493 => "000010011110101110010110",
40494 => "000010010001011111001000",
40495 => "111111100011100101011110",
40496 => "111100100000000011110010",
40497 => "111011011111010100111010",
40498 => "111100000101110011101010",
40499 => "111101101001100110111111",
40500 => "111111010100111000010001",
40501 => "000000011000110101010010",
40502 => "000000110111010110101110",
40503 => "000000101001001111010011",
40504 => "000000000101000001011000",
40505 => "000000000001011001011001",
40506 => "000001000010000001111010",
40507 => "000011000111111011000000",
40508 => "000101001101101110101111",
40509 => "000110011110100110101010",
40510 => "000111010111001011100001",
40511 => "000111111010001111000010",
40512 => "000111101010101111011101",
40513 => "000110100111000011001110",
40514 => "000101000001001000001010",
40515 => "000011001010001011111101",
40516 => "000000111111010001111110",
40517 => "111111001000001111100110",
40518 => "111110011111100110100000",
40519 => "111110000110010001100101",
40520 => "111100110011110101011101",
40521 => "111011101010100010001010",
40522 => "111011101111010111100111",
40523 => "111101000111011100111101",
40524 => "111111111000001010111111",
40525 => "000011011101011101001111",
40526 => "000110110100010010000010",
40527 => "001001100101001001001100",
40528 => "001100000010001100001010",
40529 => "001110010011111011000010",
40530 => "001111010110010000111010",
40531 => "001110001111111000100110",
40532 => "001011100100011100111000",
40533 => "000111101000111110100111",
40534 => "000010101110110010110100",
40535 => "111101011010010101100100",
40536 => "111000000100011101010011",
40537 => "110100000000100110100100",
40538 => "110010001010000110011010",
40539 => "110001110100101000101110",
40540 => "110010110000100110101000",
40541 => "110101110101011100000110",
40542 => "111011000010010100011111",
40543 => "000000110000111101000011",
40544 => "000101100010011000010010",
40545 => "001001000000101110000110",
40546 => "001100010001001110100110",
40547 => "001111101110111100100110",
40548 => "010001001010010011010110",
40549 => "001111101111101100010000",
40550 => "001101010110100101001010",
40551 => "001011001101010010010111",
40552 => "001001101000111001011101",
40553 => "001000110011110100011001",
40554 => "001001101001000110111111",
40555 => "001011011001101010000111",
40556 => "001011010000011010101110",
40557 => "001001100001101000111010",
40558 => "001000000010001111111111",
40559 => "000111110001010010001110",
40560 => "001000110001100101001110",
40561 => "001000000110011100110111",
40562 => "000100101101100101101010",
40563 => "000000001010111101001001",
40564 => "111001111010110111110001",
40565 => "110011001000111000110100",
40566 => "101111000010110001101010",
40567 => "101110101100100010101000",
40568 => "110010000010010110000000",
40569 => "110111101011011011001111",
40570 => "111100111011010101111010",
40571 => "000000101101001101010001",
40572 => "000011110101101111001001",
40573 => "000111000000010001000000",
40574 => "001000101010011100111010",
40575 => "000110110101001000110011",
40576 => "000011000100001011001100",
40577 => "111111011100000011011001",
40578 => "111100000010111000001000",
40579 => "111001111101100010100101",
40580 => "111001001000101100110010",
40581 => "110111111010010100001100",
40582 => "110101111010001110010011",
40583 => "110011100010010001100100",
40584 => "110011000011011111100100",
40585 => "110101010100001000010110",
40586 => "110110111101100110011010",
40587 => "110111001110101010011110",
40588 => "111000011000000101011101",
40589 => "111010110100111010001010",
40590 => "111101110100100101101110",
40591 => "000000101010111011000001",
40592 => "000011011001000100110111",
40593 => "000110110111111100100011",
40594 => "001011101101000111011010",
40595 => "010000101010011110101000",
40596 => "010011010011111100011000",
40597 => "010011001101001110001000",
40598 => "010001100101111101101100",
40599 => "001110100111100101101010",
40600 => "001001111000010111110110",
40601 => "000100011001110001110100",
40602 => "000000011001011100011111",
40603 => "111110101111001100011110",
40604 => "111110000101001101111000",
40605 => "111101011001000010100111",
40606 => "111100111101100010111111",
40607 => "111100100111011111100110",
40608 => "111011110000011000101111",
40609 => "111010001110010001111100",
40610 => "111000001110100010101001",
40611 => "110110111101111101000111",
40612 => "110111001111000000100011",
40613 => "111000111011011111001101",
40614 => "111100011100011110110111",
40615 => "000001000101101100101100",
40616 => "000101100110010011010001",
40617 => "001001010001100001111010",
40618 => "001011011111100000100011",
40619 => "001100010100011010101000",
40620 => "001010110000001000111101",
40621 => "000101110110111101000101",
40622 => "111110011101101100010000",
40623 => "110101001011000110111100",
40624 => "101100010000110001101000",
40625 => "100110011010110111100111",
40626 => "100011101000111011001000",
40627 => "100011101010000110111001",
40628 => "100110011001101101001010",
40629 => "101011010101110111100010",
40630 => "110001000100110011100110",
40631 => "110101111111110101010001",
40632 => "111010011101000100010001",
40633 => "111110010111000001010001",
40634 => "000000100000101010101010",
40635 => "000000111101011100000111",
40636 => "000000100101011000110110",
40637 => "000000010001101010000001",
40638 => "000000001001101001000010",
40639 => "000000001011000010110011",
40640 => "000000101101101000111111",
40641 => "000001011000011111010110",
40642 => "000010000110110000101010",
40643 => "000011010110010001100011",
40644 => "000100110001110011111001",
40645 => "000101110110111101011111",
40646 => "000110010011000100000111",
40647 => "000101111011000110110000",
40648 => "000100111100001010011010",
40649 => "000011111011000001000111",
40650 => "000011010010111010111111",
40651 => "000010111011000111011100",
40652 => "000010011111111111010110",
40653 => "000010000101101100001110",
40654 => "000001101101000000010011",
40655 => "000001000110101100100110",
40656 => "000000110101001001110011",
40657 => "000001100111000000000000",
40658 => "000011001110000101000010",
40659 => "000101001011101011000011",
40660 => "000110111010101101110100",
40661 => "001000011011111011100100",
40662 => "001010011010100111100101",
40663 => "001100000100110000001100",
40664 => "001100000101101001111100",
40665 => "001010110111101011000111",
40666 => "001001100111010111100100",
40667 => "001000100001111110100110",
40668 => "000110111101010000011100",
40669 => "000100101110000100000001",
40670 => "000001110010001101000100",
40671 => "111110001011010100101111",
40672 => "111011010010010110101101",
40673 => "111001110011010111110110",
40674 => "111000011100111000010110",
40675 => "110110100001110010010011",
40676 => "110011111111110101100000",
40677 => "110001011001001011101010",
40678 => "110000011100001001101010",
40679 => "110001100001100001001100",
40680 => "110011001001101100011000",
40681 => "110100010101010110110000",
40682 => "110101011100101010001010",
40683 => "110111010010000110110110",
40684 => "111010000010011100000000",
40685 => "111110000111001100100101",
40686 => "000011001100001100001111",
40687 => "000111010110011101000011",
40688 => "001001100110001000100111",
40689 => "001001111011000010111110",
40690 => "001001000010001000011000",
40691 => "001000000001110110000000",
40692 => "000101111011001010001111",
40693 => "000010000000101001100101",
40694 => "111110000110100001110010",
40695 => "111011110000101110010111",
40696 => "111010101111001011001111",
40697 => "111001111111011000001010",
40698 => "111001000010110011000000",
40699 => "110111011011011010110000",
40700 => "110101100110101100110110",
40701 => "110101100011001001011011",
40702 => "110111010010000001110100",
40703 => "111001010011110111000000",
40704 => "111010101110101000101110",
40705 => "111011010111100001101001",
40706 => "111100100011100110011000",
40707 => "111111000110100111110011",
40708 => "000011000000110000000000",
40709 => "001000010100110110010101",
40710 => "001101010101000011110100",
40711 => "010000110010000011001010",
40712 => "010011011101001110010100",
40713 => "010101011111110110100100",
40714 => "010110100111101001011100",
40715 => "010110101001101001101010",
40716 => "010100111111010001010110",
40717 => "010001110000011101101000",
40718 => "001110001000110111000110",
40719 => "001011011111001001001001",
40720 => "001001101110010011100101",
40721 => "000111100111101000000011",
40722 => "000110011000110100110010",
40723 => "000111000000110100110111",
40724 => "000111001000111110100110",
40725 => "000110011111010110000010",
40726 => "000110001101101100100010",
40727 => "000101101100000100101101",
40728 => "000100010110001010001011",
40729 => "000001011011111110010010",
40730 => "111110011101011010000111",
40731 => "111101110000000101101101",
40732 => "111101111011000101001100",
40733 => "111110000111000001110101",
40734 => "111111001110101000101111",
40735 => "000001001010010101101000",
40736 => "000010101000001000111010",
40737 => "000010010110001111111101",
40738 => "000001010000110100111011",
40739 => "111111111101011011000011",
40740 => "111101010110000100100110",
40741 => "111000110011001110111000",
40742 => "110010001010111111000110",
40743 => "101011010111011101110000",
40744 => "100111000010110101111001",
40745 => "100101111111010001100100",
40746 => "100111011101001000101001",
40747 => "101001011101011110001010",
40748 => "101011101101111001101010",
40749 => "101111110000010010110010",
40750 => "110101011011001111100011",
40751 => "111011000011010000111111",
40752 => "111111011110100100100111",
40753 => "000011000010100011000011",
40754 => "000110010100011010100110",
40755 => "001010000011011010110001",
40756 => "001110101110010110111000",
40757 => "010001111111100110010010",
40758 => "010001000110011110111010",
40759 => "001100111000001010110110",
40760 => "001000011001101010110000",
40761 => "000100101111001110010100",
40762 => "000000110000000011011001",
40763 => "111100110111011001101110",
40764 => "111010010010111001110110",
40765 => "111000110101101111111000",
40766 => "110111101111000111100101",
40767 => "110110110111010110110001",
40768 => "110110111010000111100001",
40769 => "110111100011101011000010",
40770 => "111000010111001001111001",
40771 => "111010000101110011110010",
40772 => "111100111000001000110110",
40773 => "000000101000101010011011",
40774 => "000101100100111100000011",
40775 => "001010100011111111010000",
40776 => "001101001000100110111100",
40777 => "001100101000001011000010",
40778 => "001011011110110111000100",
40779 => "001010111100100111111001",
40780 => "001001100100110100011110",
40781 => "000110000111111000101011",
40782 => "000000111001011100010000",
40783 => "111011011100001001101110",
40784 => "110110101111111101000111",
40785 => "110011000101111110100010",
40786 => "110000100111001001100110",
40787 => "101111001101100111110010",
40788 => "101111001101101011100100",
40789 => "110000011010000011111010",
40790 => "110010010001110111010010",
40791 => "110100101000111101100001",
40792 => "110110101010000000011001",
40793 => "110111111011011101010000",
40794 => "111000110010011001010001",
40795 => "111001110111110101001101",
40796 => "111011110100011100111010",
40797 => "111101110010110110101111",
40798 => "111110110000100110100011",
40799 => "111110110100100110110101",
40800 => "111110011111000001110000",
40801 => "111110001110101101110100",
40802 => "111101100110101010101101",
40803 => "111100000000111101001100",
40804 => "111010100101100011110100",
40805 => "111010010111010111101000",
40806 => "111010100101010111010101",
40807 => "111010111011111000100100",
40808 => "111100010001011010000001",
40809 => "111110011100100000010000",
40810 => "000000011011101000010000",
40811 => "000001111001010101101001",
40812 => "000011000110110111100100",
40813 => "000011111111110100110100",
40814 => "000100000110000001001101",
40815 => "000010110110011100010111",
40816 => "000000011101100100010100",
40817 => "111110101001101101100010",
40818 => "111110010100111110100101",
40819 => "111110110110110100001010",
40820 => "000000011100100111000011",
40821 => "000010111100001010101110",
40822 => "000101011011111111000101",
40823 => "001000000110101101000101",
40824 => "001010111111000011111110",
40825 => "001101000101101100110110",
40826 => "001101010110010000100110",
40827 => "001011101010000001011111",
40828 => "001000110000110010101000",
40829 => "000101101110111101000111",
40830 => "000011011011010000000110",
40831 => "000000111001011110001110",
40832 => "111101000100111000011011",
40833 => "111001011011100110110101",
40834 => "110111100101000110110110",
40835 => "110110111101001100100100",
40836 => "110110010111111101001000",
40837 => "110101111000011111100010",
40838 => "110110001101111101010110",
40839 => "110111101001101010000111",
40840 => "111001101000110101001111",
40841 => "111011010010000100011110",
40842 => "111100111111010110101100",
40843 => "111111100101000000100011",
40844 => "000010010011010110011110",
40845 => "000100001100101011000110",
40846 => "000101001001000111011101",
40847 => "000101011001001010111010",
40848 => "000100110110110100111110",
40849 => "000011001110010001100110",
40850 => "000001001001011100101110",
40851 => "111111011011101010100101",
40852 => "111110010000001100110110",
40853 => "111101101111111010001111",
40854 => "111101101010111011100110",
40855 => "111101100000011001000101",
40856 => "111100111010110000100110",
40857 => "111011110011001101101001",
40858 => "111010111000101101100010",
40859 => "111011001100001111011111",
40860 => "111100011101011100001110",
40861 => "111101101101000010101100",
40862 => "111110110010101101011001",
40863 => "000000110010100001101011",
40864 => "000100011110101011111000",
40865 => "001000011101101111010111",
40866 => "001011010101010101010100",
40867 => "001101100001011001011110",
40868 => "001110011100000000001000",
40869 => "001101000101111000110010",
40870 => "001010001011001110100000",
40871 => "000110011001010001111010",
40872 => "000010101000101001001010",
40873 => "111111111111001010001010",
40874 => "111110101101011101100111",
40875 => "111110111011111100001100",
40876 => "000000011000101000111011",
40877 => "000010110011110110000000",
40878 => "000110011000110000000010",
40879 => "001010100010100001111001",
40880 => "001111001110111111000010",
40881 => "010011111010111000101000",
40882 => "010110101010010010011100",
40883 => "011000000110001011111011",
40884 => "011000100011110100001011",
40885 => "010110110100001101111100",
40886 => "010100101101100001000100",
40887 => "010010010100100001010110",
40888 => "001110011110010110100100",
40889 => "001011011011100110011010",
40890 => "001001101011011100111010",
40891 => "001000110110000011010100",
40892 => "001000110110011100000100",
40893 => "001000101101110110001000",
40894 => "001000011000110001011101",
40895 => "000101111110111000011001",
40896 => "000001111111110011001001",
40897 => "111110100100111011010110",
40898 => "111001010001001011010111",
40899 => "110011001010010111011100",
40900 => "101111000001000001011010",
40901 => "101011101111001111011100",
40902 => "101010010001101100011110",
40903 => "101011110010001011010000",
40904 => "110000010111101100011110",
40905 => "110111001100011110001100",
40906 => "111101101011101100111111",
40907 => "000010111011010111001110",
40908 => "000110010000010100110010",
40909 => "000111101101100011000000",
40910 => "001000100001001100111010",
40911 => "001000010101110110110010",
40912 => "000110101111101100011110",
40913 => "000011011101011011011101",
40914 => "111111011010000110100010",
40915 => "111100011111000001111001",
40916 => "111011001001010011100011",
40917 => "111010011011101001111111",
40918 => "110111101110111001100000",
40919 => "110010100111100110010110",
40920 => "101101100100010101000100",
40921 => "101001110100111111111110",
40922 => "100111111001000001010001",
40923 => "100111010001001000100001",
40924 => "101000001001010001011010",
40925 => "101100000101010100110110",
40926 => "110010110011100101011110",
40927 => "111011101001010000100001",
40928 => "000101011111100101000100",
40929 => "001110010011011110011100",
40930 => "010100111111111101000010",
40931 => "011000110111101110000111",
40932 => "011010001001000100100001",
40933 => "011001101010110100101110",
40934 => "010111001111100010110010",
40935 => "010001110000110100111110",
40936 => "001001000011111010011100",
40937 => "111111110111001110101001",
40938 => "111000111011100001110011",
40939 => "110100010111111010011110",
40940 => "110001100010100100110110",
40941 => "110000010000100100101100",
40942 => "110000110001011010010110",
40943 => "110010100111111101010100",
40944 => "110100101110100101101110",
40945 => "110110110010000000100001",
40946 => "111000100100011010101110",
40947 => "111001101100011000000110",
40948 => "111010011111100111011010",
40949 => "111011111100001010100010",
40950 => "111110100100101001011100",
40951 => "000001111010000011001010",
40952 => "000101010001011010101101",
40953 => "000111101000110101110001",
40954 => "000111101011011101000010",
40955 => "000110000111011001110010",
40956 => "000100101011010111011110",
40957 => "000011000011100100101010",
40958 => "000000010100101010010000",
40959 => "111100101100010101000110",
40960 => "111001001000010010110010",
40961 => "110110011111110000001111",
40962 => "110100010111001110101010",
40963 => "110010011000100011101010",
40964 => "110001010110100001110110",
40965 => "110001101101011110011000",
40966 => "110011010101110001111010",
40967 => "110101101001010010111110",
40968 => "111000000110110100101010",
40969 => "111010100100011000101001",
40970 => "111100010101011110101011",
40971 => "111101000110101001100100",
40972 => "111101101000011110111110",
40973 => "111110110100110000000001",
40974 => "000000001100110110000100",
40975 => "000000001101001000111000",
40976 => "111110101000101101001110",
40977 => "111100001100110110011100",
40978 => "111001110110101111011011",
40979 => "111000010111001000100101",
40980 => "110111010010111000100100",
40981 => "110110110110011010110011",
40982 => "110111100001111011011110",
40983 => "111001000111111100011110",
40984 => "111011010010101011001010",
40985 => "111101100110000101111110",
40986 => "000000011010110101110111",
40987 => "000011000011010101100011",
40988 => "000100001001010000001110",
40989 => "000100110001000110111101",
40990 => "000101001010010010101010",
40991 => "000100010110011000001100",
40992 => "000010101101111110010011",
40993 => "000000111010101000110010",
40994 => "111111010111011101110110",
40995 => "111101100110101110001101",
40996 => "111011011100110100010000",
40997 => "111010001000111011001110",
40998 => "111001111111110001011000",
40999 => "111010110011000000110010",
41000 => "111100011011000101101011",
41001 => "111110011000011010000111",
41002 => "000000111000000010000111",
41003 => "000011101001011110001111",
41004 => "000101100110011001100010",
41005 => "000110110001011001000100",
41006 => "000111011010100110110110",
41007 => "000111010000100110000011",
41008 => "000110011010100011000001",
41009 => "000100101000000011001111",
41010 => "000010001000110010101100",
41011 => "000000100101101001001110",
41012 => "000000010101001111000000",
41013 => "000000001110111101100011",
41014 => "000000000010100001001001",
41015 => "000000010100111010110111",
41016 => "000001001111001001100110",
41017 => "000010001001110000101010",
41018 => "000010101101010011010111",
41019 => "000010111000100001111111",
41020 => "000010100011101101100111",
41021 => "000010000111001110111101",
41022 => "000001111111000010000001",
41023 => "000010001101000111110011",
41024 => "000010011110100010010010",
41025 => "000010000100100101000010",
41026 => "000001001100001001010001",
41027 => "000000110111100101111100",
41028 => "000000111000000111111011",
41029 => "000000011001110010111001",
41030 => "000000001110111000010010",
41031 => "000010000011001111010111",
41032 => "000101101001100100100000",
41033 => "001000110101010100011101",
41034 => "001010100110111000001100",
41035 => "001011100110011110101110",
41036 => "001011111111010111111010",
41037 => "001011010001101001100101",
41038 => "001000101010001011110101",
41039 => "000100011111111011100110",
41040 => "000000011001010001110111",
41041 => "111100110101001001101100",
41042 => "111010011001100101111000",
41043 => "111001100100100100000111",
41044 => "111001001101100000100111",
41045 => "111001101011110101010001",
41046 => "111011111011000000001001",
41047 => "111111010100001000001111",
41048 => "000011010100010100101101",
41049 => "000110101101111001001000",
41050 => "001000001000101000110110",
41051 => "000111111100111011001110",
41052 => "000111101111010101100110",
41053 => "000111111001100001111100",
41054 => "000110111111000010010001",
41055 => "000101000100111010000011",
41056 => "000011101000011000010000",
41057 => "000010100000111110100110",
41058 => "000000101111010110000010",
41059 => "111110000000011110100111",
41060 => "111011000101101010111000",
41061 => "111001010011001101111110",
41062 => "111001100011000001011000",
41063 => "111010000000011001100000",
41064 => "111000100011010111100101",
41065 => "110111011100110101100001",
41066 => "110111101111101001101100",
41067 => "111000000101000010111110",
41068 => "111001000011101100010110",
41069 => "111010000100000110111001",
41070 => "111011001001000101001011",
41071 => "111101111110101101101010",
41072 => "000010010010100101111111",
41073 => "000111011111111110011001",
41074 => "001100011001000010001100",
41075 => "001111101101011001110010",
41076 => "010001010101001110000000",
41077 => "010001101010001110001000",
41078 => "010010001011111001000110",
41079 => "010001111000000001101100",
41080 => "001110100001110011001100",
41081 => "001001001000110101100010",
41082 => "000011011111101100101100",
41083 => "111110110011000110110110",
41084 => "111011001001001110001000",
41085 => "111000101000011000010100",
41086 => "111000011111000001011000",
41087 => "111010111001011110111110",
41088 => "111110101001001100111000",
41089 => "000001011010101011010101",
41090 => "000010110100010101000100",
41091 => "000100110111010101011100",
41092 => "000111101100101011101110",
41093 => "001010011101111001100101",
41094 => "001100011001111001000000",
41095 => "001100101111000000000100",
41096 => "001011011011011101011010",
41097 => "001000101110001001010000",
41098 => "000101110011001010110100",
41099 => "000010110110100100010111",
41100 => "111111111111010100110111",
41101 => "111111001000100000101011",
41102 => "111111000010110011101010",
41103 => "111101110101001011011011",
41104 => "111101000011000000000011",
41105 => "111101000100011000111001",
41106 => "111101011000001011000101",
41107 => "111110010100111101101100",
41108 => "111111110110100101100101",
41109 => "000010001010110010101101",
41110 => "000100110010001110010101",
41111 => "000110101011110001011101",
41112 => "000111101111000000000111",
41113 => "000110110011100000100111",
41114 => "000010110110000010001010",
41115 => "111101011100101010100001",
41116 => "111000111000110100000100",
41117 => "110101111100101110101100",
41118 => "110100000011001100111000",
41119 => "110011011001110100001000",
41120 => "110101010010001011110011",
41121 => "111001001001111101001001",
41122 => "111101101011100001101111",
41123 => "000001101111101100110101",
41124 => "000011111010111101011111",
41125 => "000100101100111111100110",
41126 => "000100100001110100011100",
41127 => "000001111101011000010100",
41128 => "111101000010000000000111",
41129 => "110110111010011010111010",
41130 => "110001000101110100111100",
41131 => "101101111111001100100100",
41132 => "101101111000111111101100",
41133 => "101110111100000101000100",
41134 => "110000111000000001000110",
41135 => "110011110001111110010010",
41136 => "110110011010100011011110",
41137 => "111000110100100010011111",
41138 => "111011001100110011111100",
41139 => "111011110101001011110101",
41140 => "111010000101011101101011",
41141 => "110111101100100010001000",
41142 => "110110011000110101101111",
41143 => "110110010001101101101010",
41144 => "110110110011111110100110",
41145 => "110111110110011100100110",
41146 => "111001001001100011110000",
41147 => "111011000111011010001000",
41148 => "111101111000110111110101",
41149 => "000000000011100011111011",
41150 => "000001000101110110111001",
41151 => "000000111010010101101001",
41152 => "111110111110001100011111",
41153 => "111100001100100111111110",
41154 => "111001100011100101111010",
41155 => "110111010000001101001110",
41156 => "110101111010111011111111",
41157 => "110101000011101000010100",
41158 => "110011100010001010100110",
41159 => "110010010010001100101000",
41160 => "110011010001011001110100",
41161 => "110111010101010011010100",
41162 => "111101011010101001000101",
41163 => "000011000010110110001001",
41164 => "000110110011011000100111",
41165 => "001001001100000110001100",
41166 => "001011001000011111001011",
41167 => "001101000011100010000010",
41168 => "001101111010010101011000",
41169 => "001100011010110111110110",
41170 => "001001101100111000100101",
41171 => "000111111011000010110100",
41172 => "000110111110000110011001",
41173 => "000100111101001111101010",
41174 => "000001101110101101100001",
41175 => "111111001101100011101101",
41176 => "111110100001010001000011",
41177 => "111111000010110101010010",
41178 => "111111111010110111001001",
41179 => "000001001011101100011100",
41180 => "000010111110110001000110",
41181 => "000100110111011001011111",
41182 => "000110001111100010110010",
41183 => "000110110101011101011100",
41184 => "000111010000111111110101",
41185 => "000111101111011001000010",
41186 => "000111001110100111000110",
41187 => "000101100110010010000001",
41188 => "000011101111000101101101",
41189 => "000010010110001011111001",
41190 => "000001111100001101110101",
41191 => "000010100111110000110110",
41192 => "000100001001100100011100",
41193 => "000110000111011011010101",
41194 => "001000001000101110110010",
41195 => "001010000011001000101011",
41196 => "001011110001011001110000",
41197 => "001100101000100111010000",
41198 => "001011001101111010111001",
41199 => "000111100110000000100111",
41200 => "000011111111010011111100",
41201 => "000010000110001010100111",
41202 => "000001110100101001010010",
41203 => "000010000101000011111010",
41204 => "000001111111111111000101",
41205 => "000001011000001110100110",
41206 => "000000011000100100011001",
41207 => "111111001101101111110101",
41208 => "111101010101010000011101",
41209 => "111010011110111010001011",
41210 => "110111100001001111111010",
41211 => "110100010100010001100101",
41212 => "110000011000100011011010",
41213 => "101101001111010101001110",
41214 => "101100110110011110111110",
41215 => "101111000111101010001010",
41216 => "110001111101000111000100",
41217 => "110011111101010101110000",
41218 => "110101111100001011111101",
41219 => "111000000001110111000001",
41220 => "111000111110011001101110",
41221 => "111000110001110011010110",
41222 => "111000100010101011100010",
41223 => "111001000101110001100000",
41224 => "111001100001010000111011",
41225 => "111000010011000100001100",
41226 => "110110110001010110000110",
41227 => "110111010000001100011000",
41228 => "111001100101010000010111",
41229 => "111011111100010101011110",
41230 => "111101101000011000111010",
41231 => "111111011010011100010011",
41232 => "000000011011000111001100",
41233 => "000000010010101111001010",
41234 => "000000001110001110000111",
41235 => "111110111100101010101010",
41236 => "111100110000111001100110",
41237 => "111100010000000011111001",
41238 => "111101010000110101110100",
41239 => "000000000010100011100101",
41240 => "000100111111101101011011",
41241 => "001001110101010010011110",
41242 => "001101011010010101111100",
41243 => "010000110111111000110010",
41244 => "010011100100000011111010",
41245 => "010011001111011001111010",
41246 => "010000111111111111111110",
41247 => "001111011001100100111110",
41248 => "001110011111100000101010",
41249 => "001101110101001111011000",
41250 => "001100010111110011111100",
41251 => "001001110011011001010110",
41252 => "001000000111001010010001",
41253 => "000111101011010110101011",
41254 => "000111010011110000011111",
41255 => "000110110010001100010110",
41256 => "000111000000000110111111",
41257 => "001000011010011000111010",
41258 => "001001101101011111010010",
41259 => "001001111000001010111101",
41260 => "001000111100100010000000",
41261 => "001000001001000001001100",
41262 => "001000111101010101010001",
41263 => "001010001111111101111101",
41264 => "001010110010100000000000",
41265 => "001011001011011010011010",
41266 => "001011101100101011001100",
41267 => "001011111110000001010101",
41268 => "001011001011000011101011",
41269 => "001001100000010010011001",
41270 => "000111111010100110110101",
41271 => "000110001111001110111000",
41272 => "000100010010001011111011",
41273 => "000001101010011101110010",
41274 => "111100111001110100011111",
41275 => "110101100111011010101001",
41276 => "101110000011001111101100",
41277 => "101000110010000100111110",
41278 => "100110011011101010100101",
41279 => "100110111100101110101011",
41280 => "101010000101111111110100",
41281 => "101111001001110001010000",
41282 => "110101100011001111101001",
41283 => "111100010010011111100001",
41284 => "000010010110100101111111",
41285 => "000110111100001100111010",
41286 => "001001001011111001101101",
41287 => "001001011100011010110010",
41288 => "001000011011100000010110",
41289 => "000110000101101100000100",
41290 => "000010100100011010000001",
41291 => "111101111000001100010001",
41292 => "110111111111011010001111",
41293 => "110010001011111100010110",
41294 => "101110011101001010010100",
41295 => "101101010100110110110010",
41296 => "101101010001100010110100",
41297 => "101101001010101100011110",
41298 => "101101010010101010100100",
41299 => "101101100011000001100110",
41300 => "101110000011110101001010",
41301 => "101111110000010001100010",
41302 => "110010010100000010100110",
41303 => "110100111110011010110110",
41304 => "111000001011010110011000",
41305 => "111100010100110000111001",
41306 => "000001000000100100000110",
41307 => "000101001011011100110100",
41308 => "000111101010010010001000",
41309 => "001000010111100100010110",
41310 => "001000000101100100000101",
41311 => "000111001101000111000100",
41312 => "000110000101101000110110",
41313 => "000101000000100011011110",
41314 => "000010110010000000011010",
41315 => "111110110000100011010010",
41316 => "111010110010100011011110",
41317 => "111000001110010111001100",
41318 => "110110011000111100001100",
41319 => "110100110010000110110100",
41320 => "110100000110010100110010",
41321 => "110101010001010111001101",
41322 => "111000010100011000001100",
41323 => "111100100001011001011010",
41324 => "000001001100011100010100",
41325 => "000101111101010000010110",
41326 => "001010101101010101001010",
41327 => "001111000001000010000010",
41328 => "010010010010001010010110",
41329 => "010100110010110000110000",
41330 => "010110100100010100110100",
41331 => "010110001100111101010110",
41332 => "010011000011110000011010",
41333 => "001110000000011111010010",
41334 => "001000010010100110000000",
41335 => "000011100111010111001010",
41336 => "000000000011110010010010",
41337 => "111100011000110001111110",
41338 => "111001110001100011110000",
41339 => "111001100110111100011100",
41340 => "111011010111100011000100",
41341 => "111110100000000001101010",
41342 => "000010010100111111011010",
41343 => "000110011111001111101110",
41344 => "001010100110010111000001",
41345 => "001101010010010100010010",
41346 => "001110001011011110010100",
41347 => "001101110011011000001110",
41348 => "001100011001001110110000",
41349 => "001010101011010101001000",
41350 => "001001010001000101111000",
41351 => "001000000011100110111010",
41352 => "000110110100011110110000",
41353 => "000101110101101100100010",
41354 => "000101100111111001101011",
41355 => "000101011100100100000111",
41356 => "000100001001101101111010",
41357 => "000010011101110110000110",
41358 => "000010001101110011100100",
41359 => "000011110001100001100111",
41360 => "000101001110100100111010",
41361 => "000100110001011110001000",
41362 => "000011001010100100110010",
41363 => "000001101111110010001000",
41364 => "000000111001100001010011",
41365 => "000001000110100001001101",
41366 => "000001110000110010010001",
41367 => "000001111011000000001111",
41368 => "000010010001111111011011",
41369 => "000010101000011001111011",
41370 => "000010101000000000011001",
41371 => "000011110011010101111011",
41372 => "000101000010101100101010",
41373 => "000011111101110010101110",
41374 => "000001100111000010011111",
41375 => "111110011100101000111010",
41376 => "111001110111000010001100",
41377 => "110100000011100010010110",
41378 => "101100001001100000001000",
41379 => "100100010110110001110001",
41380 => "100001001110100100010101",
41381 => "100001100010000000011111",
41382 => "100010000101110001110000",
41383 => "100010110100011001101001",
41384 => "100100001001100111111001",
41385 => "100111100010001011011001",
41386 => "101101110100111000010000",
41387 => "110101001111100010101001",
41388 => "111100100001101100111001",
41389 => "000010100110000010100100",
41390 => "000101101011010111000101",
41391 => "000101101111000111010110",
41392 => "000011100100010000011010",
41393 => "111111110011101001100000",
41394 => "111011100010011110000011",
41395 => "110111100010101111100001",
41396 => "110100111111101000110010",
41397 => "110100111011010001010100",
41398 => "110110101010101100011010",
41399 => "111010000101010101101001",
41400 => "111110100111111100001111",
41401 => "000001000100110011111010",
41402 => "000000010000101111110110",
41403 => "111110001111000011001100",
41404 => "111100010011001001111100",
41405 => "111010110111110000010111",
41406 => "111001111000100010110010",
41407 => "111001100001111100111011",
41408 => "111011001000111011010110",
41409 => "111111000100110101010110",
41410 => "000100011011011001001111",
41411 => "001010100000101010111100",
41412 => "010000111111011111011010",
41413 => "010110101111100110011100",
41414 => "011001100000001001000011",
41415 => "011001000011110110100001",
41416 => "010111101111000100110000",
41417 => "010110011111001011010100",
41418 => "010100100110111110011110",
41419 => "010001010001000111001000",
41420 => "001100011101101101110000",
41421 => "001000001110100101000001",
41422 => "000110000100010111110110",
41423 => "000100011100101001010110",
41424 => "000010001000101101110001",
41425 => "000000010011100011001010",
41426 => "111111011011111100010111",
41427 => "111110011010011100000100",
41428 => "111100111011110111011000",
41429 => "111100101001101111100101",
41430 => "111111010011110011101101",
41431 => "000011100010100010011000",
41432 => "000110011011011111010101",
41433 => "000111111111110100000000",
41434 => "001010010000100000011000",
41435 => "001101100011011011000100",
41436 => "001111101100001101111110",
41437 => "001110111000110111001000",
41438 => "001100011110011010001100",
41439 => "001001110111101111011110",
41440 => "000110100100100101000000",
41441 => "000010111000111110110111",
41442 => "111111110111010001000000",
41443 => "111101110010000010000101",
41444 => "111100100001110000010111",
41445 => "111011011110110111010101",
41446 => "111010011001001011000000",
41447 => "111001100111001111111000",
41448 => "111000100101111011000001",
41449 => "110110110111111010010010",
41450 => "110101010101010110101110",
41451 => "110100010100000001110111",
41452 => "110010101110001100011110",
41453 => "101111110000010001010010",
41454 => "101100001001010110000010",
41455 => "101001011101000000001000",
41456 => "101000101011101110010010",
41457 => "101010010000010101100000",
41458 => "101110000010111000100000",
41459 => "110010101000011010000010",
41460 => "110110011111001110010101",
41461 => "111001110111010101110000",
41462 => "111101100110100010001000",
41463 => "000001010000001101011000",
41464 => "000011011111111101110100",
41465 => "000011101000101100011000",
41466 => "000010011001100111100011",
41467 => "000000110011010010101110",
41468 => "111110100100110001001000",
41469 => "111011001010100100010001",
41470 => "110111001010111011111010",
41471 => "110011101001111101001000",
41472 => "110001000000110110001100",
41473 => "101111010011001111111000",
41474 => "101111000101001100011010",
41475 => "110000101110010001101110",
41476 => "110011010100010011110000",
41477 => "110101100010101101101000",
41478 => "110111001010010001100110",
41479 => "111000111000000110000101",
41480 => "111010111110110101010101",
41481 => "111101000000101111011010",
41482 => "111110110011100001010101",
41483 => "000000111011001111110001",
41484 => "000011110110101000000100",
41485 => "000111010001111001000000",
41486 => "001010011100001110100000",
41487 => "001100110111010101010110",
41488 => "001110001110001100001110",
41489 => "001110001100100110110110",
41490 => "001101010010010111111100",
41491 => "001100011100111011000010",
41492 => "001011001000100001001111",
41493 => "000111101000011010000100",
41494 => "000010011010010110000100",
41495 => "111110001010000001011101",
41496 => "111011111011101000100000",
41497 => "111010011111100110000001",
41498 => "111001010010011110100000",
41499 => "111001011001001100001001",
41500 => "111011101000110001110110",
41501 => "111111010000111001111001",
41502 => "000010101110011010110100",
41503 => "000101101011100101011101",
41504 => "001001001111000110001011",
41505 => "001101001111011011101100",
41506 => "001111101001100111101000",
41507 => "010000000111100011101000",
41508 => "010000011110001010100100",
41509 => "010000100100000101000000",
41510 => "001110010101001010100010",
41511 => "001001101101000100101100",
41512 => "000100100101011001111110",
41513 => "000000001111000001101110",
41514 => "111100100001111100010111",
41515 => "111000111110111110111101",
41516 => "110110011000101001010111",
41517 => "110110001110111100001000",
41518 => "111000101000010010001101",
41519 => "111100111011100001100110",
41520 => "000010110000111100011101",
41521 => "001000111001011001000001",
41522 => "001101101001010111111000",
41523 => "010000011101101110001010",
41524 => "010001111011010101100000",
41525 => "010010101111001111111100",
41526 => "010010100001010010011010",
41527 => "010000010000000011110100",
41528 => "001100000111001111001100",
41529 => "000111101001111011111100",
41530 => "000100011110000000111101",
41531 => "000010101010001001011000",
41532 => "000000111000001000011110",
41533 => "111111000010101010110100",
41534 => "111110101111010100101001",
41535 => "000000001011001111001011",
41536 => "000001101001010100010000",
41537 => "000001111111110101000100",
41538 => "000010000110101011111010",
41539 => "000010110110000101011000",
41540 => "000010010000001110001100",
41541 => "111110011100011111100011",
41542 => "111001110010011110000111",
41543 => "110111011001000011110101",
41544 => "110110011010100000110000",
41545 => "110100001101000001001001",
41546 => "110000101100010001000010",
41547 => "101110011101011110111000",
41548 => "101110101101010111011100",
41549 => "110000000011010001010110",
41550 => "110001100001110000110010",
41551 => "110011010110100111111100",
41552 => "110101110101001001011100",
41553 => "111000110001111101101100",
41554 => "111011000110000000001101",
41555 => "111100110101100001110111",
41556 => "111111011110010101000011",
41557 => "000010001010010110110101",
41558 => "000011001010110100110110",
41559 => "000011001101000110110101",
41560 => "000011010001111010010011",
41561 => "000011001011000101000011",
41562 => "000010000010001000101100",
41563 => "111111000111100100001001",
41564 => "111011100101001110011010",
41565 => "111001010101111100011011",
41566 => "111000101010100101001111",
41567 => "111001001010001001111010",
41568 => "111010110100111011100111",
41569 => "111101100010100100000000",
41570 => "000000000100011011111101",
41571 => "000000110110111101100001",
41572 => "000000111100001101001010",
41573 => "000001111000010110110000",
41574 => "000010010000001010101010",
41575 => "000001001100111111100101",
41576 => "000000001010111011101110",
41577 => "000000010010011100101100",
41578 => "000010011101000010111001",
41579 => "000101111111100001110011",
41580 => "001000110010010100010001",
41581 => "001011001110011110000000",
41582 => "001101110011010001111000",
41583 => "001110001000000111001010",
41584 => "001011001010000010000010",
41585 => "000110101100101101010101",
41586 => "000010110111011011011010",
41587 => "000000000110001110010101",
41588 => "111100101010110110110001",
41589 => "111000011110111010100110",
41590 => "110110010110110110011110",
41591 => "110111010000101101101110",
41592 => "111001111011000101000010",
41593 => "111101101110101010001110",
41594 => "000010000011010101001100",
41595 => "000101110100000011001000",
41596 => "001000001100100100000101",
41597 => "001000110111100110101100",
41598 => "001000010100111100001010",
41599 => "000111001001110001010100",
41600 => "000101011111000000110011",
41601 => "000011101110101110011000",
41602 => "000010101100110001011100",
41603 => "000011010011001001111000",
41604 => "000101011101100000110011",
41605 => "000111011100100001100111",
41606 => "000111101110110100010000",
41607 => "000110101100110001010000",
41608 => "000101111100101000100101",
41609 => "000110010101100110110011",
41610 => "000110100001011111011101",
41611 => "000100111100111111111011",
41612 => "000010010000011001010001",
41613 => "111111010110111010101111",
41614 => "111100011100100110110111",
41615 => "111010101101100100010011",
41616 => "111011000110100000010001",
41617 => "111100010001000100010100",
41618 => "111100101111001000101000",
41619 => "111101000110110100111100",
41620 => "111110000010010100101011",
41621 => "111110100100111010111110",
41622 => "111110000110111100000001",
41623 => "111101010111000110001001",
41624 => "111100111101001011100110",
41625 => "111101001000011000011011",
41626 => "111110000001011100101010",
41627 => "111111001111000101001101",
41628 => "000000010100011100110110",
41629 => "000001000001011011001011",
41630 => "000000100100110111011111",
41631 => "111101111001101100011011",
41632 => "111000110110001110111010",
41633 => "110010111111001001010110",
41634 => "101110001101111100111100",
41635 => "101010100011000011110010",
41636 => "100111000101011010100111",
41637 => "100100010010110001010111",
41638 => "100011011111100010001001",
41639 => "100101101101111100110001",
41640 => "101011001111110001000110",
41641 => "110010110001101110111100",
41642 => "111010001110010100000111",
41643 => "000000110100000010100111",
41644 => "000110111011000010010010",
41645 => "001100001101100110100010",
41646 => "001111011000010101110010",
41647 => "001111100111110000000010",
41648 => "001101010100010110111010",
41649 => "001001000100010000100110",
41650 => "000011001101000110101011",
41651 => "111101000011011000010100",
41652 => "111000100010101110000011",
41653 => "110101100100010010100100",
41654 => "110010101110100101001010",
41655 => "110000101011010001101110",
41656 => "110000111011001001101010",
41657 => "110011000101011100111110",
41658 => "110110001111110101000110",
41659 => "111010000010010001001101",
41660 => "111101011101001101011110",
41661 => "111111110000101101001000",
41662 => "000001111000010011010000",
41663 => "000101000111100100000100",
41664 => "001001001011100100011001",
41665 => "001100100111000001010010",
41666 => "001110101011101111001100",
41667 => "001111100000010111000100",
41668 => "001111000101111000000000",
41669 => "001101111111011110011000",
41670 => "001101001011101010001000",
41671 => "001100001111100100110000",
41672 => "001001110000111000101100",
41673 => "000101111111011010110101",
41674 => "000010101111111001100101",
41675 => "000000011000011000110100",
41676 => "111101101001001111101100",
41677 => "111010111001111101001111",
41678 => "111010001000111100101001",
41679 => "111100000100110110100010",
41680 => "111111101111010100111011",
41681 => "000011110000100100011100",
41682 => "000111011100001101111010",
41683 => "001010110101010010001101",
41684 => "001101101010000010101010",
41685 => "001111101110010000111110",
41686 => "010001100011110101100100",
41687 => "010010110110001001001000",
41688 => "010010011011000000010000",
41689 => "001111111000000110101010",
41690 => "001011011010100100011100",
41691 => "000110000000111110110011",
41692 => "000001001101000111110010",
41693 => "111101001010001110111100",
41694 => "111001001010000101011100",
41695 => "110101101101000101101010",
41696 => "110100001011101110000010",
41697 => "110101000110100100100010",
41698 => "110111101010111101000110",
41699 => "111010111101011111111000",
41700 => "111110001110011100010110",
41701 => "000000000011010111011101",
41702 => "111111110110011110010111",
41703 => "111111010100100111101111",
41704 => "111111110001000111100111",
41705 => "000000001101010111111111",
41706 => "111111101101011011001000",
41707 => "111110110010011111101101",
41708 => "111101111010010101001110",
41709 => "111101000011101111101101",
41710 => "111101001011100000001011",
41711 => "111111011010010111111011",
41712 => "000010110000110110101111",
41713 => "000101001010110101000010",
41714 => "000101101100111000001011",
41715 => "000100010101010011111011",
41716 => "000001100000000101000001",
41717 => "111101101111111000011010",
41718 => "111001010100110100011000",
41719 => "110101000100010110101001",
41720 => "110001111011000010100100",
41721 => "101111110010110000110000",
41722 => "101110101001001110101100",
41723 => "101110101001010000100000",
41724 => "101111100001110011000010",
41725 => "110001110000110001101100",
41726 => "110101110111000101101100",
41727 => "111010110011000101100101",
41728 => "111111110101111101001001",
41729 => "000101011100011001001111",
41730 => "001010110011101011101100",
41731 => "001101110100011110111000",
41732 => "001101110001111110000000",
41733 => "001011100001111011110101",
41734 => "000111100000100111111011",
41735 => "000010100100000010111000",
41736 => "111110111000110111010100",
41737 => "111101010110000011100100",
41738 => "111100101000101010000101",
41739 => "111011110111101001011101",
41740 => "111010110010011000110011",
41741 => "111001011010111100111011",
41742 => "111000100110001000100101",
41743 => "111000000100011011110011",
41744 => "110110101110011101101111",
41745 => "110101010011111101101000",
41746 => "110100111100011101100110",
41747 => "110101011001010001111110",
41748 => "110110101000101010000111",
41749 => "111000011110001100001010",
41750 => "111010101110011100010101",
41751 => "111110111100110001001011",
41752 => "000101011100001100011110",
41753 => "001011000001101101000000",
41754 => "001101011011011100101110",
41755 => "001101100000011111000100",
41756 => "001100010000100011100010",
41757 => "001001011110001010110110",
41758 => "000101000010110000101001",
41759 => "111111111010101110111010",
41760 => "111011110001011110000100",
41761 => "111001100110100011111100",
41762 => "111000111001011001110111",
41763 => "111000111001100100100010",
41764 => "111001111001001100101000",
41765 => "111100010011100011110011",
41766 => "111111100101001010111110",
41767 => "000010101001100000110100",
41768 => "000100011100110101011000",
41769 => "000100111001001100101011",
41770 => "000101100111001001101101",
41771 => "000111011000010000101011",
41772 => "001000100100101001011110",
41773 => "001000100110010011111011",
41774 => "001001001100010110011010",
41775 => "001011101000000010100100",
41776 => "001111010100001011001110",
41777 => "010010010011000101000110",
41778 => "010011010001110010000100",
41779 => "010011000101110010111010",
41780 => "010010000101011010111100",
41781 => "001111001010100101011010",
41782 => "001010101001101000000101",
41783 => "000101111111010110100100",
41784 => "000001111111100000001110",
41785 => "111111010011010000010010",
41786 => "111110001011100001000111",
41787 => "111110010010100011010110",
41788 => "111111011100100110010011",
41789 => "000001011100010100110011",
41790 => "000011110100100100010000",
41791 => "000101110111010000110000",
41792 => "000110110000101001111001",
41793 => "000110100000001111010110",
41794 => "000101100001100000111001",
41795 => "000011110110001010011011",
41796 => "000001110000101001010010",
41797 => "000000001110000001000000",
41798 => "000000001010011101100000",
41799 => "000001010000111010000001",
41800 => "000001111010001100100100",
41801 => "000001101111010000101110",
41802 => "000001111010000101010111",
41803 => "000010011101000010011001",
41804 => "000010100100110001111100",
41805 => "000001110000101001011100",
41806 => "111111011011001100001110",
41807 => "111100000010111111110111",
41808 => "111001000100111111000000",
41809 => "110111000100001100001110",
41810 => "110101111011111101001011",
41811 => "110100101101001001001010",
41812 => "110001001100100111110000",
41813 => "101011110101000111010010",
41814 => "101000010111110111111000",
41815 => "101000101000011001100110",
41816 => "101010111101101100100010",
41817 => "101101100011010111001010",
41818 => "101111011111110110111000",
41819 => "110001010111110111010100",
41820 => "110101010111100100010000",
41821 => "111011101010001011100000",
41822 => "000001100110100001000101",
41823 => "000110001001000100000111",
41824 => "001001110001011010000100",
41825 => "001011110100010011000010",
41826 => "001100001110010000001010",
41827 => "001011101001110100010101",
41828 => "001001000111100101011000",
41829 => "000011111111101111100001",
41830 => "111101110100010010010100",
41831 => "111000011011011110011110",
41832 => "110101000110011100010111",
41833 => "110011101100111010001110",
41834 => "110010101010110001001010",
41835 => "110010001000100100010000",
41836 => "110011111111100100000010",
41837 => "111000001101001011000101",
41838 => "111101011110110110110100",
41839 => "000011110000010100100110",
41840 => "001010001000111111000010",
41841 => "001110010010100111111110",
41842 => "010000001000100111101010",
41843 => "010001111011111110110110",
41844 => "010100011101000101110000",
41845 => "010110010011011111101010",
41846 => "010101110010111010001000",
41847 => "010010101100100011110010",
41848 => "001111001011100001011100",
41849 => "001100111001111100111010",
41850 => "001010010101101001111011",
41851 => "000101110011111010100101",
41852 => "000000010001100110111010",
41853 => "111011110010110101101110",
41854 => "111001010111111001101000",
41855 => "110111111011011001110110",
41856 => "110110001001000111111111",
41857 => "110100111001001001010011",
41858 => "110101001010011001111011",
41859 => "110110001111010100101011",
41860 => "110111111110111010111111",
41861 => "111010111110011111001101",
41862 => "111110001101101111100110",
41863 => "000000000110100000001001",
41864 => "000001010110001000111001",
41865 => "000011111100001110000111",
41866 => "000111001111110011111010",
41867 => "001000100101100000000000",
41868 => "000111100100000101011110",
41869 => "000101101111011000001110",
41870 => "000011001110000100010110",
41871 => "111111001010010101110111",
41872 => "111010011000001001101100",
41873 => "110110110011001111011001",
41874 => "110100100000111011001110",
41875 => "110010001010000111100000",
41876 => "110000101001101010000000",
41877 => "110010010010101110010100",
41878 => "110111000000111101001111",
41879 => "111101010101100110010110",
41880 => "000011111101001101011011",
41881 => "001001010100010101110010",
41882 => "001100111100100001110010",
41883 => "001111000000001101000100",
41884 => "001101111001110010110110",
41885 => "001000011001110010111010",
41886 => "000000011001010110110000",
41887 => "111000100111101001101110",
41888 => "110010000101111100111110",
41889 => "101101000110000010011000",
41890 => "101010011101100110111010",
41891 => "101010110111100010010100",
41892 => "101101110100010110011100",
41893 => "110010011011001011101010",
41894 => "111000011101110000110100",
41895 => "111111011100111101111100",
41896 => "000101010101011100000100",
41897 => "001000010001001010001111",
41898 => "001001010011101111000111",
41899 => "001010010110001010010101",
41900 => "001010010101110001011111",
41901 => "000111011001010100100001",
41902 => "000010011011000100010010",
41903 => "111101001101110010100101",
41904 => "111000001001000101110010",
41905 => "110011111101001001000010",
41906 => "110010010100110111110010",
41907 => "110011101101001100001010",
41908 => "110110111000100101111100",
41909 => "111001111010010010110011",
41910 => "111011001000110110001100",
41911 => "111011001000110101010111",
41912 => "111011110011010000101110",
41913 => "111100011110111011111110",
41914 => "111011001000111000100000",
41915 => "111000100000011001110010",
41916 => "110110101010010111010101",
41917 => "110110001000111111100000",
41918 => "110110110000110011100100",
41919 => "111000001000100111000111",
41920 => "111001111110010100101010",
41921 => "111100110110000010001110",
41922 => "000000100010001110011100",
41923 => "000011110101000010111001",
41924 => "000110101001100010010010",
41925 => "001001000010101110110011",
41926 => "001001110000001011011000",
41927 => "001000000101100111111001",
41928 => "000100011100000111100110",
41929 => "111111010000100111001111",
41930 => "111001110100011111101100",
41931 => "110101111011111001010111",
41932 => "110100000001100100000010",
41933 => "110011011110101000010100",
41934 => "110100010001011011110100",
41935 => "110110101100111101111101",
41936 => "111010100100000100101000",
41937 => "111110111101000010111000",
41938 => "000010100101010011110010",
41939 => "000101001001001000100000",
41940 => "000111101001111000101001",
41941 => "001010010111000011101100",
41942 => "001100001101010010001100",
41943 => "001100111001111011101010",
41944 => "001101001001010001110110",
41945 => "001101001011000001110100",
41946 => "001100110000000111001100",
41947 => "001011110111010111010001",
41948 => "001010110110000101011111",
41949 => "001001110111100100110110",
41950 => "001000100000110100100011",
41951 => "000110100010101001001101",
41952 => "000100101001010001000000",
41953 => "000011011011001000101101",
41954 => "000010101000101010100010",
41955 => "000010001001001010111110",
41956 => "000010000101111101010001",
41957 => "000010000000001000110111",
41958 => "000001100101000011001000",
41959 => "000001100010010001110100",
41960 => "000001110001011010100011",
41961 => "000001000000011000001101",
41962 => "111111010100110000110010",
41963 => "111110001101001110111100",
41964 => "111110001101011110001011",
41965 => "111110111010111010000111",
41966 => "000000000011011100111110",
41967 => "000001101000111011000110",
41968 => "000011110001111011100100",
41969 => "000110001010000011001001",
41970 => "001000000110000100100001",
41971 => "001001000100101010110011",
41972 => "001000101001101001011101",
41973 => "000110111000000111110111",
41974 => "000100010010100111010100",
41975 => "000000101001001011010010",
41976 => "111011101010011011101111",
41977 => "110110101111111111111011",
41978 => "110011101001001000111110",
41979 => "110010110110000011100100",
41980 => "110011111101001011111000",
41981 => "110110000001110011100100",
41982 => "111000011011001011110101",
41983 => "111011011000111111010110",
41984 => "111110110010111001101001",
41985 => "000001110110111110110010",
41986 => "000100001000101110110100",
41987 => "000101010011000100011000",
41988 => "000101010110011000011001",
41989 => "000101010001100010011000",
41990 => "000101010110011100001010",
41991 => "000011111111101010000110",
41992 => "000000000110111010001001",
41993 => "111011000101100000110111",
41994 => "110111011001110011001110",
41995 => "110110011110110101111010",
41996 => "111000010101101101110001",
41997 => "111011110110111101111111",
41998 => "111111011001001010100011",
41999 => "000010100000110101001111",
42000 => "000110001100000010101000",
42001 => "001010101000101101101001",
42002 => "001111000011100111101010",
42003 => "010010110101110100011010",
42004 => "010101011010110110011100",
42005 => "010110100010000111001000",
42006 => "010110101000000110011110",
42007 => "010101110001001000010110",
42008 => "010011110000001010101010",
42009 => "010001000100010010001010",
42010 => "001101111010100001101010",
42011 => "001001110011110010001010",
42012 => "000101001100110010001000",
42013 => "000001110001011000111100",
42014 => "000000011011111111111011",
42015 => "000000000010010011111110",
42016 => "111111000010111111110111",
42017 => "111101111111100000000100",
42018 => "111110100001000111000100",
42019 => "000000100001000100110000",
42020 => "000001101010111010100000",
42021 => "000000011110010001111001",
42022 => "111110101000111110111101",
42023 => "111110000111010100110100",
42024 => "111101111100101010001001",
42025 => "111101010110011101100011",
42026 => "111101101100000001000100",
42027 => "111111100001101110101101",
42028 => "000001100111111100110011",
42029 => "000011000000100001011011",
42030 => "000100010010001001011110",
42031 => "000101111110011011011110",
42032 => "000110010111110100100010",
42033 => "000100001110010101111000",
42034 => "000001011100001110100110",
42035 => "111111011100010100000100",
42036 => "111100111010101111111101",
42037 => "111001000111000000110010",
42038 => "110101011010101000110110",
42039 => "110011100010101111011110",
42040 => "110011110010010011000100",
42041 => "110101010001001010001010",
42042 => "110111110111110001010010",
42043 => "111100010111000110010000",
42044 => "000001111001100000110111",
42045 => "000101111110111111110100",
42046 => "000111011100100110110001",
42047 => "000111010100100011001111",
42048 => "000110101000110010000011",
42049 => "000101011000010001101100",
42050 => "000011101101001111011010",
42051 => "000010000101011110011000",
42052 => "000000110010010110100101",
42053 => "111111101010010010010011",
42054 => "111100110101100010010001",
42055 => "110111011000010001010110",
42056 => "110010101111100100101110",
42057 => "110001000001101100010110",
42058 => "101111111010110100001000",
42059 => "101111011010001001100100",
42060 => "110001100011001111110010",
42061 => "110101001010101110010010",
42062 => "110111110100001010110111",
42063 => "111000101111000110010011",
42064 => "111001001101011010001010",
42065 => "111011011110101000110111",
42066 => "111111001000001000001001",
42067 => "000001101100110100011010",
42068 => "000010110110010011100101",
42069 => "000010111111100110000111",
42070 => "000001011001011000111111",
42071 => "111110101100101111000101",
42072 => "111101000110011010111101",
42073 => "111101000101000101000100",
42074 => "111101000101101110110011",
42075 => "111100101111001111010110",
42076 => "111100111010001011011110",
42077 => "111100111000011100101011",
42078 => "111011101111000111011011",
42079 => "111010000101001111101111",
42080 => "110111100101101110001111",
42081 => "110100001011101010000010",
42082 => "110001110000011000110000",
42083 => "110000100010001010010100",
42084 => "101111011100011000000110",
42085 => "101111010011000001101100",
42086 => "110000110110000101100100",
42087 => "110011110011101101000000",
42088 => "111000000101111001111000",
42089 => "111101001101101000011010",
42090 => "000010111100100001110101",
42091 => "001001000111000011101110",
42092 => "001101011011011101101010",
42093 => "001101101010001000001000",
42094 => "001010100110011001001010",
42095 => "000110011011101010110001",
42096 => "000010100110010010110011",
42097 => "111111001101010111011000",
42098 => "111011010010010000010011",
42099 => "110110110011100011110101",
42100 => "110011101110110111100100",
42101 => "110011010110110000110110",
42102 => "110011111011000000100010",
42103 => "110011101110010000011100",
42104 => "110100011011100100111000",
42105 => "110111100010101000101100",
42106 => "111011100011110010011010",
42107 => "111110101000110100001000",
42108 => "000000000011101011110101",
42109 => "000000011100011101101001",
42110 => "000001000101000010011001",
42111 => "000001110111110110110011",
42112 => "000010101010010000010110",
42113 => "000100100000010000000111",
42114 => "000111100000001000100100",
42115 => "001010011001000001110110",
42116 => "001100000011010100001100",
42117 => "001011111100111000000110",
42118 => "001010100010011101111000",
42119 => "001000111001010001010110",
42120 => "000110111011110110011010",
42121 => "000011010010111111101011",
42122 => "111101111000000000101111",
42123 => "111000101011101011011010",
42124 => "110101010111010101111101",
42125 => "110011110001100110000000",
42126 => "110011011111010000111110",
42127 => "110100100101010001010010",
42128 => "110110110010010100110000",
42129 => "111001100001100010111110",
42130 => "111100010101111011010111",
42131 => "111111001010001010010110",
42132 => "000010000010101110010110",
42133 => "000100001100010000001000",
42134 => "000101001011000000111111",
42135 => "000101111110011101010100",
42136 => "000110101100010110101110",
42137 => "000110101101001000000011",
42138 => "000110011111101000100111",
42139 => "000110011010010010000000",
42140 => "000101111100100001000011",
42141 => "000100101000100101100000",
42142 => "000010110001000000110111",
42143 => "000000110001101001011000",
42144 => "111110001001011010101101",
42145 => "111010111001011100001011",
42146 => "111000011010010101110111",
42147 => "110111011001100110000001",
42148 => "110111010111011111101110",
42149 => "111000010001000010001110",
42150 => "111011001100000001001011",
42151 => "000000000010100010110011",
42152 => "000100011000001001011101",
42153 => "000110111000110011011010",
42154 => "001000101010000101001010",
42155 => "001010010000000101001100",
42156 => "001010111001110110110110",
42157 => "001010010011010110101010",
42158 => "001001100111010101000001",
42159 => "001010000000000001011100",
42160 => "001010110110111110100010",
42161 => "001011001111110110000010",
42162 => "001011100110111101001110",
42163 => "001100011100101100010010",
42164 => "001101000000111011001110",
42165 => "001100101101010111111000",
42166 => "001100001101011101011110",
42167 => "001011111111111111111111",
42168 => "001011011100110001000101",
42169 => "001010100010001011000111",
42170 => "001010011011011111011100",
42171 => "001010110110101001101110",
42172 => "001001100100110100011110",
42173 => "000101101101100101110110",
42174 => "000000101111110010100000",
42175 => "111101000010001100111010",
42176 => "111100000011110010000000",
42177 => "111100110011110000100110",
42178 => "111101011110110100101010",
42179 => "111110000001111100001101",
42180 => "111111011011100101001110",
42181 => "000001111100110000111011",
42182 => "000100010010000100001001",
42183 => "000101001001001111111000",
42184 => "000100111100110101110110",
42185 => "000100001101010010110100",
42186 => "000011000010011010111011",
42187 => "000010000011001010111010",
42188 => "000001001101010110101011",
42189 => "111111010111001011010110",
42190 => "111011011011110110011010",
42191 => "110110001110111011001011",
42192 => "110010100010110100110110",
42193 => "110001101010101111000100",
42194 => "110010010110010111001010",
42195 => "110011110110111110000110",
42196 => "110110000001001100110100",
42197 => "110111100111100111100010",
42198 => "111000001110011110000101",
42199 => "111001000111110100011101",
42200 => "111011000010101101101011",
42201 => "111101001000011111010010",
42202 => "111110110000010100011101",
42203 => "000000101111111110010011",
42204 => "000011100111001110001110",
42205 => "000110000001101000111010",
42206 => "000110100101000101010110",
42207 => "000101011101001110111010",
42208 => "000100000010010011111101",
42209 => "000011001000011000001010",
42210 => "000010011101100100111101",
42211 => "000010001111000101010110",
42212 => "000010100000010110000110",
42213 => "000010001010001111010111",
42214 => "000000111001011001101000",
42215 => "111111100010110011010110",
42216 => "111110110010000110111000",
42217 => "111110101111110101101010",
42218 => "111110110100011111001111",
42219 => "111110111101100000101011",
42220 => "000000011001110101011110",
42221 => "000011111000001111100101",
42222 => "001000100000001011110100",
42223 => "001100100101111000111100",
42224 => "001111001110110101011100",
42225 => "010000001010010000111000",
42226 => "001111000001110010011100",
42227 => "001100100001110010100100",
42228 => "001001100000100001001000",
42229 => "000101000001111010011001",
42230 => "111110001101111111111101",
42231 => "110101110011010000000000",
42232 => "101101111110000011110010",
42233 => "101001111110100001010010",
42234 => "101010011101011010010010",
42235 => "101100110101000100001110",
42236 => "110000010011110110101110",
42237 => "110101110100110110010100",
42238 => "111100110110100110100011",
42239 => "000011111011100001101101",
42240 => "001001101001001101010110",
42241 => "001101110011011111110110",
42242 => "010000011111011001101010",
42243 => "010000011101101000001100",
42244 => "001101101100011000110010",
42245 => "001001110001010100111101",
42246 => "000110010100010010110001",
42247 => "000011111100000010111100",
42248 => "000001000110001101001101",
42249 => "111101110011010010110111",
42250 => "111011010101010000011001",
42251 => "111000001101011110010110",
42252 => "110100111001111111010110",
42253 => "110011101010110001001100",
42254 => "110011000100100011010000",
42255 => "110010000011010001100110",
42256 => "110001110111110000111010",
42257 => "110011010010010000001100",
42258 => "110110111110101010111100",
42259 => "111100101001001000101100",
42260 => "000010010010011100100100",
42261 => "000110101010110110101110",
42262 => "001010010000110111000010",
42263 => "001101000001011101100000",
42264 => "001101010011000010001110",
42265 => "001010101101010011101000",
42266 => "000110110101100011100000",
42267 => "000010101110110111001111",
42268 => "111110010010001011011101",
42269 => "111000110000010010011100",
42270 => "110010100010111110111010",
42271 => "101110100000111010100110",
42272 => "101110100000010011010010",
42273 => "110000010010101000011110",
42274 => "110001100100111100110110",
42275 => "110011011000001110110110",
42276 => "110110000011101111000110",
42277 => "111000010111011110011100",
42278 => "111010011111111110011100",
42279 => "111100100000001011001110",
42280 => "111110001011111010110011",
42281 => "000000001110101101100110",
42282 => "000001110010001001010101",
42283 => "000001111110110110111000",
42284 => "000001110011000100001101",
42285 => "000001110101001000001001",
42286 => "000010001101100010001010",
42287 => "000010101000011001100011",
42288 => "000010000100100101011011",
42289 => "000000101100110010111001",
42290 => "111110111001000001001100",
42291 => "111011001111011000111101",
42292 => "110101100010101000100000",
42293 => "110000110010011100111100",
42294 => "101111001011010010000000",
42295 => "110000000110101110010000",
42296 => "110010111101010100111110",
42297 => "110111010001000101110100",
42298 => "111011010110011111110001",
42299 => "111110001011110111111010",
42300 => "000000011111010011000000",
42301 => "000010101011101101100010",
42302 => "000100001111101100101011",
42303 => "000100101100110001010111",
42304 => "000011011101010110000111",
42305 => "000000110010110010011100",
42306 => "111110010000000001001110",
42307 => "111100010001110110001010",
42308 => "111010110101110101000000",
42309 => "111010111110100101101100",
42310 => "111100101010111001110101",
42311 => "111110111010000101100000",
42312 => "000001101000110010011100",
42313 => "000100011110010010010110",
42314 => "000101110110001011011000",
42315 => "000100111010100001000001",
42316 => "000010011101101100101110",
42317 => "111111111101010010011001",
42318 => "111110100111000001000100",
42319 => "111110101110101111111101",
42320 => "111111111000101000111101",
42321 => "000001110001111111110010",
42322 => "000100001110100111110100",
42323 => "000110111001111101111000",
42324 => "001001101011010000111111",
42325 => "001100100010011100001000",
42326 => "001111000101000101011110",
42327 => "010000011110011011111000",
42328 => "010000101101000111110010",
42329 => "010000100010101110110000",
42330 => "010000011011010001111010",
42331 => "010000011111111100101100",
42332 => "010000010001100101111010",
42333 => "001110110100110011000000",
42334 => "001100001101100111110100",
42335 => "001001011011010011001001",
42336 => "000111010010011101101100",
42337 => "000101100100000100001100",
42338 => "000011100000001011001010",
42339 => "000001010011001001101000",
42340 => "111111110110001010000011",
42341 => "111111101000011111010111",
42342 => "000000000101010110110000",
42343 => "000000100110111100000011",
42344 => "000001101010111101110011",
42345 => "000010111000111011110000",
42346 => "000010111110010010011010",
42347 => "000010001000000000001100",
42348 => "000001101101001100010000",
42349 => "000010011000001100110111",
42350 => "000011010001000101111101",
42351 => "000011000110011111100101",
42352 => "000001101011110111101011",
42353 => "111111010001010111100010",
42354 => "111011101001001001111100",
42355 => "110110111101101111101000",
42356 => "110011000110111010101100",
42357 => "110001101111000000000010",
42358 => "110010000100101001001110",
42359 => "110010110100000100011100",
42360 => "110011010010101101000100",
42361 => "110011101010100101100000",
42362 => "110101000100100011001101",
42363 => "110111111100110110111110",
42364 => "111100001100100011011010",
42365 => "000001010000110001100110",
42366 => "000101100111100111111011",
42367 => "001000010100110110111101",
42368 => "001001010011110010110010",
42369 => "001000110111111001001111",
42370 => "000110111011000011010011",
42371 => "000011010000010011101110",
42372 => "111111011000001011100101",
42373 => "111100100100000111010111",
42374 => "111011001111011011100110",
42375 => "111011101000001110011010",
42376 => "111100000011000011001000",
42377 => "111011110000001111111001",
42378 => "111011101000100110001000",
42379 => "111011110101101001111001",
42380 => "111101001000001001100101",
42381 => "111111000100100111111111",
42382 => "000000010111111000010000",
42383 => "000001111011011110110001",
42384 => "000100000100100110101110",
42385 => "000110000000001000111100",
42386 => "000111011001001000000111",
42387 => "001000100010101001100101",
42388 => "001010100111111111110001",
42389 => "001101000100101100101110",
42390 => "001110011001000010011100",
42391 => "001110110001001101111100",
42392 => "001110000011001000000010",
42393 => "001100001111100000011010",
42394 => "001001110101000010101111",
42395 => "000101101101000011000001",
42396 => "111111110000011001011110",
42397 => "111010000100101010010011",
42398 => "110101101001101011101011",
42399 => "110001111101000000001100",
42400 => "101110111101011110100100",
42401 => "101101010110001100000100",
42402 => "101101010110100100011010",
42403 => "101111000001011110000000",
42404 => "110010111110100001001010",
42405 => "111001001101000100101110",
42406 => "000000011111101111111110",
42407 => "001000000101010101110000",
42408 => "001111000110011101100110",
42409 => "010011101100011000001000",
42410 => "010100110011111110101000",
42411 => "010010001111110010001010",
42412 => "001100011010110101100100",
42413 => "000101001010001111000001",
42414 => "111101101111011110101111",
42415 => "110110010101111100110100",
42416 => "101111100100100111010000",
42417 => "101010101101000000010000",
42418 => "101001010011101111011000",
42419 => "101011100100110111000010",
42420 => "110000001111101100100100",
42421 => "110101110101110110011011",
42422 => "111010111010101011001110",
42423 => "111111101101100110100100",
42424 => "000100000010001000001100",
42425 => "000100111111111110111100",
42426 => "000010001111010110011001",
42427 => "111110011110001000010011",
42428 => "111011000011001010000000",
42429 => "111000011101010100011011",
42430 => "110110111011111111011010",
42431 => "110110110110111100000000",
42432 => "111001011111110100111110",
42433 => "111110010100001010001010",
42434 => "000010110010100010000010",
42435 => "000101101100100101001010",
42436 => "000111001100100111000010",
42437 => "000111101101111101100100",
42438 => "000111001100001001010100",
42439 => "000100101001001000010000",
42440 => "000000010001001111000000",
42441 => "111011101011111100010010",
42442 => "110111111101010000111000",
42443 => "110101011001000001001001",
42444 => "110011011110101110000110",
42445 => "110010000100111101010010",
42446 => "110001110110101010100100",
42447 => "110010011010011011000110",
42448 => "110011111011000111000110",
42449 => "110111001000110100011101",
42450 => "111011000100001011111000",
42451 => "111111010101100110010001",
42452 => "000011111001101100001001",
42453 => "000111001111010100010110",
42454 => "001000110000101101110011",
42455 => "001001001111100111100000",
42456 => "001010000000110011000110",
42457 => "001011100000011101011100",
42458 => "001100001011110100101000",
42459 => "001011001001011011001001",
42460 => "001000100110011100000111",
42461 => "000100110010011101001110",
42462 => "000000101001011000001010",
42463 => "111100110001110010100101",
42464 => "111001011000001001111110",
42465 => "110111000110011001110010",
42466 => "110110001001000110001000",
42467 => "110110001010110011011110",
42468 => "110111000010100100000000",
42469 => "111000101110011011011101",
42470 => "111011001000001010111010",
42471 => "111101110100010010011000",
42472 => "111111111011010110101101",
42473 => "000001011111001011010110",
42474 => "000011011011111001100110",
42475 => "000101011100011011110000",
42476 => "000110100110010110100010",
42477 => "000111000001101000010011",
42478 => "000111100101011010000101",
42479 => "001001001010111000111010",
42480 => "001011000110111110110111",
42481 => "001100001111011111011000",
42482 => "001100011100100011110000",
42483 => "001011011000010001100011",
42484 => "001001011111110111011011",
42485 => "000111100000000010100110",
42486 => "000100111000110101001101",
42487 => "000001110000100110011100",
42488 => "111110100010000010001001",
42489 => "111100001001011010001111",
42490 => "111011110100101111000000",
42491 => "111101010010010010100001",
42492 => "000000101110110001111011",
42493 => "000101110010111011010011",
42494 => "001010011000000001010110",
42495 => "001101110000111110001100",
42496 => "001111110010001101000010",
42497 => "010000001101000100110010",
42498 => "001110110100110101111000",
42499 => "001010010100000010000110",
42500 => "000011111001011111110000",
42501 => "111111000101000100111101",
42502 => "111100100110000011100010",
42503 => "111011100100000111101000",
42504 => "111011011100011111001111",
42505 => "111011100001011100101000",
42506 => "111011101110100101000010",
42507 => "111100011001010111110100",
42508 => "111101000110000001010100",
42509 => "111101100100111010001111",
42510 => "111110101000010001111011",
42511 => "000000100010100010011000",
42512 => "000001111101001011111100",
42513 => "000001010100010100110001",
42514 => "111111011010111011100010",
42515 => "111110010001011111011101",
42516 => "111101110101110111101010",
42517 => "111101101111110011110000",
42518 => "111110011101011111010101",
42519 => "111111010010111100110010",
42520 => "111111001001000101100000",
42521 => "111101100011001010111101",
42522 => "111011111011101110001110",
42523 => "111100100100010011010000",
42524 => "111110100111111110010100",
42525 => "000000100001000111010010",
42526 => "000010110001110101111010",
42527 => "000101111011101010111101",
42528 => "001000111111101011110111",
42529 => "001001010111111010111011",
42530 => "000111001001010011011010",
42531 => "000101010110010110101011",
42532 => "000011011111110111001010",
42533 => "000000010100001011111110",
42534 => "111101001101101010101010",
42535 => "111010011001011000001100",
42536 => "110111011101111111001100",
42537 => "110100101101100111001110",
42538 => "110010011111110100000000",
42539 => "110001111010001111000010",
42540 => "110011010110110111010100",
42541 => "110110001100001000010010",
42542 => "111001011011010100100100",
42543 => "111100000111111010011010",
42544 => "111110101101011001101110",
42545 => "000001111001111101111101",
42546 => "000101010111110011001111",
42547 => "001000011111011000110001",
42548 => "001010101100000100111110",
42549 => "001100001001110011011010",
42550 => "001101001000100010101110",
42551 => "001100101010100011101100",
42552 => "001010100010101000001111",
42553 => "000111010010010010001000",
42554 => "000010011111100110110110",
42555 => "111101010100100011100010",
42556 => "111010101010001010110100",
42557 => "111011001100110100001010",
42558 => "111101001011100111100000",
42559 => "111110111110011010000110",
42560 => "000000010111011101011000",
42561 => "000001111110000100110100",
42562 => "000011101100111010010010",
42563 => "000100110001000110000110",
42564 => "000100111111100110100110",
42565 => "000100101111111111011110",
42566 => "000011011001110110000011",
42567 => "000000000100110001001101",
42568 => "111011111100101010000100",
42569 => "111001010011001001000110",
42570 => "111000110111110011100010",
42571 => "111000111111100100001011",
42572 => "111000000001011000000000",
42573 => "110111010101001011011011",
42574 => "111000100101100001001110",
42575 => "111010111001010000011010",
42576 => "111100011100101110000110",
42577 => "111100101001100001001101",
42578 => "111101001010101011100101",
42579 => "111110010001110010010110",
42580 => "111101101111000101101100",
42581 => "111011111101101000101001",
42582 => "111010101000101101010100",
42583 => "111010000000010101011001",
42584 => "111001111110111001001101",
42585 => "111001110000101001001101",
42586 => "111001111010101010110110",
42587 => "111011100000011111001100",
42588 => "111101111010001001011011",
42589 => "000000101101101011110110",
42590 => "000010100000111011000011",
42591 => "000010001011100010111000",
42592 => "000000001101111011001100",
42593 => "111100100101110010010110",
42594 => "111000110011101011001111",
42595 => "110101110000010111110010",
42596 => "110010000110010010111100",
42597 => "101110101000111001110100",
42598 => "101100010111010011001000",
42599 => "101100000001000010001000",
42600 => "101111000101001100001010",
42601 => "110100100110101101101011",
42602 => "111011100010111010011100",
42603 => "000011111000110111000110",
42604 => "001100001000101000011110",
42605 => "010001111011011011011010",
42606 => "010011001000010101011100",
42607 => "010000000101011001011100",
42608 => "001010111100110001010110",
42609 => "000100100110110001000001",
42610 => "111101101011101001000010",
42611 => "110111000011111001000110",
42612 => "110001111101111000111100",
42613 => "101111111011110110010000",
42614 => "110000010101110100001110",
42615 => "110001011110001100011010",
42616 => "110011100110101000101110",
42617 => "110111111001001100000111",
42618 => "111101111001101000100100",
42619 => "000011111110001111110010",
42620 => "001000110001100000111011",
42621 => "001011110000110001001110",
42622 => "001101100011110001111100",
42623 => "001110011100110000111000",
42624 => "001101010110111000111000",
42625 => "001010101000110001011000",
42626 => "001000001101000111000101",
42627 => "000110110010011111110111",
42628 => "000101100111011101000101",
42629 => "000011101011001001101111",
42630 => "000001000110101101010111",
42631 => "111110111110010100101101",
42632 => "111101110100000001111111",
42633 => "111101000011110011101100",
42634 => "111011110001000101100001",
42635 => "111010100000101100011111",
42636 => "111010100110111011010100",
42637 => "111011100001011101001101",
42638 => "111100000100011000110010",
42639 => "111100011011101000011000",
42640 => "111101011110011011101000",
42641 => "111111011000001001100110",
42642 => "000001010101010001000011",
42643 => "000010101100010101101001",
42644 => "000011110110111100001000",
42645 => "000101001010001011100100",
42646 => "000101101101001100101100",
42647 => "000100110101101100001001",
42648 => "000011011011011111100110",
42649 => "000010101100010000001110",
42650 => "000011000011010111101001",
42651 => "000011110000110010000100",
42652 => "000011101010110101110101",
42653 => "000010110110011110101110",
42654 => "000010000100110011100000",
42655 => "000001010011111001001101",
42656 => "111111111100101010001101",
42657 => "111110000110110000001101",
42658 => "111100011001000111100100",
42659 => "111010101001110010110000",
42660 => "111001001001011001100100",
42661 => "111000111010011111010010",
42662 => "111010001000010000011101",
42663 => "111100001011111001101101",
42664 => "111110001101110111011010",
42665 => "111111110011010011001110",
42666 => "000001001011000011000110",
42667 => "000010001100010000001111",
42668 => "000010010101011011000101",
42669 => "000000011110001110110110",
42670 => "111100001111100110010110",
42671 => "110111110011110110011011",
42672 => "110101010011001111111110",
42673 => "110101001001100111011100",
42674 => "110110101001110100011110",
42675 => "111000100100011101111010",
42676 => "111010110110100001101101",
42677 => "111110000001111011110010",
42678 => "000001110100001110001000");
signal count : std_logic_vector(16 -1 downto 0) := (others => '0');
begin
	getRomData: process (count)
	begin
		case count is
		when "0000000000000000" => data_out <= rom_array(0);
		when "0000000000000001" => data_out <= rom_array(1);
		when "0000000000000010" => data_out <= rom_array(2);
		when "0000000000000011" => data_out <= rom_array(3);
		when "0000000000000100" => data_out <= rom_array(4);
		when "0000000000000101" => data_out <= rom_array(5);
		when "0000000000000110" => data_out <= rom_array(6);
		when "0000000000000111" => data_out <= rom_array(7);
		when "0000000000001000" => data_out <= rom_array(8);
		when "0000000000001001" => data_out <= rom_array(9);
		when "0000000000001010" => data_out <= rom_array(10);
		when "0000000000001011" => data_out <= rom_array(11);
		when "0000000000001100" => data_out <= rom_array(12);
		when "0000000000001101" => data_out <= rom_array(13);
		when "0000000000001110" => data_out <= rom_array(14);
		when "0000000000001111" => data_out <= rom_array(15);
		when "0000000000010000" => data_out <= rom_array(16);
		when "0000000000010001" => data_out <= rom_array(17);
		when "0000000000010010" => data_out <= rom_array(18);
		when "0000000000010011" => data_out <= rom_array(19);
		when "0000000000010100" => data_out <= rom_array(20);
		when "0000000000010101" => data_out <= rom_array(21);
		when "0000000000010110" => data_out <= rom_array(22);
		when "0000000000010111" => data_out <= rom_array(23);
		when "0000000000011000" => data_out <= rom_array(24);
		when "0000000000011001" => data_out <= rom_array(25);
		when "0000000000011010" => data_out <= rom_array(26);
		when "0000000000011011" => data_out <= rom_array(27);
		when "0000000000011100" => data_out <= rom_array(28);
		when "0000000000011101" => data_out <= rom_array(29);
		when "0000000000011110" => data_out <= rom_array(30);
		when "0000000000011111" => data_out <= rom_array(31);
		when "0000000000100000" => data_out <= rom_array(32);
		when "0000000000100001" => data_out <= rom_array(33);
		when "0000000000100010" => data_out <= rom_array(34);
		when "0000000000100011" => data_out <= rom_array(35);
		when "0000000000100100" => data_out <= rom_array(36);
		when "0000000000100101" => data_out <= rom_array(37);
		when "0000000000100110" => data_out <= rom_array(38);
		when "0000000000100111" => data_out <= rom_array(39);
		when "0000000000101000" => data_out <= rom_array(40);
		when "0000000000101001" => data_out <= rom_array(41);
		when "0000000000101010" => data_out <= rom_array(42);
		when "0000000000101011" => data_out <= rom_array(43);
		when "0000000000101100" => data_out <= rom_array(44);
		when "0000000000101101" => data_out <= rom_array(45);
		when "0000000000101110" => data_out <= rom_array(46);
		when "0000000000101111" => data_out <= rom_array(47);
		when "0000000000110000" => data_out <= rom_array(48);
		when "0000000000110001" => data_out <= rom_array(49);
		when "0000000000110010" => data_out <= rom_array(50);
		when "0000000000110011" => data_out <= rom_array(51);
		when "0000000000110100" => data_out <= rom_array(52);
		when "0000000000110101" => data_out <= rom_array(53);
		when "0000000000110110" => data_out <= rom_array(54);
		when "0000000000110111" => data_out <= rom_array(55);
		when "0000000000111000" => data_out <= rom_array(56);
		when "0000000000111001" => data_out <= rom_array(57);
		when "0000000000111010" => data_out <= rom_array(58);
		when "0000000000111011" => data_out <= rom_array(59);
		when "0000000000111100" => data_out <= rom_array(60);
		when "0000000000111101" => data_out <= rom_array(61);
		when "0000000000111110" => data_out <= rom_array(62);
		when "0000000000111111" => data_out <= rom_array(63);
		when "0000000001000000" => data_out <= rom_array(64);
		when "0000000001000001" => data_out <= rom_array(65);
		when "0000000001000010" => data_out <= rom_array(66);
		when "0000000001000011" => data_out <= rom_array(67);
		when "0000000001000100" => data_out <= rom_array(68);
		when "0000000001000101" => data_out <= rom_array(69);
		when "0000000001000110" => data_out <= rom_array(70);
		when "0000000001000111" => data_out <= rom_array(71);
		when "0000000001001000" => data_out <= rom_array(72);
		when "0000000001001001" => data_out <= rom_array(73);
		when "0000000001001010" => data_out <= rom_array(74);
		when "0000000001001011" => data_out <= rom_array(75);
		when "0000000001001100" => data_out <= rom_array(76);
		when "0000000001001101" => data_out <= rom_array(77);
		when "0000000001001110" => data_out <= rom_array(78);
		when "0000000001001111" => data_out <= rom_array(79);
		when "0000000001010000" => data_out <= rom_array(80);
		when "0000000001010001" => data_out <= rom_array(81);
		when "0000000001010010" => data_out <= rom_array(82);
		when "0000000001010011" => data_out <= rom_array(83);
		when "0000000001010100" => data_out <= rom_array(84);
		when "0000000001010101" => data_out <= rom_array(85);
		when "0000000001010110" => data_out <= rom_array(86);
		when "0000000001010111" => data_out <= rom_array(87);
		when "0000000001011000" => data_out <= rom_array(88);
		when "0000000001011001" => data_out <= rom_array(89);
		when "0000000001011010" => data_out <= rom_array(90);
		when "0000000001011011" => data_out <= rom_array(91);
		when "0000000001011100" => data_out <= rom_array(92);
		when "0000000001011101" => data_out <= rom_array(93);
		when "0000000001011110" => data_out <= rom_array(94);
		when "0000000001011111" => data_out <= rom_array(95);
		when "0000000001100000" => data_out <= rom_array(96);
		when "0000000001100001" => data_out <= rom_array(97);
		when "0000000001100010" => data_out <= rom_array(98);
		when "0000000001100011" => data_out <= rom_array(99);
		when "0000000001100100" => data_out <= rom_array(100);
		when "0000000001100101" => data_out <= rom_array(101);
		when "0000000001100110" => data_out <= rom_array(102);
		when "0000000001100111" => data_out <= rom_array(103);
		when "0000000001101000" => data_out <= rom_array(104);
		when "0000000001101001" => data_out <= rom_array(105);
		when "0000000001101010" => data_out <= rom_array(106);
		when "0000000001101011" => data_out <= rom_array(107);
		when "0000000001101100" => data_out <= rom_array(108);
		when "0000000001101101" => data_out <= rom_array(109);
		when "0000000001101110" => data_out <= rom_array(110);
		when "0000000001101111" => data_out <= rom_array(111);
		when "0000000001110000" => data_out <= rom_array(112);
		when "0000000001110001" => data_out <= rom_array(113);
		when "0000000001110010" => data_out <= rom_array(114);
		when "0000000001110011" => data_out <= rom_array(115);
		when "0000000001110100" => data_out <= rom_array(116);
		when "0000000001110101" => data_out <= rom_array(117);
		when "0000000001110110" => data_out <= rom_array(118);
		when "0000000001110111" => data_out <= rom_array(119);
		when "0000000001111000" => data_out <= rom_array(120);
		when "0000000001111001" => data_out <= rom_array(121);
		when "0000000001111010" => data_out <= rom_array(122);
		when "0000000001111011" => data_out <= rom_array(123);
		when "0000000001111100" => data_out <= rom_array(124);
		when "0000000001111101" => data_out <= rom_array(125);
		when "0000000001111110" => data_out <= rom_array(126);
		when "0000000001111111" => data_out <= rom_array(127);
		when "0000000010000000" => data_out <= rom_array(128);
		when "0000000010000001" => data_out <= rom_array(129);
		when "0000000010000010" => data_out <= rom_array(130);
		when "0000000010000011" => data_out <= rom_array(131);
		when "0000000010000100" => data_out <= rom_array(132);
		when "0000000010000101" => data_out <= rom_array(133);
		when "0000000010000110" => data_out <= rom_array(134);
		when "0000000010000111" => data_out <= rom_array(135);
		when "0000000010001000" => data_out <= rom_array(136);
		when "0000000010001001" => data_out <= rom_array(137);
		when "0000000010001010" => data_out <= rom_array(138);
		when "0000000010001011" => data_out <= rom_array(139);
		when "0000000010001100" => data_out <= rom_array(140);
		when "0000000010001101" => data_out <= rom_array(141);
		when "0000000010001110" => data_out <= rom_array(142);
		when "0000000010001111" => data_out <= rom_array(143);
		when "0000000010010000" => data_out <= rom_array(144);
		when "0000000010010001" => data_out <= rom_array(145);
		when "0000000010010010" => data_out <= rom_array(146);
		when "0000000010010011" => data_out <= rom_array(147);
		when "0000000010010100" => data_out <= rom_array(148);
		when "0000000010010101" => data_out <= rom_array(149);
		when "0000000010010110" => data_out <= rom_array(150);
		when "0000000010010111" => data_out <= rom_array(151);
		when "0000000010011000" => data_out <= rom_array(152);
		when "0000000010011001" => data_out <= rom_array(153);
		when "0000000010011010" => data_out <= rom_array(154);
		when "0000000010011011" => data_out <= rom_array(155);
		when "0000000010011100" => data_out <= rom_array(156);
		when "0000000010011101" => data_out <= rom_array(157);
		when "0000000010011110" => data_out <= rom_array(158);
		when "0000000010011111" => data_out <= rom_array(159);
		when "0000000010100000" => data_out <= rom_array(160);
		when "0000000010100001" => data_out <= rom_array(161);
		when "0000000010100010" => data_out <= rom_array(162);
		when "0000000010100011" => data_out <= rom_array(163);
		when "0000000010100100" => data_out <= rom_array(164);
		when "0000000010100101" => data_out <= rom_array(165);
		when "0000000010100110" => data_out <= rom_array(166);
		when "0000000010100111" => data_out <= rom_array(167);
		when "0000000010101000" => data_out <= rom_array(168);
		when "0000000010101001" => data_out <= rom_array(169);
		when "0000000010101010" => data_out <= rom_array(170);
		when "0000000010101011" => data_out <= rom_array(171);
		when "0000000010101100" => data_out <= rom_array(172);
		when "0000000010101101" => data_out <= rom_array(173);
		when "0000000010101110" => data_out <= rom_array(174);
		when "0000000010101111" => data_out <= rom_array(175);
		when "0000000010110000" => data_out <= rom_array(176);
		when "0000000010110001" => data_out <= rom_array(177);
		when "0000000010110010" => data_out <= rom_array(178);
		when "0000000010110011" => data_out <= rom_array(179);
		when "0000000010110100" => data_out <= rom_array(180);
		when "0000000010110101" => data_out <= rom_array(181);
		when "0000000010110110" => data_out <= rom_array(182);
		when "0000000010110111" => data_out <= rom_array(183);
		when "0000000010111000" => data_out <= rom_array(184);
		when "0000000010111001" => data_out <= rom_array(185);
		when "0000000010111010" => data_out <= rom_array(186);
		when "0000000010111011" => data_out <= rom_array(187);
		when "0000000010111100" => data_out <= rom_array(188);
		when "0000000010111101" => data_out <= rom_array(189);
		when "0000000010111110" => data_out <= rom_array(190);
		when "0000000010111111" => data_out <= rom_array(191);
		when "0000000011000000" => data_out <= rom_array(192);
		when "0000000011000001" => data_out <= rom_array(193);
		when "0000000011000010" => data_out <= rom_array(194);
		when "0000000011000011" => data_out <= rom_array(195);
		when "0000000011000100" => data_out <= rom_array(196);
		when "0000000011000101" => data_out <= rom_array(197);
		when "0000000011000110" => data_out <= rom_array(198);
		when "0000000011000111" => data_out <= rom_array(199);
		when "0000000011001000" => data_out <= rom_array(200);
		when "0000000011001001" => data_out <= rom_array(201);
		when "0000000011001010" => data_out <= rom_array(202);
		when "0000000011001011" => data_out <= rom_array(203);
		when "0000000011001100" => data_out <= rom_array(204);
		when "0000000011001101" => data_out <= rom_array(205);
		when "0000000011001110" => data_out <= rom_array(206);
		when "0000000011001111" => data_out <= rom_array(207);
		when "0000000011010000" => data_out <= rom_array(208);
		when "0000000011010001" => data_out <= rom_array(209);
		when "0000000011010010" => data_out <= rom_array(210);
		when "0000000011010011" => data_out <= rom_array(211);
		when "0000000011010100" => data_out <= rom_array(212);
		when "0000000011010101" => data_out <= rom_array(213);
		when "0000000011010110" => data_out <= rom_array(214);
		when "0000000011010111" => data_out <= rom_array(215);
		when "0000000011011000" => data_out <= rom_array(216);
		when "0000000011011001" => data_out <= rom_array(217);
		when "0000000011011010" => data_out <= rom_array(218);
		when "0000000011011011" => data_out <= rom_array(219);
		when "0000000011011100" => data_out <= rom_array(220);
		when "0000000011011101" => data_out <= rom_array(221);
		when "0000000011011110" => data_out <= rom_array(222);
		when "0000000011011111" => data_out <= rom_array(223);
		when "0000000011100000" => data_out <= rom_array(224);
		when "0000000011100001" => data_out <= rom_array(225);
		when "0000000011100010" => data_out <= rom_array(226);
		when "0000000011100011" => data_out <= rom_array(227);
		when "0000000011100100" => data_out <= rom_array(228);
		when "0000000011100101" => data_out <= rom_array(229);
		when "0000000011100110" => data_out <= rom_array(230);
		when "0000000011100111" => data_out <= rom_array(231);
		when "0000000011101000" => data_out <= rom_array(232);
		when "0000000011101001" => data_out <= rom_array(233);
		when "0000000011101010" => data_out <= rom_array(234);
		when "0000000011101011" => data_out <= rom_array(235);
		when "0000000011101100" => data_out <= rom_array(236);
		when "0000000011101101" => data_out <= rom_array(237);
		when "0000000011101110" => data_out <= rom_array(238);
		when "0000000011101111" => data_out <= rom_array(239);
		when "0000000011110000" => data_out <= rom_array(240);
		when "0000000011110001" => data_out <= rom_array(241);
		when "0000000011110010" => data_out <= rom_array(242);
		when "0000000011110011" => data_out <= rom_array(243);
		when "0000000011110100" => data_out <= rom_array(244);
		when "0000000011110101" => data_out <= rom_array(245);
		when "0000000011110110" => data_out <= rom_array(246);
		when "0000000011110111" => data_out <= rom_array(247);
		when "0000000011111000" => data_out <= rom_array(248);
		when "0000000011111001" => data_out <= rom_array(249);
		when "0000000011111010" => data_out <= rom_array(250);
		when "0000000011111011" => data_out <= rom_array(251);
		when "0000000011111100" => data_out <= rom_array(252);
		when "0000000011111101" => data_out <= rom_array(253);
		when "0000000011111110" => data_out <= rom_array(254);
		when "0000000011111111" => data_out <= rom_array(255);
		when "0000000100000000" => data_out <= rom_array(256);
		when "0000000100000001" => data_out <= rom_array(257);
		when "0000000100000010" => data_out <= rom_array(258);
		when "0000000100000011" => data_out <= rom_array(259);
		when "0000000100000100" => data_out <= rom_array(260);
		when "0000000100000101" => data_out <= rom_array(261);
		when "0000000100000110" => data_out <= rom_array(262);
		when "0000000100000111" => data_out <= rom_array(263);
		when "0000000100001000" => data_out <= rom_array(264);
		when "0000000100001001" => data_out <= rom_array(265);
		when "0000000100001010" => data_out <= rom_array(266);
		when "0000000100001011" => data_out <= rom_array(267);
		when "0000000100001100" => data_out <= rom_array(268);
		when "0000000100001101" => data_out <= rom_array(269);
		when "0000000100001110" => data_out <= rom_array(270);
		when "0000000100001111" => data_out <= rom_array(271);
		when "0000000100010000" => data_out <= rom_array(272);
		when "0000000100010001" => data_out <= rom_array(273);
		when "0000000100010010" => data_out <= rom_array(274);
		when "0000000100010011" => data_out <= rom_array(275);
		when "0000000100010100" => data_out <= rom_array(276);
		when "0000000100010101" => data_out <= rom_array(277);
		when "0000000100010110" => data_out <= rom_array(278);
		when "0000000100010111" => data_out <= rom_array(279);
		when "0000000100011000" => data_out <= rom_array(280);
		when "0000000100011001" => data_out <= rom_array(281);
		when "0000000100011010" => data_out <= rom_array(282);
		when "0000000100011011" => data_out <= rom_array(283);
		when "0000000100011100" => data_out <= rom_array(284);
		when "0000000100011101" => data_out <= rom_array(285);
		when "0000000100011110" => data_out <= rom_array(286);
		when "0000000100011111" => data_out <= rom_array(287);
		when "0000000100100000" => data_out <= rom_array(288);
		when "0000000100100001" => data_out <= rom_array(289);
		when "0000000100100010" => data_out <= rom_array(290);
		when "0000000100100011" => data_out <= rom_array(291);
		when "0000000100100100" => data_out <= rom_array(292);
		when "0000000100100101" => data_out <= rom_array(293);
		when "0000000100100110" => data_out <= rom_array(294);
		when "0000000100100111" => data_out <= rom_array(295);
		when "0000000100101000" => data_out <= rom_array(296);
		when "0000000100101001" => data_out <= rom_array(297);
		when "0000000100101010" => data_out <= rom_array(298);
		when "0000000100101011" => data_out <= rom_array(299);
		when "0000000100101100" => data_out <= rom_array(300);
		when "0000000100101101" => data_out <= rom_array(301);
		when "0000000100101110" => data_out <= rom_array(302);
		when "0000000100101111" => data_out <= rom_array(303);
		when "0000000100110000" => data_out <= rom_array(304);
		when "0000000100110001" => data_out <= rom_array(305);
		when "0000000100110010" => data_out <= rom_array(306);
		when "0000000100110011" => data_out <= rom_array(307);
		when "0000000100110100" => data_out <= rom_array(308);
		when "0000000100110101" => data_out <= rom_array(309);
		when "0000000100110110" => data_out <= rom_array(310);
		when "0000000100110111" => data_out <= rom_array(311);
		when "0000000100111000" => data_out <= rom_array(312);
		when "0000000100111001" => data_out <= rom_array(313);
		when "0000000100111010" => data_out <= rom_array(314);
		when "0000000100111011" => data_out <= rom_array(315);
		when "0000000100111100" => data_out <= rom_array(316);
		when "0000000100111101" => data_out <= rom_array(317);
		when "0000000100111110" => data_out <= rom_array(318);
		when "0000000100111111" => data_out <= rom_array(319);
		when "0000000101000000" => data_out <= rom_array(320);
		when "0000000101000001" => data_out <= rom_array(321);
		when "0000000101000010" => data_out <= rom_array(322);
		when "0000000101000011" => data_out <= rom_array(323);
		when "0000000101000100" => data_out <= rom_array(324);
		when "0000000101000101" => data_out <= rom_array(325);
		when "0000000101000110" => data_out <= rom_array(326);
		when "0000000101000111" => data_out <= rom_array(327);
		when "0000000101001000" => data_out <= rom_array(328);
		when "0000000101001001" => data_out <= rom_array(329);
		when "0000000101001010" => data_out <= rom_array(330);
		when "0000000101001011" => data_out <= rom_array(331);
		when "0000000101001100" => data_out <= rom_array(332);
		when "0000000101001101" => data_out <= rom_array(333);
		when "0000000101001110" => data_out <= rom_array(334);
		when "0000000101001111" => data_out <= rom_array(335);
		when "0000000101010000" => data_out <= rom_array(336);
		when "0000000101010001" => data_out <= rom_array(337);
		when "0000000101010010" => data_out <= rom_array(338);
		when "0000000101010011" => data_out <= rom_array(339);
		when "0000000101010100" => data_out <= rom_array(340);
		when "0000000101010101" => data_out <= rom_array(341);
		when "0000000101010110" => data_out <= rom_array(342);
		when "0000000101010111" => data_out <= rom_array(343);
		when "0000000101011000" => data_out <= rom_array(344);
		when "0000000101011001" => data_out <= rom_array(345);
		when "0000000101011010" => data_out <= rom_array(346);
		when "0000000101011011" => data_out <= rom_array(347);
		when "0000000101011100" => data_out <= rom_array(348);
		when "0000000101011101" => data_out <= rom_array(349);
		when "0000000101011110" => data_out <= rom_array(350);
		when "0000000101011111" => data_out <= rom_array(351);
		when "0000000101100000" => data_out <= rom_array(352);
		when "0000000101100001" => data_out <= rom_array(353);
		when "0000000101100010" => data_out <= rom_array(354);
		when "0000000101100011" => data_out <= rom_array(355);
		when "0000000101100100" => data_out <= rom_array(356);
		when "0000000101100101" => data_out <= rom_array(357);
		when "0000000101100110" => data_out <= rom_array(358);
		when "0000000101100111" => data_out <= rom_array(359);
		when "0000000101101000" => data_out <= rom_array(360);
		when "0000000101101001" => data_out <= rom_array(361);
		when "0000000101101010" => data_out <= rom_array(362);
		when "0000000101101011" => data_out <= rom_array(363);
		when "0000000101101100" => data_out <= rom_array(364);
		when "0000000101101101" => data_out <= rom_array(365);
		when "0000000101101110" => data_out <= rom_array(366);
		when "0000000101101111" => data_out <= rom_array(367);
		when "0000000101110000" => data_out <= rom_array(368);
		when "0000000101110001" => data_out <= rom_array(369);
		when "0000000101110010" => data_out <= rom_array(370);
		when "0000000101110011" => data_out <= rom_array(371);
		when "0000000101110100" => data_out <= rom_array(372);
		when "0000000101110101" => data_out <= rom_array(373);
		when "0000000101110110" => data_out <= rom_array(374);
		when "0000000101110111" => data_out <= rom_array(375);
		when "0000000101111000" => data_out <= rom_array(376);
		when "0000000101111001" => data_out <= rom_array(377);
		when "0000000101111010" => data_out <= rom_array(378);
		when "0000000101111011" => data_out <= rom_array(379);
		when "0000000101111100" => data_out <= rom_array(380);
		when "0000000101111101" => data_out <= rom_array(381);
		when "0000000101111110" => data_out <= rom_array(382);
		when "0000000101111111" => data_out <= rom_array(383);
		when "0000000110000000" => data_out <= rom_array(384);
		when "0000000110000001" => data_out <= rom_array(385);
		when "0000000110000010" => data_out <= rom_array(386);
		when "0000000110000011" => data_out <= rom_array(387);
		when "0000000110000100" => data_out <= rom_array(388);
		when "0000000110000101" => data_out <= rom_array(389);
		when "0000000110000110" => data_out <= rom_array(390);
		when "0000000110000111" => data_out <= rom_array(391);
		when "0000000110001000" => data_out <= rom_array(392);
		when "0000000110001001" => data_out <= rom_array(393);
		when "0000000110001010" => data_out <= rom_array(394);
		when "0000000110001011" => data_out <= rom_array(395);
		when "0000000110001100" => data_out <= rom_array(396);
		when "0000000110001101" => data_out <= rom_array(397);
		when "0000000110001110" => data_out <= rom_array(398);
		when "0000000110001111" => data_out <= rom_array(399);
		when "0000000110010000" => data_out <= rom_array(400);
		when "0000000110010001" => data_out <= rom_array(401);
		when "0000000110010010" => data_out <= rom_array(402);
		when "0000000110010011" => data_out <= rom_array(403);
		when "0000000110010100" => data_out <= rom_array(404);
		when "0000000110010101" => data_out <= rom_array(405);
		when "0000000110010110" => data_out <= rom_array(406);
		when "0000000110010111" => data_out <= rom_array(407);
		when "0000000110011000" => data_out <= rom_array(408);
		when "0000000110011001" => data_out <= rom_array(409);
		when "0000000110011010" => data_out <= rom_array(410);
		when "0000000110011011" => data_out <= rom_array(411);
		when "0000000110011100" => data_out <= rom_array(412);
		when "0000000110011101" => data_out <= rom_array(413);
		when "0000000110011110" => data_out <= rom_array(414);
		when "0000000110011111" => data_out <= rom_array(415);
		when "0000000110100000" => data_out <= rom_array(416);
		when "0000000110100001" => data_out <= rom_array(417);
		when "0000000110100010" => data_out <= rom_array(418);
		when "0000000110100011" => data_out <= rom_array(419);
		when "0000000110100100" => data_out <= rom_array(420);
		when "0000000110100101" => data_out <= rom_array(421);
		when "0000000110100110" => data_out <= rom_array(422);
		when "0000000110100111" => data_out <= rom_array(423);
		when "0000000110101000" => data_out <= rom_array(424);
		when "0000000110101001" => data_out <= rom_array(425);
		when "0000000110101010" => data_out <= rom_array(426);
		when "0000000110101011" => data_out <= rom_array(427);
		when "0000000110101100" => data_out <= rom_array(428);
		when "0000000110101101" => data_out <= rom_array(429);
		when "0000000110101110" => data_out <= rom_array(430);
		when "0000000110101111" => data_out <= rom_array(431);
		when "0000000110110000" => data_out <= rom_array(432);
		when "0000000110110001" => data_out <= rom_array(433);
		when "0000000110110010" => data_out <= rom_array(434);
		when "0000000110110011" => data_out <= rom_array(435);
		when "0000000110110100" => data_out <= rom_array(436);
		when "0000000110110101" => data_out <= rom_array(437);
		when "0000000110110110" => data_out <= rom_array(438);
		when "0000000110110111" => data_out <= rom_array(439);
		when "0000000110111000" => data_out <= rom_array(440);
		when "0000000110111001" => data_out <= rom_array(441);
		when "0000000110111010" => data_out <= rom_array(442);
		when "0000000110111011" => data_out <= rom_array(443);
		when "0000000110111100" => data_out <= rom_array(444);
		when "0000000110111101" => data_out <= rom_array(445);
		when "0000000110111110" => data_out <= rom_array(446);
		when "0000000110111111" => data_out <= rom_array(447);
		when "0000000111000000" => data_out <= rom_array(448);
		when "0000000111000001" => data_out <= rom_array(449);
		when "0000000111000010" => data_out <= rom_array(450);
		when "0000000111000011" => data_out <= rom_array(451);
		when "0000000111000100" => data_out <= rom_array(452);
		when "0000000111000101" => data_out <= rom_array(453);
		when "0000000111000110" => data_out <= rom_array(454);
		when "0000000111000111" => data_out <= rom_array(455);
		when "0000000111001000" => data_out <= rom_array(456);
		when "0000000111001001" => data_out <= rom_array(457);
		when "0000000111001010" => data_out <= rom_array(458);
		when "0000000111001011" => data_out <= rom_array(459);
		when "0000000111001100" => data_out <= rom_array(460);
		when "0000000111001101" => data_out <= rom_array(461);
		when "0000000111001110" => data_out <= rom_array(462);
		when "0000000111001111" => data_out <= rom_array(463);
		when "0000000111010000" => data_out <= rom_array(464);
		when "0000000111010001" => data_out <= rom_array(465);
		when "0000000111010010" => data_out <= rom_array(466);
		when "0000000111010011" => data_out <= rom_array(467);
		when "0000000111010100" => data_out <= rom_array(468);
		when "0000000111010101" => data_out <= rom_array(469);
		when "0000000111010110" => data_out <= rom_array(470);
		when "0000000111010111" => data_out <= rom_array(471);
		when "0000000111011000" => data_out <= rom_array(472);
		when "0000000111011001" => data_out <= rom_array(473);
		when "0000000111011010" => data_out <= rom_array(474);
		when "0000000111011011" => data_out <= rom_array(475);
		when "0000000111011100" => data_out <= rom_array(476);
		when "0000000111011101" => data_out <= rom_array(477);
		when "0000000111011110" => data_out <= rom_array(478);
		when "0000000111011111" => data_out <= rom_array(479);
		when "0000000111100000" => data_out <= rom_array(480);
		when "0000000111100001" => data_out <= rom_array(481);
		when "0000000111100010" => data_out <= rom_array(482);
		when "0000000111100011" => data_out <= rom_array(483);
		when "0000000111100100" => data_out <= rom_array(484);
		when "0000000111100101" => data_out <= rom_array(485);
		when "0000000111100110" => data_out <= rom_array(486);
		when "0000000111100111" => data_out <= rom_array(487);
		when "0000000111101000" => data_out <= rom_array(488);
		when "0000000111101001" => data_out <= rom_array(489);
		when "0000000111101010" => data_out <= rom_array(490);
		when "0000000111101011" => data_out <= rom_array(491);
		when "0000000111101100" => data_out <= rom_array(492);
		when "0000000111101101" => data_out <= rom_array(493);
		when "0000000111101110" => data_out <= rom_array(494);
		when "0000000111101111" => data_out <= rom_array(495);
		when "0000000111110000" => data_out <= rom_array(496);
		when "0000000111110001" => data_out <= rom_array(497);
		when "0000000111110010" => data_out <= rom_array(498);
		when "0000000111110011" => data_out <= rom_array(499);
		when "0000000111110100" => data_out <= rom_array(500);
		when "0000000111110101" => data_out <= rom_array(501);
		when "0000000111110110" => data_out <= rom_array(502);
		when "0000000111110111" => data_out <= rom_array(503);
		when "0000000111111000" => data_out <= rom_array(504);
		when "0000000111111001" => data_out <= rom_array(505);
		when "0000000111111010" => data_out <= rom_array(506);
		when "0000000111111011" => data_out <= rom_array(507);
		when "0000000111111100" => data_out <= rom_array(508);
		when "0000000111111101" => data_out <= rom_array(509);
		when "0000000111111110" => data_out <= rom_array(510);
		when "0000000111111111" => data_out <= rom_array(511);
		when "0000001000000000" => data_out <= rom_array(512);
		when "0000001000000001" => data_out <= rom_array(513);
		when "0000001000000010" => data_out <= rom_array(514);
		when "0000001000000011" => data_out <= rom_array(515);
		when "0000001000000100" => data_out <= rom_array(516);
		when "0000001000000101" => data_out <= rom_array(517);
		when "0000001000000110" => data_out <= rom_array(518);
		when "0000001000000111" => data_out <= rom_array(519);
		when "0000001000001000" => data_out <= rom_array(520);
		when "0000001000001001" => data_out <= rom_array(521);
		when "0000001000001010" => data_out <= rom_array(522);
		when "0000001000001011" => data_out <= rom_array(523);
		when "0000001000001100" => data_out <= rom_array(524);
		when "0000001000001101" => data_out <= rom_array(525);
		when "0000001000001110" => data_out <= rom_array(526);
		when "0000001000001111" => data_out <= rom_array(527);
		when "0000001000010000" => data_out <= rom_array(528);
		when "0000001000010001" => data_out <= rom_array(529);
		when "0000001000010010" => data_out <= rom_array(530);
		when "0000001000010011" => data_out <= rom_array(531);
		when "0000001000010100" => data_out <= rom_array(532);
		when "0000001000010101" => data_out <= rom_array(533);
		when "0000001000010110" => data_out <= rom_array(534);
		when "0000001000010111" => data_out <= rom_array(535);
		when "0000001000011000" => data_out <= rom_array(536);
		when "0000001000011001" => data_out <= rom_array(537);
		when "0000001000011010" => data_out <= rom_array(538);
		when "0000001000011011" => data_out <= rom_array(539);
		when "0000001000011100" => data_out <= rom_array(540);
		when "0000001000011101" => data_out <= rom_array(541);
		when "0000001000011110" => data_out <= rom_array(542);
		when "0000001000011111" => data_out <= rom_array(543);
		when "0000001000100000" => data_out <= rom_array(544);
		when "0000001000100001" => data_out <= rom_array(545);
		when "0000001000100010" => data_out <= rom_array(546);
		when "0000001000100011" => data_out <= rom_array(547);
		when "0000001000100100" => data_out <= rom_array(548);
		when "0000001000100101" => data_out <= rom_array(549);
		when "0000001000100110" => data_out <= rom_array(550);
		when "0000001000100111" => data_out <= rom_array(551);
		when "0000001000101000" => data_out <= rom_array(552);
		when "0000001000101001" => data_out <= rom_array(553);
		when "0000001000101010" => data_out <= rom_array(554);
		when "0000001000101011" => data_out <= rom_array(555);
		when "0000001000101100" => data_out <= rom_array(556);
		when "0000001000101101" => data_out <= rom_array(557);
		when "0000001000101110" => data_out <= rom_array(558);
		when "0000001000101111" => data_out <= rom_array(559);
		when "0000001000110000" => data_out <= rom_array(560);
		when "0000001000110001" => data_out <= rom_array(561);
		when "0000001000110010" => data_out <= rom_array(562);
		when "0000001000110011" => data_out <= rom_array(563);
		when "0000001000110100" => data_out <= rom_array(564);
		when "0000001000110101" => data_out <= rom_array(565);
		when "0000001000110110" => data_out <= rom_array(566);
		when "0000001000110111" => data_out <= rom_array(567);
		when "0000001000111000" => data_out <= rom_array(568);
		when "0000001000111001" => data_out <= rom_array(569);
		when "0000001000111010" => data_out <= rom_array(570);
		when "0000001000111011" => data_out <= rom_array(571);
		when "0000001000111100" => data_out <= rom_array(572);
		when "0000001000111101" => data_out <= rom_array(573);
		when "0000001000111110" => data_out <= rom_array(574);
		when "0000001000111111" => data_out <= rom_array(575);
		when "0000001001000000" => data_out <= rom_array(576);
		when "0000001001000001" => data_out <= rom_array(577);
		when "0000001001000010" => data_out <= rom_array(578);
		when "0000001001000011" => data_out <= rom_array(579);
		when "0000001001000100" => data_out <= rom_array(580);
		when "0000001001000101" => data_out <= rom_array(581);
		when "0000001001000110" => data_out <= rom_array(582);
		when "0000001001000111" => data_out <= rom_array(583);
		when "0000001001001000" => data_out <= rom_array(584);
		when "0000001001001001" => data_out <= rom_array(585);
		when "0000001001001010" => data_out <= rom_array(586);
		when "0000001001001011" => data_out <= rom_array(587);
		when "0000001001001100" => data_out <= rom_array(588);
		when "0000001001001101" => data_out <= rom_array(589);
		when "0000001001001110" => data_out <= rom_array(590);
		when "0000001001001111" => data_out <= rom_array(591);
		when "0000001001010000" => data_out <= rom_array(592);
		when "0000001001010001" => data_out <= rom_array(593);
		when "0000001001010010" => data_out <= rom_array(594);
		when "0000001001010011" => data_out <= rom_array(595);
		when "0000001001010100" => data_out <= rom_array(596);
		when "0000001001010101" => data_out <= rom_array(597);
		when "0000001001010110" => data_out <= rom_array(598);
		when "0000001001010111" => data_out <= rom_array(599);
		when "0000001001011000" => data_out <= rom_array(600);
		when "0000001001011001" => data_out <= rom_array(601);
		when "0000001001011010" => data_out <= rom_array(602);
		when "0000001001011011" => data_out <= rom_array(603);
		when "0000001001011100" => data_out <= rom_array(604);
		when "0000001001011101" => data_out <= rom_array(605);
		when "0000001001011110" => data_out <= rom_array(606);
		when "0000001001011111" => data_out <= rom_array(607);
		when "0000001001100000" => data_out <= rom_array(608);
		when "0000001001100001" => data_out <= rom_array(609);
		when "0000001001100010" => data_out <= rom_array(610);
		when "0000001001100011" => data_out <= rom_array(611);
		when "0000001001100100" => data_out <= rom_array(612);
		when "0000001001100101" => data_out <= rom_array(613);
		when "0000001001100110" => data_out <= rom_array(614);
		when "0000001001100111" => data_out <= rom_array(615);
		when "0000001001101000" => data_out <= rom_array(616);
		when "0000001001101001" => data_out <= rom_array(617);
		when "0000001001101010" => data_out <= rom_array(618);
		when "0000001001101011" => data_out <= rom_array(619);
		when "0000001001101100" => data_out <= rom_array(620);
		when "0000001001101101" => data_out <= rom_array(621);
		when "0000001001101110" => data_out <= rom_array(622);
		when "0000001001101111" => data_out <= rom_array(623);
		when "0000001001110000" => data_out <= rom_array(624);
		when "0000001001110001" => data_out <= rom_array(625);
		when "0000001001110010" => data_out <= rom_array(626);
		when "0000001001110011" => data_out <= rom_array(627);
		when "0000001001110100" => data_out <= rom_array(628);
		when "0000001001110101" => data_out <= rom_array(629);
		when "0000001001110110" => data_out <= rom_array(630);
		when "0000001001110111" => data_out <= rom_array(631);
		when "0000001001111000" => data_out <= rom_array(632);
		when "0000001001111001" => data_out <= rom_array(633);
		when "0000001001111010" => data_out <= rom_array(634);
		when "0000001001111011" => data_out <= rom_array(635);
		when "0000001001111100" => data_out <= rom_array(636);
		when "0000001001111101" => data_out <= rom_array(637);
		when "0000001001111110" => data_out <= rom_array(638);
		when "0000001001111111" => data_out <= rom_array(639);
		when "0000001010000000" => data_out <= rom_array(640);
		when "0000001010000001" => data_out <= rom_array(641);
		when "0000001010000010" => data_out <= rom_array(642);
		when "0000001010000011" => data_out <= rom_array(643);
		when "0000001010000100" => data_out <= rom_array(644);
		when "0000001010000101" => data_out <= rom_array(645);
		when "0000001010000110" => data_out <= rom_array(646);
		when "0000001010000111" => data_out <= rom_array(647);
		when "0000001010001000" => data_out <= rom_array(648);
		when "0000001010001001" => data_out <= rom_array(649);
		when "0000001010001010" => data_out <= rom_array(650);
		when "0000001010001011" => data_out <= rom_array(651);
		when "0000001010001100" => data_out <= rom_array(652);
		when "0000001010001101" => data_out <= rom_array(653);
		when "0000001010001110" => data_out <= rom_array(654);
		when "0000001010001111" => data_out <= rom_array(655);
		when "0000001010010000" => data_out <= rom_array(656);
		when "0000001010010001" => data_out <= rom_array(657);
		when "0000001010010010" => data_out <= rom_array(658);
		when "0000001010010011" => data_out <= rom_array(659);
		when "0000001010010100" => data_out <= rom_array(660);
		when "0000001010010101" => data_out <= rom_array(661);
		when "0000001010010110" => data_out <= rom_array(662);
		when "0000001010010111" => data_out <= rom_array(663);
		when "0000001010011000" => data_out <= rom_array(664);
		when "0000001010011001" => data_out <= rom_array(665);
		when "0000001010011010" => data_out <= rom_array(666);
		when "0000001010011011" => data_out <= rom_array(667);
		when "0000001010011100" => data_out <= rom_array(668);
		when "0000001010011101" => data_out <= rom_array(669);
		when "0000001010011110" => data_out <= rom_array(670);
		when "0000001010011111" => data_out <= rom_array(671);
		when "0000001010100000" => data_out <= rom_array(672);
		when "0000001010100001" => data_out <= rom_array(673);
		when "0000001010100010" => data_out <= rom_array(674);
		when "0000001010100011" => data_out <= rom_array(675);
		when "0000001010100100" => data_out <= rom_array(676);
		when "0000001010100101" => data_out <= rom_array(677);
		when "0000001010100110" => data_out <= rom_array(678);
		when "0000001010100111" => data_out <= rom_array(679);
		when "0000001010101000" => data_out <= rom_array(680);
		when "0000001010101001" => data_out <= rom_array(681);
		when "0000001010101010" => data_out <= rom_array(682);
		when "0000001010101011" => data_out <= rom_array(683);
		when "0000001010101100" => data_out <= rom_array(684);
		when "0000001010101101" => data_out <= rom_array(685);
		when "0000001010101110" => data_out <= rom_array(686);
		when "0000001010101111" => data_out <= rom_array(687);
		when "0000001010110000" => data_out <= rom_array(688);
		when "0000001010110001" => data_out <= rom_array(689);
		when "0000001010110010" => data_out <= rom_array(690);
		when "0000001010110011" => data_out <= rom_array(691);
		when "0000001010110100" => data_out <= rom_array(692);
		when "0000001010110101" => data_out <= rom_array(693);
		when "0000001010110110" => data_out <= rom_array(694);
		when "0000001010110111" => data_out <= rom_array(695);
		when "0000001010111000" => data_out <= rom_array(696);
		when "0000001010111001" => data_out <= rom_array(697);
		when "0000001010111010" => data_out <= rom_array(698);
		when "0000001010111011" => data_out <= rom_array(699);
		when "0000001010111100" => data_out <= rom_array(700);
		when "0000001010111101" => data_out <= rom_array(701);
		when "0000001010111110" => data_out <= rom_array(702);
		when "0000001010111111" => data_out <= rom_array(703);
		when "0000001011000000" => data_out <= rom_array(704);
		when "0000001011000001" => data_out <= rom_array(705);
		when "0000001011000010" => data_out <= rom_array(706);
		when "0000001011000011" => data_out <= rom_array(707);
		when "0000001011000100" => data_out <= rom_array(708);
		when "0000001011000101" => data_out <= rom_array(709);
		when "0000001011000110" => data_out <= rom_array(710);
		when "0000001011000111" => data_out <= rom_array(711);
		when "0000001011001000" => data_out <= rom_array(712);
		when "0000001011001001" => data_out <= rom_array(713);
		when "0000001011001010" => data_out <= rom_array(714);
		when "0000001011001011" => data_out <= rom_array(715);
		when "0000001011001100" => data_out <= rom_array(716);
		when "0000001011001101" => data_out <= rom_array(717);
		when "0000001011001110" => data_out <= rom_array(718);
		when "0000001011001111" => data_out <= rom_array(719);
		when "0000001011010000" => data_out <= rom_array(720);
		when "0000001011010001" => data_out <= rom_array(721);
		when "0000001011010010" => data_out <= rom_array(722);
		when "0000001011010011" => data_out <= rom_array(723);
		when "0000001011010100" => data_out <= rom_array(724);
		when "0000001011010101" => data_out <= rom_array(725);
		when "0000001011010110" => data_out <= rom_array(726);
		when "0000001011010111" => data_out <= rom_array(727);
		when "0000001011011000" => data_out <= rom_array(728);
		when "0000001011011001" => data_out <= rom_array(729);
		when "0000001011011010" => data_out <= rom_array(730);
		when "0000001011011011" => data_out <= rom_array(731);
		when "0000001011011100" => data_out <= rom_array(732);
		when "0000001011011101" => data_out <= rom_array(733);
		when "0000001011011110" => data_out <= rom_array(734);
		when "0000001011011111" => data_out <= rom_array(735);
		when "0000001011100000" => data_out <= rom_array(736);
		when "0000001011100001" => data_out <= rom_array(737);
		when "0000001011100010" => data_out <= rom_array(738);
		when "0000001011100011" => data_out <= rom_array(739);
		when "0000001011100100" => data_out <= rom_array(740);
		when "0000001011100101" => data_out <= rom_array(741);
		when "0000001011100110" => data_out <= rom_array(742);
		when "0000001011100111" => data_out <= rom_array(743);
		when "0000001011101000" => data_out <= rom_array(744);
		when "0000001011101001" => data_out <= rom_array(745);
		when "0000001011101010" => data_out <= rom_array(746);
		when "0000001011101011" => data_out <= rom_array(747);
		when "0000001011101100" => data_out <= rom_array(748);
		when "0000001011101101" => data_out <= rom_array(749);
		when "0000001011101110" => data_out <= rom_array(750);
		when "0000001011101111" => data_out <= rom_array(751);
		when "0000001011110000" => data_out <= rom_array(752);
		when "0000001011110001" => data_out <= rom_array(753);
		when "0000001011110010" => data_out <= rom_array(754);
		when "0000001011110011" => data_out <= rom_array(755);
		when "0000001011110100" => data_out <= rom_array(756);
		when "0000001011110101" => data_out <= rom_array(757);
		when "0000001011110110" => data_out <= rom_array(758);
		when "0000001011110111" => data_out <= rom_array(759);
		when "0000001011111000" => data_out <= rom_array(760);
		when "0000001011111001" => data_out <= rom_array(761);
		when "0000001011111010" => data_out <= rom_array(762);
		when "0000001011111011" => data_out <= rom_array(763);
		when "0000001011111100" => data_out <= rom_array(764);
		when "0000001011111101" => data_out <= rom_array(765);
		when "0000001011111110" => data_out <= rom_array(766);
		when "0000001011111111" => data_out <= rom_array(767);
		when "0000001100000000" => data_out <= rom_array(768);
		when "0000001100000001" => data_out <= rom_array(769);
		when "0000001100000010" => data_out <= rom_array(770);
		when "0000001100000011" => data_out <= rom_array(771);
		when "0000001100000100" => data_out <= rom_array(772);
		when "0000001100000101" => data_out <= rom_array(773);
		when "0000001100000110" => data_out <= rom_array(774);
		when "0000001100000111" => data_out <= rom_array(775);
		when "0000001100001000" => data_out <= rom_array(776);
		when "0000001100001001" => data_out <= rom_array(777);
		when "0000001100001010" => data_out <= rom_array(778);
		when "0000001100001011" => data_out <= rom_array(779);
		when "0000001100001100" => data_out <= rom_array(780);
		when "0000001100001101" => data_out <= rom_array(781);
		when "0000001100001110" => data_out <= rom_array(782);
		when "0000001100001111" => data_out <= rom_array(783);
		when "0000001100010000" => data_out <= rom_array(784);
		when "0000001100010001" => data_out <= rom_array(785);
		when "0000001100010010" => data_out <= rom_array(786);
		when "0000001100010011" => data_out <= rom_array(787);
		when "0000001100010100" => data_out <= rom_array(788);
		when "0000001100010101" => data_out <= rom_array(789);
		when "0000001100010110" => data_out <= rom_array(790);
		when "0000001100010111" => data_out <= rom_array(791);
		when "0000001100011000" => data_out <= rom_array(792);
		when "0000001100011001" => data_out <= rom_array(793);
		when "0000001100011010" => data_out <= rom_array(794);
		when "0000001100011011" => data_out <= rom_array(795);
		when "0000001100011100" => data_out <= rom_array(796);
		when "0000001100011101" => data_out <= rom_array(797);
		when "0000001100011110" => data_out <= rom_array(798);
		when "0000001100011111" => data_out <= rom_array(799);
		when "0000001100100000" => data_out <= rom_array(800);
		when "0000001100100001" => data_out <= rom_array(801);
		when "0000001100100010" => data_out <= rom_array(802);
		when "0000001100100011" => data_out <= rom_array(803);
		when "0000001100100100" => data_out <= rom_array(804);
		when "0000001100100101" => data_out <= rom_array(805);
		when "0000001100100110" => data_out <= rom_array(806);
		when "0000001100100111" => data_out <= rom_array(807);
		when "0000001100101000" => data_out <= rom_array(808);
		when "0000001100101001" => data_out <= rom_array(809);
		when "0000001100101010" => data_out <= rom_array(810);
		when "0000001100101011" => data_out <= rom_array(811);
		when "0000001100101100" => data_out <= rom_array(812);
		when "0000001100101101" => data_out <= rom_array(813);
		when "0000001100101110" => data_out <= rom_array(814);
		when "0000001100101111" => data_out <= rom_array(815);
		when "0000001100110000" => data_out <= rom_array(816);
		when "0000001100110001" => data_out <= rom_array(817);
		when "0000001100110010" => data_out <= rom_array(818);
		when "0000001100110011" => data_out <= rom_array(819);
		when "0000001100110100" => data_out <= rom_array(820);
		when "0000001100110101" => data_out <= rom_array(821);
		when "0000001100110110" => data_out <= rom_array(822);
		when "0000001100110111" => data_out <= rom_array(823);
		when "0000001100111000" => data_out <= rom_array(824);
		when "0000001100111001" => data_out <= rom_array(825);
		when "0000001100111010" => data_out <= rom_array(826);
		when "0000001100111011" => data_out <= rom_array(827);
		when "0000001100111100" => data_out <= rom_array(828);
		when "0000001100111101" => data_out <= rom_array(829);
		when "0000001100111110" => data_out <= rom_array(830);
		when "0000001100111111" => data_out <= rom_array(831);
		when "0000001101000000" => data_out <= rom_array(832);
		when "0000001101000001" => data_out <= rom_array(833);
		when "0000001101000010" => data_out <= rom_array(834);
		when "0000001101000011" => data_out <= rom_array(835);
		when "0000001101000100" => data_out <= rom_array(836);
		when "0000001101000101" => data_out <= rom_array(837);
		when "0000001101000110" => data_out <= rom_array(838);
		when "0000001101000111" => data_out <= rom_array(839);
		when "0000001101001000" => data_out <= rom_array(840);
		when "0000001101001001" => data_out <= rom_array(841);
		when "0000001101001010" => data_out <= rom_array(842);
		when "0000001101001011" => data_out <= rom_array(843);
		when "0000001101001100" => data_out <= rom_array(844);
		when "0000001101001101" => data_out <= rom_array(845);
		when "0000001101001110" => data_out <= rom_array(846);
		when "0000001101001111" => data_out <= rom_array(847);
		when "0000001101010000" => data_out <= rom_array(848);
		when "0000001101010001" => data_out <= rom_array(849);
		when "0000001101010010" => data_out <= rom_array(850);
		when "0000001101010011" => data_out <= rom_array(851);
		when "0000001101010100" => data_out <= rom_array(852);
		when "0000001101010101" => data_out <= rom_array(853);
		when "0000001101010110" => data_out <= rom_array(854);
		when "0000001101010111" => data_out <= rom_array(855);
		when "0000001101011000" => data_out <= rom_array(856);
		when "0000001101011001" => data_out <= rom_array(857);
		when "0000001101011010" => data_out <= rom_array(858);
		when "0000001101011011" => data_out <= rom_array(859);
		when "0000001101011100" => data_out <= rom_array(860);
		when "0000001101011101" => data_out <= rom_array(861);
		when "0000001101011110" => data_out <= rom_array(862);
		when "0000001101011111" => data_out <= rom_array(863);
		when "0000001101100000" => data_out <= rom_array(864);
		when "0000001101100001" => data_out <= rom_array(865);
		when "0000001101100010" => data_out <= rom_array(866);
		when "0000001101100011" => data_out <= rom_array(867);
		when "0000001101100100" => data_out <= rom_array(868);
		when "0000001101100101" => data_out <= rom_array(869);
		when "0000001101100110" => data_out <= rom_array(870);
		when "0000001101100111" => data_out <= rom_array(871);
		when "0000001101101000" => data_out <= rom_array(872);
		when "0000001101101001" => data_out <= rom_array(873);
		when "0000001101101010" => data_out <= rom_array(874);
		when "0000001101101011" => data_out <= rom_array(875);
		when "0000001101101100" => data_out <= rom_array(876);
		when "0000001101101101" => data_out <= rom_array(877);
		when "0000001101101110" => data_out <= rom_array(878);
		when "0000001101101111" => data_out <= rom_array(879);
		when "0000001101110000" => data_out <= rom_array(880);
		when "0000001101110001" => data_out <= rom_array(881);
		when "0000001101110010" => data_out <= rom_array(882);
		when "0000001101110011" => data_out <= rom_array(883);
		when "0000001101110100" => data_out <= rom_array(884);
		when "0000001101110101" => data_out <= rom_array(885);
		when "0000001101110110" => data_out <= rom_array(886);
		when "0000001101110111" => data_out <= rom_array(887);
		when "0000001101111000" => data_out <= rom_array(888);
		when "0000001101111001" => data_out <= rom_array(889);
		when "0000001101111010" => data_out <= rom_array(890);
		when "0000001101111011" => data_out <= rom_array(891);
		when "0000001101111100" => data_out <= rom_array(892);
		when "0000001101111101" => data_out <= rom_array(893);
		when "0000001101111110" => data_out <= rom_array(894);
		when "0000001101111111" => data_out <= rom_array(895);
		when "0000001110000000" => data_out <= rom_array(896);
		when "0000001110000001" => data_out <= rom_array(897);
		when "0000001110000010" => data_out <= rom_array(898);
		when "0000001110000011" => data_out <= rom_array(899);
		when "0000001110000100" => data_out <= rom_array(900);
		when "0000001110000101" => data_out <= rom_array(901);
		when "0000001110000110" => data_out <= rom_array(902);
		when "0000001110000111" => data_out <= rom_array(903);
		when "0000001110001000" => data_out <= rom_array(904);
		when "0000001110001001" => data_out <= rom_array(905);
		when "0000001110001010" => data_out <= rom_array(906);
		when "0000001110001011" => data_out <= rom_array(907);
		when "0000001110001100" => data_out <= rom_array(908);
		when "0000001110001101" => data_out <= rom_array(909);
		when "0000001110001110" => data_out <= rom_array(910);
		when "0000001110001111" => data_out <= rom_array(911);
		when "0000001110010000" => data_out <= rom_array(912);
		when "0000001110010001" => data_out <= rom_array(913);
		when "0000001110010010" => data_out <= rom_array(914);
		when "0000001110010011" => data_out <= rom_array(915);
		when "0000001110010100" => data_out <= rom_array(916);
		when "0000001110010101" => data_out <= rom_array(917);
		when "0000001110010110" => data_out <= rom_array(918);
		when "0000001110010111" => data_out <= rom_array(919);
		when "0000001110011000" => data_out <= rom_array(920);
		when "0000001110011001" => data_out <= rom_array(921);
		when "0000001110011010" => data_out <= rom_array(922);
		when "0000001110011011" => data_out <= rom_array(923);
		when "0000001110011100" => data_out <= rom_array(924);
		when "0000001110011101" => data_out <= rom_array(925);
		when "0000001110011110" => data_out <= rom_array(926);
		when "0000001110011111" => data_out <= rom_array(927);
		when "0000001110100000" => data_out <= rom_array(928);
		when "0000001110100001" => data_out <= rom_array(929);
		when "0000001110100010" => data_out <= rom_array(930);
		when "0000001110100011" => data_out <= rom_array(931);
		when "0000001110100100" => data_out <= rom_array(932);
		when "0000001110100101" => data_out <= rom_array(933);
		when "0000001110100110" => data_out <= rom_array(934);
		when "0000001110100111" => data_out <= rom_array(935);
		when "0000001110101000" => data_out <= rom_array(936);
		when "0000001110101001" => data_out <= rom_array(937);
		when "0000001110101010" => data_out <= rom_array(938);
		when "0000001110101011" => data_out <= rom_array(939);
		when "0000001110101100" => data_out <= rom_array(940);
		when "0000001110101101" => data_out <= rom_array(941);
		when "0000001110101110" => data_out <= rom_array(942);
		when "0000001110101111" => data_out <= rom_array(943);
		when "0000001110110000" => data_out <= rom_array(944);
		when "0000001110110001" => data_out <= rom_array(945);
		when "0000001110110010" => data_out <= rom_array(946);
		when "0000001110110011" => data_out <= rom_array(947);
		when "0000001110110100" => data_out <= rom_array(948);
		when "0000001110110101" => data_out <= rom_array(949);
		when "0000001110110110" => data_out <= rom_array(950);
		when "0000001110110111" => data_out <= rom_array(951);
		when "0000001110111000" => data_out <= rom_array(952);
		when "0000001110111001" => data_out <= rom_array(953);
		when "0000001110111010" => data_out <= rom_array(954);
		when "0000001110111011" => data_out <= rom_array(955);
		when "0000001110111100" => data_out <= rom_array(956);
		when "0000001110111101" => data_out <= rom_array(957);
		when "0000001110111110" => data_out <= rom_array(958);
		when "0000001110111111" => data_out <= rom_array(959);
		when "0000001111000000" => data_out <= rom_array(960);
		when "0000001111000001" => data_out <= rom_array(961);
		when "0000001111000010" => data_out <= rom_array(962);
		when "0000001111000011" => data_out <= rom_array(963);
		when "0000001111000100" => data_out <= rom_array(964);
		when "0000001111000101" => data_out <= rom_array(965);
		when "0000001111000110" => data_out <= rom_array(966);
		when "0000001111000111" => data_out <= rom_array(967);
		when "0000001111001000" => data_out <= rom_array(968);
		when "0000001111001001" => data_out <= rom_array(969);
		when "0000001111001010" => data_out <= rom_array(970);
		when "0000001111001011" => data_out <= rom_array(971);
		when "0000001111001100" => data_out <= rom_array(972);
		when "0000001111001101" => data_out <= rom_array(973);
		when "0000001111001110" => data_out <= rom_array(974);
		when "0000001111001111" => data_out <= rom_array(975);
		when "0000001111010000" => data_out <= rom_array(976);
		when "0000001111010001" => data_out <= rom_array(977);
		when "0000001111010010" => data_out <= rom_array(978);
		when "0000001111010011" => data_out <= rom_array(979);
		when "0000001111010100" => data_out <= rom_array(980);
		when "0000001111010101" => data_out <= rom_array(981);
		when "0000001111010110" => data_out <= rom_array(982);
		when "0000001111010111" => data_out <= rom_array(983);
		when "0000001111011000" => data_out <= rom_array(984);
		when "0000001111011001" => data_out <= rom_array(985);
		when "0000001111011010" => data_out <= rom_array(986);
		when "0000001111011011" => data_out <= rom_array(987);
		when "0000001111011100" => data_out <= rom_array(988);
		when "0000001111011101" => data_out <= rom_array(989);
		when "0000001111011110" => data_out <= rom_array(990);
		when "0000001111011111" => data_out <= rom_array(991);
		when "0000001111100000" => data_out <= rom_array(992);
		when "0000001111100001" => data_out <= rom_array(993);
		when "0000001111100010" => data_out <= rom_array(994);
		when "0000001111100011" => data_out <= rom_array(995);
		when "0000001111100100" => data_out <= rom_array(996);
		when "0000001111100101" => data_out <= rom_array(997);
		when "0000001111100110" => data_out <= rom_array(998);
		when "0000001111100111" => data_out <= rom_array(999);
		when "0000001111101000" => data_out <= rom_array(1000);
		when "0000001111101001" => data_out <= rom_array(1001);
		when "0000001111101010" => data_out <= rom_array(1002);
		when "0000001111101011" => data_out <= rom_array(1003);
		when "0000001111101100" => data_out <= rom_array(1004);
		when "0000001111101101" => data_out <= rom_array(1005);
		when "0000001111101110" => data_out <= rom_array(1006);
		when "0000001111101111" => data_out <= rom_array(1007);
		when "0000001111110000" => data_out <= rom_array(1008);
		when "0000001111110001" => data_out <= rom_array(1009);
		when "0000001111110010" => data_out <= rom_array(1010);
		when "0000001111110011" => data_out <= rom_array(1011);
		when "0000001111110100" => data_out <= rom_array(1012);
		when "0000001111110101" => data_out <= rom_array(1013);
		when "0000001111110110" => data_out <= rom_array(1014);
		when "0000001111110111" => data_out <= rom_array(1015);
		when "0000001111111000" => data_out <= rom_array(1016);
		when "0000001111111001" => data_out <= rom_array(1017);
		when "0000001111111010" => data_out <= rom_array(1018);
		when "0000001111111011" => data_out <= rom_array(1019);
		when "0000001111111100" => data_out <= rom_array(1020);
		when "0000001111111101" => data_out <= rom_array(1021);
		when "0000001111111110" => data_out <= rom_array(1022);
		when "0000001111111111" => data_out <= rom_array(1023);
		when "0000010000000000" => data_out <= rom_array(1024);
		when "0000010000000001" => data_out <= rom_array(1025);
		when "0000010000000010" => data_out <= rom_array(1026);
		when "0000010000000011" => data_out <= rom_array(1027);
		when "0000010000000100" => data_out <= rom_array(1028);
		when "0000010000000101" => data_out <= rom_array(1029);
		when "0000010000000110" => data_out <= rom_array(1030);
		when "0000010000000111" => data_out <= rom_array(1031);
		when "0000010000001000" => data_out <= rom_array(1032);
		when "0000010000001001" => data_out <= rom_array(1033);
		when "0000010000001010" => data_out <= rom_array(1034);
		when "0000010000001011" => data_out <= rom_array(1035);
		when "0000010000001100" => data_out <= rom_array(1036);
		when "0000010000001101" => data_out <= rom_array(1037);
		when "0000010000001110" => data_out <= rom_array(1038);
		when "0000010000001111" => data_out <= rom_array(1039);
		when "0000010000010000" => data_out <= rom_array(1040);
		when "0000010000010001" => data_out <= rom_array(1041);
		when "0000010000010010" => data_out <= rom_array(1042);
		when "0000010000010011" => data_out <= rom_array(1043);
		when "0000010000010100" => data_out <= rom_array(1044);
		when "0000010000010101" => data_out <= rom_array(1045);
		when "0000010000010110" => data_out <= rom_array(1046);
		when "0000010000010111" => data_out <= rom_array(1047);
		when "0000010000011000" => data_out <= rom_array(1048);
		when "0000010000011001" => data_out <= rom_array(1049);
		when "0000010000011010" => data_out <= rom_array(1050);
		when "0000010000011011" => data_out <= rom_array(1051);
		when "0000010000011100" => data_out <= rom_array(1052);
		when "0000010000011101" => data_out <= rom_array(1053);
		when "0000010000011110" => data_out <= rom_array(1054);
		when "0000010000011111" => data_out <= rom_array(1055);
		when "0000010000100000" => data_out <= rom_array(1056);
		when "0000010000100001" => data_out <= rom_array(1057);
		when "0000010000100010" => data_out <= rom_array(1058);
		when "0000010000100011" => data_out <= rom_array(1059);
		when "0000010000100100" => data_out <= rom_array(1060);
		when "0000010000100101" => data_out <= rom_array(1061);
		when "0000010000100110" => data_out <= rom_array(1062);
		when "0000010000100111" => data_out <= rom_array(1063);
		when "0000010000101000" => data_out <= rom_array(1064);
		when "0000010000101001" => data_out <= rom_array(1065);
		when "0000010000101010" => data_out <= rom_array(1066);
		when "0000010000101011" => data_out <= rom_array(1067);
		when "0000010000101100" => data_out <= rom_array(1068);
		when "0000010000101101" => data_out <= rom_array(1069);
		when "0000010000101110" => data_out <= rom_array(1070);
		when "0000010000101111" => data_out <= rom_array(1071);
		when "0000010000110000" => data_out <= rom_array(1072);
		when "0000010000110001" => data_out <= rom_array(1073);
		when "0000010000110010" => data_out <= rom_array(1074);
		when "0000010000110011" => data_out <= rom_array(1075);
		when "0000010000110100" => data_out <= rom_array(1076);
		when "0000010000110101" => data_out <= rom_array(1077);
		when "0000010000110110" => data_out <= rom_array(1078);
		when "0000010000110111" => data_out <= rom_array(1079);
		when "0000010000111000" => data_out <= rom_array(1080);
		when "0000010000111001" => data_out <= rom_array(1081);
		when "0000010000111010" => data_out <= rom_array(1082);
		when "0000010000111011" => data_out <= rom_array(1083);
		when "0000010000111100" => data_out <= rom_array(1084);
		when "0000010000111101" => data_out <= rom_array(1085);
		when "0000010000111110" => data_out <= rom_array(1086);
		when "0000010000111111" => data_out <= rom_array(1087);
		when "0000010001000000" => data_out <= rom_array(1088);
		when "0000010001000001" => data_out <= rom_array(1089);
		when "0000010001000010" => data_out <= rom_array(1090);
		when "0000010001000011" => data_out <= rom_array(1091);
		when "0000010001000100" => data_out <= rom_array(1092);
		when "0000010001000101" => data_out <= rom_array(1093);
		when "0000010001000110" => data_out <= rom_array(1094);
		when "0000010001000111" => data_out <= rom_array(1095);
		when "0000010001001000" => data_out <= rom_array(1096);
		when "0000010001001001" => data_out <= rom_array(1097);
		when "0000010001001010" => data_out <= rom_array(1098);
		when "0000010001001011" => data_out <= rom_array(1099);
		when "0000010001001100" => data_out <= rom_array(1100);
		when "0000010001001101" => data_out <= rom_array(1101);
		when "0000010001001110" => data_out <= rom_array(1102);
		when "0000010001001111" => data_out <= rom_array(1103);
		when "0000010001010000" => data_out <= rom_array(1104);
		when "0000010001010001" => data_out <= rom_array(1105);
		when "0000010001010010" => data_out <= rom_array(1106);
		when "0000010001010011" => data_out <= rom_array(1107);
		when "0000010001010100" => data_out <= rom_array(1108);
		when "0000010001010101" => data_out <= rom_array(1109);
		when "0000010001010110" => data_out <= rom_array(1110);
		when "0000010001010111" => data_out <= rom_array(1111);
		when "0000010001011000" => data_out <= rom_array(1112);
		when "0000010001011001" => data_out <= rom_array(1113);
		when "0000010001011010" => data_out <= rom_array(1114);
		when "0000010001011011" => data_out <= rom_array(1115);
		when "0000010001011100" => data_out <= rom_array(1116);
		when "0000010001011101" => data_out <= rom_array(1117);
		when "0000010001011110" => data_out <= rom_array(1118);
		when "0000010001011111" => data_out <= rom_array(1119);
		when "0000010001100000" => data_out <= rom_array(1120);
		when "0000010001100001" => data_out <= rom_array(1121);
		when "0000010001100010" => data_out <= rom_array(1122);
		when "0000010001100011" => data_out <= rom_array(1123);
		when "0000010001100100" => data_out <= rom_array(1124);
		when "0000010001100101" => data_out <= rom_array(1125);
		when "0000010001100110" => data_out <= rom_array(1126);
		when "0000010001100111" => data_out <= rom_array(1127);
		when "0000010001101000" => data_out <= rom_array(1128);
		when "0000010001101001" => data_out <= rom_array(1129);
		when "0000010001101010" => data_out <= rom_array(1130);
		when "0000010001101011" => data_out <= rom_array(1131);
		when "0000010001101100" => data_out <= rom_array(1132);
		when "0000010001101101" => data_out <= rom_array(1133);
		when "0000010001101110" => data_out <= rom_array(1134);
		when "0000010001101111" => data_out <= rom_array(1135);
		when "0000010001110000" => data_out <= rom_array(1136);
		when "0000010001110001" => data_out <= rom_array(1137);
		when "0000010001110010" => data_out <= rom_array(1138);
		when "0000010001110011" => data_out <= rom_array(1139);
		when "0000010001110100" => data_out <= rom_array(1140);
		when "0000010001110101" => data_out <= rom_array(1141);
		when "0000010001110110" => data_out <= rom_array(1142);
		when "0000010001110111" => data_out <= rom_array(1143);
		when "0000010001111000" => data_out <= rom_array(1144);
		when "0000010001111001" => data_out <= rom_array(1145);
		when "0000010001111010" => data_out <= rom_array(1146);
		when "0000010001111011" => data_out <= rom_array(1147);
		when "0000010001111100" => data_out <= rom_array(1148);
		when "0000010001111101" => data_out <= rom_array(1149);
		when "0000010001111110" => data_out <= rom_array(1150);
		when "0000010001111111" => data_out <= rom_array(1151);
		when "0000010010000000" => data_out <= rom_array(1152);
		when "0000010010000001" => data_out <= rom_array(1153);
		when "0000010010000010" => data_out <= rom_array(1154);
		when "0000010010000011" => data_out <= rom_array(1155);
		when "0000010010000100" => data_out <= rom_array(1156);
		when "0000010010000101" => data_out <= rom_array(1157);
		when "0000010010000110" => data_out <= rom_array(1158);
		when "0000010010000111" => data_out <= rom_array(1159);
		when "0000010010001000" => data_out <= rom_array(1160);
		when "0000010010001001" => data_out <= rom_array(1161);
		when "0000010010001010" => data_out <= rom_array(1162);
		when "0000010010001011" => data_out <= rom_array(1163);
		when "0000010010001100" => data_out <= rom_array(1164);
		when "0000010010001101" => data_out <= rom_array(1165);
		when "0000010010001110" => data_out <= rom_array(1166);
		when "0000010010001111" => data_out <= rom_array(1167);
		when "0000010010010000" => data_out <= rom_array(1168);
		when "0000010010010001" => data_out <= rom_array(1169);
		when "0000010010010010" => data_out <= rom_array(1170);
		when "0000010010010011" => data_out <= rom_array(1171);
		when "0000010010010100" => data_out <= rom_array(1172);
		when "0000010010010101" => data_out <= rom_array(1173);
		when "0000010010010110" => data_out <= rom_array(1174);
		when "0000010010010111" => data_out <= rom_array(1175);
		when "0000010010011000" => data_out <= rom_array(1176);
		when "0000010010011001" => data_out <= rom_array(1177);
		when "0000010010011010" => data_out <= rom_array(1178);
		when "0000010010011011" => data_out <= rom_array(1179);
		when "0000010010011100" => data_out <= rom_array(1180);
		when "0000010010011101" => data_out <= rom_array(1181);
		when "0000010010011110" => data_out <= rom_array(1182);
		when "0000010010011111" => data_out <= rom_array(1183);
		when "0000010010100000" => data_out <= rom_array(1184);
		when "0000010010100001" => data_out <= rom_array(1185);
		when "0000010010100010" => data_out <= rom_array(1186);
		when "0000010010100011" => data_out <= rom_array(1187);
		when "0000010010100100" => data_out <= rom_array(1188);
		when "0000010010100101" => data_out <= rom_array(1189);
		when "0000010010100110" => data_out <= rom_array(1190);
		when "0000010010100111" => data_out <= rom_array(1191);
		when "0000010010101000" => data_out <= rom_array(1192);
		when "0000010010101001" => data_out <= rom_array(1193);
		when "0000010010101010" => data_out <= rom_array(1194);
		when "0000010010101011" => data_out <= rom_array(1195);
		when "0000010010101100" => data_out <= rom_array(1196);
		when "0000010010101101" => data_out <= rom_array(1197);
		when "0000010010101110" => data_out <= rom_array(1198);
		when "0000010010101111" => data_out <= rom_array(1199);
		when "0000010010110000" => data_out <= rom_array(1200);
		when "0000010010110001" => data_out <= rom_array(1201);
		when "0000010010110010" => data_out <= rom_array(1202);
		when "0000010010110011" => data_out <= rom_array(1203);
		when "0000010010110100" => data_out <= rom_array(1204);
		when "0000010010110101" => data_out <= rom_array(1205);
		when "0000010010110110" => data_out <= rom_array(1206);
		when "0000010010110111" => data_out <= rom_array(1207);
		when "0000010010111000" => data_out <= rom_array(1208);
		when "0000010010111001" => data_out <= rom_array(1209);
		when "0000010010111010" => data_out <= rom_array(1210);
		when "0000010010111011" => data_out <= rom_array(1211);
		when "0000010010111100" => data_out <= rom_array(1212);
		when "0000010010111101" => data_out <= rom_array(1213);
		when "0000010010111110" => data_out <= rom_array(1214);
		when "0000010010111111" => data_out <= rom_array(1215);
		when "0000010011000000" => data_out <= rom_array(1216);
		when "0000010011000001" => data_out <= rom_array(1217);
		when "0000010011000010" => data_out <= rom_array(1218);
		when "0000010011000011" => data_out <= rom_array(1219);
		when "0000010011000100" => data_out <= rom_array(1220);
		when "0000010011000101" => data_out <= rom_array(1221);
		when "0000010011000110" => data_out <= rom_array(1222);
		when "0000010011000111" => data_out <= rom_array(1223);
		when "0000010011001000" => data_out <= rom_array(1224);
		when "0000010011001001" => data_out <= rom_array(1225);
		when "0000010011001010" => data_out <= rom_array(1226);
		when "0000010011001011" => data_out <= rom_array(1227);
		when "0000010011001100" => data_out <= rom_array(1228);
		when "0000010011001101" => data_out <= rom_array(1229);
		when "0000010011001110" => data_out <= rom_array(1230);
		when "0000010011001111" => data_out <= rom_array(1231);
		when "0000010011010000" => data_out <= rom_array(1232);
		when "0000010011010001" => data_out <= rom_array(1233);
		when "0000010011010010" => data_out <= rom_array(1234);
		when "0000010011010011" => data_out <= rom_array(1235);
		when "0000010011010100" => data_out <= rom_array(1236);
		when "0000010011010101" => data_out <= rom_array(1237);
		when "0000010011010110" => data_out <= rom_array(1238);
		when "0000010011010111" => data_out <= rom_array(1239);
		when "0000010011011000" => data_out <= rom_array(1240);
		when "0000010011011001" => data_out <= rom_array(1241);
		when "0000010011011010" => data_out <= rom_array(1242);
		when "0000010011011011" => data_out <= rom_array(1243);
		when "0000010011011100" => data_out <= rom_array(1244);
		when "0000010011011101" => data_out <= rom_array(1245);
		when "0000010011011110" => data_out <= rom_array(1246);
		when "0000010011011111" => data_out <= rom_array(1247);
		when "0000010011100000" => data_out <= rom_array(1248);
		when "0000010011100001" => data_out <= rom_array(1249);
		when "0000010011100010" => data_out <= rom_array(1250);
		when "0000010011100011" => data_out <= rom_array(1251);
		when "0000010011100100" => data_out <= rom_array(1252);
		when "0000010011100101" => data_out <= rom_array(1253);
		when "0000010011100110" => data_out <= rom_array(1254);
		when "0000010011100111" => data_out <= rom_array(1255);
		when "0000010011101000" => data_out <= rom_array(1256);
		when "0000010011101001" => data_out <= rom_array(1257);
		when "0000010011101010" => data_out <= rom_array(1258);
		when "0000010011101011" => data_out <= rom_array(1259);
		when "0000010011101100" => data_out <= rom_array(1260);
		when "0000010011101101" => data_out <= rom_array(1261);
		when "0000010011101110" => data_out <= rom_array(1262);
		when "0000010011101111" => data_out <= rom_array(1263);
		when "0000010011110000" => data_out <= rom_array(1264);
		when "0000010011110001" => data_out <= rom_array(1265);
		when "0000010011110010" => data_out <= rom_array(1266);
		when "0000010011110011" => data_out <= rom_array(1267);
		when "0000010011110100" => data_out <= rom_array(1268);
		when "0000010011110101" => data_out <= rom_array(1269);
		when "0000010011110110" => data_out <= rom_array(1270);
		when "0000010011110111" => data_out <= rom_array(1271);
		when "0000010011111000" => data_out <= rom_array(1272);
		when "0000010011111001" => data_out <= rom_array(1273);
		when "0000010011111010" => data_out <= rom_array(1274);
		when "0000010011111011" => data_out <= rom_array(1275);
		when "0000010011111100" => data_out <= rom_array(1276);
		when "0000010011111101" => data_out <= rom_array(1277);
		when "0000010011111110" => data_out <= rom_array(1278);
		when "0000010011111111" => data_out <= rom_array(1279);
		when "0000010100000000" => data_out <= rom_array(1280);
		when "0000010100000001" => data_out <= rom_array(1281);
		when "0000010100000010" => data_out <= rom_array(1282);
		when "0000010100000011" => data_out <= rom_array(1283);
		when "0000010100000100" => data_out <= rom_array(1284);
		when "0000010100000101" => data_out <= rom_array(1285);
		when "0000010100000110" => data_out <= rom_array(1286);
		when "0000010100000111" => data_out <= rom_array(1287);
		when "0000010100001000" => data_out <= rom_array(1288);
		when "0000010100001001" => data_out <= rom_array(1289);
		when "0000010100001010" => data_out <= rom_array(1290);
		when "0000010100001011" => data_out <= rom_array(1291);
		when "0000010100001100" => data_out <= rom_array(1292);
		when "0000010100001101" => data_out <= rom_array(1293);
		when "0000010100001110" => data_out <= rom_array(1294);
		when "0000010100001111" => data_out <= rom_array(1295);
		when "0000010100010000" => data_out <= rom_array(1296);
		when "0000010100010001" => data_out <= rom_array(1297);
		when "0000010100010010" => data_out <= rom_array(1298);
		when "0000010100010011" => data_out <= rom_array(1299);
		when "0000010100010100" => data_out <= rom_array(1300);
		when "0000010100010101" => data_out <= rom_array(1301);
		when "0000010100010110" => data_out <= rom_array(1302);
		when "0000010100010111" => data_out <= rom_array(1303);
		when "0000010100011000" => data_out <= rom_array(1304);
		when "0000010100011001" => data_out <= rom_array(1305);
		when "0000010100011010" => data_out <= rom_array(1306);
		when "0000010100011011" => data_out <= rom_array(1307);
		when "0000010100011100" => data_out <= rom_array(1308);
		when "0000010100011101" => data_out <= rom_array(1309);
		when "0000010100011110" => data_out <= rom_array(1310);
		when "0000010100011111" => data_out <= rom_array(1311);
		when "0000010100100000" => data_out <= rom_array(1312);
		when "0000010100100001" => data_out <= rom_array(1313);
		when "0000010100100010" => data_out <= rom_array(1314);
		when "0000010100100011" => data_out <= rom_array(1315);
		when "0000010100100100" => data_out <= rom_array(1316);
		when "0000010100100101" => data_out <= rom_array(1317);
		when "0000010100100110" => data_out <= rom_array(1318);
		when "0000010100100111" => data_out <= rom_array(1319);
		when "0000010100101000" => data_out <= rom_array(1320);
		when "0000010100101001" => data_out <= rom_array(1321);
		when "0000010100101010" => data_out <= rom_array(1322);
		when "0000010100101011" => data_out <= rom_array(1323);
		when "0000010100101100" => data_out <= rom_array(1324);
		when "0000010100101101" => data_out <= rom_array(1325);
		when "0000010100101110" => data_out <= rom_array(1326);
		when "0000010100101111" => data_out <= rom_array(1327);
		when "0000010100110000" => data_out <= rom_array(1328);
		when "0000010100110001" => data_out <= rom_array(1329);
		when "0000010100110010" => data_out <= rom_array(1330);
		when "0000010100110011" => data_out <= rom_array(1331);
		when "0000010100110100" => data_out <= rom_array(1332);
		when "0000010100110101" => data_out <= rom_array(1333);
		when "0000010100110110" => data_out <= rom_array(1334);
		when "0000010100110111" => data_out <= rom_array(1335);
		when "0000010100111000" => data_out <= rom_array(1336);
		when "0000010100111001" => data_out <= rom_array(1337);
		when "0000010100111010" => data_out <= rom_array(1338);
		when "0000010100111011" => data_out <= rom_array(1339);
		when "0000010100111100" => data_out <= rom_array(1340);
		when "0000010100111101" => data_out <= rom_array(1341);
		when "0000010100111110" => data_out <= rom_array(1342);
		when "0000010100111111" => data_out <= rom_array(1343);
		when "0000010101000000" => data_out <= rom_array(1344);
		when "0000010101000001" => data_out <= rom_array(1345);
		when "0000010101000010" => data_out <= rom_array(1346);
		when "0000010101000011" => data_out <= rom_array(1347);
		when "0000010101000100" => data_out <= rom_array(1348);
		when "0000010101000101" => data_out <= rom_array(1349);
		when "0000010101000110" => data_out <= rom_array(1350);
		when "0000010101000111" => data_out <= rom_array(1351);
		when "0000010101001000" => data_out <= rom_array(1352);
		when "0000010101001001" => data_out <= rom_array(1353);
		when "0000010101001010" => data_out <= rom_array(1354);
		when "0000010101001011" => data_out <= rom_array(1355);
		when "0000010101001100" => data_out <= rom_array(1356);
		when "0000010101001101" => data_out <= rom_array(1357);
		when "0000010101001110" => data_out <= rom_array(1358);
		when "0000010101001111" => data_out <= rom_array(1359);
		when "0000010101010000" => data_out <= rom_array(1360);
		when "0000010101010001" => data_out <= rom_array(1361);
		when "0000010101010010" => data_out <= rom_array(1362);
		when "0000010101010011" => data_out <= rom_array(1363);
		when "0000010101010100" => data_out <= rom_array(1364);
		when "0000010101010101" => data_out <= rom_array(1365);
		when "0000010101010110" => data_out <= rom_array(1366);
		when "0000010101010111" => data_out <= rom_array(1367);
		when "0000010101011000" => data_out <= rom_array(1368);
		when "0000010101011001" => data_out <= rom_array(1369);
		when "0000010101011010" => data_out <= rom_array(1370);
		when "0000010101011011" => data_out <= rom_array(1371);
		when "0000010101011100" => data_out <= rom_array(1372);
		when "0000010101011101" => data_out <= rom_array(1373);
		when "0000010101011110" => data_out <= rom_array(1374);
		when "0000010101011111" => data_out <= rom_array(1375);
		when "0000010101100000" => data_out <= rom_array(1376);
		when "0000010101100001" => data_out <= rom_array(1377);
		when "0000010101100010" => data_out <= rom_array(1378);
		when "0000010101100011" => data_out <= rom_array(1379);
		when "0000010101100100" => data_out <= rom_array(1380);
		when "0000010101100101" => data_out <= rom_array(1381);
		when "0000010101100110" => data_out <= rom_array(1382);
		when "0000010101100111" => data_out <= rom_array(1383);
		when "0000010101101000" => data_out <= rom_array(1384);
		when "0000010101101001" => data_out <= rom_array(1385);
		when "0000010101101010" => data_out <= rom_array(1386);
		when "0000010101101011" => data_out <= rom_array(1387);
		when "0000010101101100" => data_out <= rom_array(1388);
		when "0000010101101101" => data_out <= rom_array(1389);
		when "0000010101101110" => data_out <= rom_array(1390);
		when "0000010101101111" => data_out <= rom_array(1391);
		when "0000010101110000" => data_out <= rom_array(1392);
		when "0000010101110001" => data_out <= rom_array(1393);
		when "0000010101110010" => data_out <= rom_array(1394);
		when "0000010101110011" => data_out <= rom_array(1395);
		when "0000010101110100" => data_out <= rom_array(1396);
		when "0000010101110101" => data_out <= rom_array(1397);
		when "0000010101110110" => data_out <= rom_array(1398);
		when "0000010101110111" => data_out <= rom_array(1399);
		when "0000010101111000" => data_out <= rom_array(1400);
		when "0000010101111001" => data_out <= rom_array(1401);
		when "0000010101111010" => data_out <= rom_array(1402);
		when "0000010101111011" => data_out <= rom_array(1403);
		when "0000010101111100" => data_out <= rom_array(1404);
		when "0000010101111101" => data_out <= rom_array(1405);
		when "0000010101111110" => data_out <= rom_array(1406);
		when "0000010101111111" => data_out <= rom_array(1407);
		when "0000010110000000" => data_out <= rom_array(1408);
		when "0000010110000001" => data_out <= rom_array(1409);
		when "0000010110000010" => data_out <= rom_array(1410);
		when "0000010110000011" => data_out <= rom_array(1411);
		when "0000010110000100" => data_out <= rom_array(1412);
		when "0000010110000101" => data_out <= rom_array(1413);
		when "0000010110000110" => data_out <= rom_array(1414);
		when "0000010110000111" => data_out <= rom_array(1415);
		when "0000010110001000" => data_out <= rom_array(1416);
		when "0000010110001001" => data_out <= rom_array(1417);
		when "0000010110001010" => data_out <= rom_array(1418);
		when "0000010110001011" => data_out <= rom_array(1419);
		when "0000010110001100" => data_out <= rom_array(1420);
		when "0000010110001101" => data_out <= rom_array(1421);
		when "0000010110001110" => data_out <= rom_array(1422);
		when "0000010110001111" => data_out <= rom_array(1423);
		when "0000010110010000" => data_out <= rom_array(1424);
		when "0000010110010001" => data_out <= rom_array(1425);
		when "0000010110010010" => data_out <= rom_array(1426);
		when "0000010110010011" => data_out <= rom_array(1427);
		when "0000010110010100" => data_out <= rom_array(1428);
		when "0000010110010101" => data_out <= rom_array(1429);
		when "0000010110010110" => data_out <= rom_array(1430);
		when "0000010110010111" => data_out <= rom_array(1431);
		when "0000010110011000" => data_out <= rom_array(1432);
		when "0000010110011001" => data_out <= rom_array(1433);
		when "0000010110011010" => data_out <= rom_array(1434);
		when "0000010110011011" => data_out <= rom_array(1435);
		when "0000010110011100" => data_out <= rom_array(1436);
		when "0000010110011101" => data_out <= rom_array(1437);
		when "0000010110011110" => data_out <= rom_array(1438);
		when "0000010110011111" => data_out <= rom_array(1439);
		when "0000010110100000" => data_out <= rom_array(1440);
		when "0000010110100001" => data_out <= rom_array(1441);
		when "0000010110100010" => data_out <= rom_array(1442);
		when "0000010110100011" => data_out <= rom_array(1443);
		when "0000010110100100" => data_out <= rom_array(1444);
		when "0000010110100101" => data_out <= rom_array(1445);
		when "0000010110100110" => data_out <= rom_array(1446);
		when "0000010110100111" => data_out <= rom_array(1447);
		when "0000010110101000" => data_out <= rom_array(1448);
		when "0000010110101001" => data_out <= rom_array(1449);
		when "0000010110101010" => data_out <= rom_array(1450);
		when "0000010110101011" => data_out <= rom_array(1451);
		when "0000010110101100" => data_out <= rom_array(1452);
		when "0000010110101101" => data_out <= rom_array(1453);
		when "0000010110101110" => data_out <= rom_array(1454);
		when "0000010110101111" => data_out <= rom_array(1455);
		when "0000010110110000" => data_out <= rom_array(1456);
		when "0000010110110001" => data_out <= rom_array(1457);
		when "0000010110110010" => data_out <= rom_array(1458);
		when "0000010110110011" => data_out <= rom_array(1459);
		when "0000010110110100" => data_out <= rom_array(1460);
		when "0000010110110101" => data_out <= rom_array(1461);
		when "0000010110110110" => data_out <= rom_array(1462);
		when "0000010110110111" => data_out <= rom_array(1463);
		when "0000010110111000" => data_out <= rom_array(1464);
		when "0000010110111001" => data_out <= rom_array(1465);
		when "0000010110111010" => data_out <= rom_array(1466);
		when "0000010110111011" => data_out <= rom_array(1467);
		when "0000010110111100" => data_out <= rom_array(1468);
		when "0000010110111101" => data_out <= rom_array(1469);
		when "0000010110111110" => data_out <= rom_array(1470);
		when "0000010110111111" => data_out <= rom_array(1471);
		when "0000010111000000" => data_out <= rom_array(1472);
		when "0000010111000001" => data_out <= rom_array(1473);
		when "0000010111000010" => data_out <= rom_array(1474);
		when "0000010111000011" => data_out <= rom_array(1475);
		when "0000010111000100" => data_out <= rom_array(1476);
		when "0000010111000101" => data_out <= rom_array(1477);
		when "0000010111000110" => data_out <= rom_array(1478);
		when "0000010111000111" => data_out <= rom_array(1479);
		when "0000010111001000" => data_out <= rom_array(1480);
		when "0000010111001001" => data_out <= rom_array(1481);
		when "0000010111001010" => data_out <= rom_array(1482);
		when "0000010111001011" => data_out <= rom_array(1483);
		when "0000010111001100" => data_out <= rom_array(1484);
		when "0000010111001101" => data_out <= rom_array(1485);
		when "0000010111001110" => data_out <= rom_array(1486);
		when "0000010111001111" => data_out <= rom_array(1487);
		when "0000010111010000" => data_out <= rom_array(1488);
		when "0000010111010001" => data_out <= rom_array(1489);
		when "0000010111010010" => data_out <= rom_array(1490);
		when "0000010111010011" => data_out <= rom_array(1491);
		when "0000010111010100" => data_out <= rom_array(1492);
		when "0000010111010101" => data_out <= rom_array(1493);
		when "0000010111010110" => data_out <= rom_array(1494);
		when "0000010111010111" => data_out <= rom_array(1495);
		when "0000010111011000" => data_out <= rom_array(1496);
		when "0000010111011001" => data_out <= rom_array(1497);
		when "0000010111011010" => data_out <= rom_array(1498);
		when "0000010111011011" => data_out <= rom_array(1499);
		when "0000010111011100" => data_out <= rom_array(1500);
		when "0000010111011101" => data_out <= rom_array(1501);
		when "0000010111011110" => data_out <= rom_array(1502);
		when "0000010111011111" => data_out <= rom_array(1503);
		when "0000010111100000" => data_out <= rom_array(1504);
		when "0000010111100001" => data_out <= rom_array(1505);
		when "0000010111100010" => data_out <= rom_array(1506);
		when "0000010111100011" => data_out <= rom_array(1507);
		when "0000010111100100" => data_out <= rom_array(1508);
		when "0000010111100101" => data_out <= rom_array(1509);
		when "0000010111100110" => data_out <= rom_array(1510);
		when "0000010111100111" => data_out <= rom_array(1511);
		when "0000010111101000" => data_out <= rom_array(1512);
		when "0000010111101001" => data_out <= rom_array(1513);
		when "0000010111101010" => data_out <= rom_array(1514);
		when "0000010111101011" => data_out <= rom_array(1515);
		when "0000010111101100" => data_out <= rom_array(1516);
		when "0000010111101101" => data_out <= rom_array(1517);
		when "0000010111101110" => data_out <= rom_array(1518);
		when "0000010111101111" => data_out <= rom_array(1519);
		when "0000010111110000" => data_out <= rom_array(1520);
		when "0000010111110001" => data_out <= rom_array(1521);
		when "0000010111110010" => data_out <= rom_array(1522);
		when "0000010111110011" => data_out <= rom_array(1523);
		when "0000010111110100" => data_out <= rom_array(1524);
		when "0000010111110101" => data_out <= rom_array(1525);
		when "0000010111110110" => data_out <= rom_array(1526);
		when "0000010111110111" => data_out <= rom_array(1527);
		when "0000010111111000" => data_out <= rom_array(1528);
		when "0000010111111001" => data_out <= rom_array(1529);
		when "0000010111111010" => data_out <= rom_array(1530);
		when "0000010111111011" => data_out <= rom_array(1531);
		when "0000010111111100" => data_out <= rom_array(1532);
		when "0000010111111101" => data_out <= rom_array(1533);
		when "0000010111111110" => data_out <= rom_array(1534);
		when "0000010111111111" => data_out <= rom_array(1535);
		when "0000011000000000" => data_out <= rom_array(1536);
		when "0000011000000001" => data_out <= rom_array(1537);
		when "0000011000000010" => data_out <= rom_array(1538);
		when "0000011000000011" => data_out <= rom_array(1539);
		when "0000011000000100" => data_out <= rom_array(1540);
		when "0000011000000101" => data_out <= rom_array(1541);
		when "0000011000000110" => data_out <= rom_array(1542);
		when "0000011000000111" => data_out <= rom_array(1543);
		when "0000011000001000" => data_out <= rom_array(1544);
		when "0000011000001001" => data_out <= rom_array(1545);
		when "0000011000001010" => data_out <= rom_array(1546);
		when "0000011000001011" => data_out <= rom_array(1547);
		when "0000011000001100" => data_out <= rom_array(1548);
		when "0000011000001101" => data_out <= rom_array(1549);
		when "0000011000001110" => data_out <= rom_array(1550);
		when "0000011000001111" => data_out <= rom_array(1551);
		when "0000011000010000" => data_out <= rom_array(1552);
		when "0000011000010001" => data_out <= rom_array(1553);
		when "0000011000010010" => data_out <= rom_array(1554);
		when "0000011000010011" => data_out <= rom_array(1555);
		when "0000011000010100" => data_out <= rom_array(1556);
		when "0000011000010101" => data_out <= rom_array(1557);
		when "0000011000010110" => data_out <= rom_array(1558);
		when "0000011000010111" => data_out <= rom_array(1559);
		when "0000011000011000" => data_out <= rom_array(1560);
		when "0000011000011001" => data_out <= rom_array(1561);
		when "0000011000011010" => data_out <= rom_array(1562);
		when "0000011000011011" => data_out <= rom_array(1563);
		when "0000011000011100" => data_out <= rom_array(1564);
		when "0000011000011101" => data_out <= rom_array(1565);
		when "0000011000011110" => data_out <= rom_array(1566);
		when "0000011000011111" => data_out <= rom_array(1567);
		when "0000011000100000" => data_out <= rom_array(1568);
		when "0000011000100001" => data_out <= rom_array(1569);
		when "0000011000100010" => data_out <= rom_array(1570);
		when "0000011000100011" => data_out <= rom_array(1571);
		when "0000011000100100" => data_out <= rom_array(1572);
		when "0000011000100101" => data_out <= rom_array(1573);
		when "0000011000100110" => data_out <= rom_array(1574);
		when "0000011000100111" => data_out <= rom_array(1575);
		when "0000011000101000" => data_out <= rom_array(1576);
		when "0000011000101001" => data_out <= rom_array(1577);
		when "0000011000101010" => data_out <= rom_array(1578);
		when "0000011000101011" => data_out <= rom_array(1579);
		when "0000011000101100" => data_out <= rom_array(1580);
		when "0000011000101101" => data_out <= rom_array(1581);
		when "0000011000101110" => data_out <= rom_array(1582);
		when "0000011000101111" => data_out <= rom_array(1583);
		when "0000011000110000" => data_out <= rom_array(1584);
		when "0000011000110001" => data_out <= rom_array(1585);
		when "0000011000110010" => data_out <= rom_array(1586);
		when "0000011000110011" => data_out <= rom_array(1587);
		when "0000011000110100" => data_out <= rom_array(1588);
		when "0000011000110101" => data_out <= rom_array(1589);
		when "0000011000110110" => data_out <= rom_array(1590);
		when "0000011000110111" => data_out <= rom_array(1591);
		when "0000011000111000" => data_out <= rom_array(1592);
		when "0000011000111001" => data_out <= rom_array(1593);
		when "0000011000111010" => data_out <= rom_array(1594);
		when "0000011000111011" => data_out <= rom_array(1595);
		when "0000011000111100" => data_out <= rom_array(1596);
		when "0000011000111101" => data_out <= rom_array(1597);
		when "0000011000111110" => data_out <= rom_array(1598);
		when "0000011000111111" => data_out <= rom_array(1599);
		when "0000011001000000" => data_out <= rom_array(1600);
		when "0000011001000001" => data_out <= rom_array(1601);
		when "0000011001000010" => data_out <= rom_array(1602);
		when "0000011001000011" => data_out <= rom_array(1603);
		when "0000011001000100" => data_out <= rom_array(1604);
		when "0000011001000101" => data_out <= rom_array(1605);
		when "0000011001000110" => data_out <= rom_array(1606);
		when "0000011001000111" => data_out <= rom_array(1607);
		when "0000011001001000" => data_out <= rom_array(1608);
		when "0000011001001001" => data_out <= rom_array(1609);
		when "0000011001001010" => data_out <= rom_array(1610);
		when "0000011001001011" => data_out <= rom_array(1611);
		when "0000011001001100" => data_out <= rom_array(1612);
		when "0000011001001101" => data_out <= rom_array(1613);
		when "0000011001001110" => data_out <= rom_array(1614);
		when "0000011001001111" => data_out <= rom_array(1615);
		when "0000011001010000" => data_out <= rom_array(1616);
		when "0000011001010001" => data_out <= rom_array(1617);
		when "0000011001010010" => data_out <= rom_array(1618);
		when "0000011001010011" => data_out <= rom_array(1619);
		when "0000011001010100" => data_out <= rom_array(1620);
		when "0000011001010101" => data_out <= rom_array(1621);
		when "0000011001010110" => data_out <= rom_array(1622);
		when "0000011001010111" => data_out <= rom_array(1623);
		when "0000011001011000" => data_out <= rom_array(1624);
		when "0000011001011001" => data_out <= rom_array(1625);
		when "0000011001011010" => data_out <= rom_array(1626);
		when "0000011001011011" => data_out <= rom_array(1627);
		when "0000011001011100" => data_out <= rom_array(1628);
		when "0000011001011101" => data_out <= rom_array(1629);
		when "0000011001011110" => data_out <= rom_array(1630);
		when "0000011001011111" => data_out <= rom_array(1631);
		when "0000011001100000" => data_out <= rom_array(1632);
		when "0000011001100001" => data_out <= rom_array(1633);
		when "0000011001100010" => data_out <= rom_array(1634);
		when "0000011001100011" => data_out <= rom_array(1635);
		when "0000011001100100" => data_out <= rom_array(1636);
		when "0000011001100101" => data_out <= rom_array(1637);
		when "0000011001100110" => data_out <= rom_array(1638);
		when "0000011001100111" => data_out <= rom_array(1639);
		when "0000011001101000" => data_out <= rom_array(1640);
		when "0000011001101001" => data_out <= rom_array(1641);
		when "0000011001101010" => data_out <= rom_array(1642);
		when "0000011001101011" => data_out <= rom_array(1643);
		when "0000011001101100" => data_out <= rom_array(1644);
		when "0000011001101101" => data_out <= rom_array(1645);
		when "0000011001101110" => data_out <= rom_array(1646);
		when "0000011001101111" => data_out <= rom_array(1647);
		when "0000011001110000" => data_out <= rom_array(1648);
		when "0000011001110001" => data_out <= rom_array(1649);
		when "0000011001110010" => data_out <= rom_array(1650);
		when "0000011001110011" => data_out <= rom_array(1651);
		when "0000011001110100" => data_out <= rom_array(1652);
		when "0000011001110101" => data_out <= rom_array(1653);
		when "0000011001110110" => data_out <= rom_array(1654);
		when "0000011001110111" => data_out <= rom_array(1655);
		when "0000011001111000" => data_out <= rom_array(1656);
		when "0000011001111001" => data_out <= rom_array(1657);
		when "0000011001111010" => data_out <= rom_array(1658);
		when "0000011001111011" => data_out <= rom_array(1659);
		when "0000011001111100" => data_out <= rom_array(1660);
		when "0000011001111101" => data_out <= rom_array(1661);
		when "0000011001111110" => data_out <= rom_array(1662);
		when "0000011001111111" => data_out <= rom_array(1663);
		when "0000011010000000" => data_out <= rom_array(1664);
		when "0000011010000001" => data_out <= rom_array(1665);
		when "0000011010000010" => data_out <= rom_array(1666);
		when "0000011010000011" => data_out <= rom_array(1667);
		when "0000011010000100" => data_out <= rom_array(1668);
		when "0000011010000101" => data_out <= rom_array(1669);
		when "0000011010000110" => data_out <= rom_array(1670);
		when "0000011010000111" => data_out <= rom_array(1671);
		when "0000011010001000" => data_out <= rom_array(1672);
		when "0000011010001001" => data_out <= rom_array(1673);
		when "0000011010001010" => data_out <= rom_array(1674);
		when "0000011010001011" => data_out <= rom_array(1675);
		when "0000011010001100" => data_out <= rom_array(1676);
		when "0000011010001101" => data_out <= rom_array(1677);
		when "0000011010001110" => data_out <= rom_array(1678);
		when "0000011010001111" => data_out <= rom_array(1679);
		when "0000011010010000" => data_out <= rom_array(1680);
		when "0000011010010001" => data_out <= rom_array(1681);
		when "0000011010010010" => data_out <= rom_array(1682);
		when "0000011010010011" => data_out <= rom_array(1683);
		when "0000011010010100" => data_out <= rom_array(1684);
		when "0000011010010101" => data_out <= rom_array(1685);
		when "0000011010010110" => data_out <= rom_array(1686);
		when "0000011010010111" => data_out <= rom_array(1687);
		when "0000011010011000" => data_out <= rom_array(1688);
		when "0000011010011001" => data_out <= rom_array(1689);
		when "0000011010011010" => data_out <= rom_array(1690);
		when "0000011010011011" => data_out <= rom_array(1691);
		when "0000011010011100" => data_out <= rom_array(1692);
		when "0000011010011101" => data_out <= rom_array(1693);
		when "0000011010011110" => data_out <= rom_array(1694);
		when "0000011010011111" => data_out <= rom_array(1695);
		when "0000011010100000" => data_out <= rom_array(1696);
		when "0000011010100001" => data_out <= rom_array(1697);
		when "0000011010100010" => data_out <= rom_array(1698);
		when "0000011010100011" => data_out <= rom_array(1699);
		when "0000011010100100" => data_out <= rom_array(1700);
		when "0000011010100101" => data_out <= rom_array(1701);
		when "0000011010100110" => data_out <= rom_array(1702);
		when "0000011010100111" => data_out <= rom_array(1703);
		when "0000011010101000" => data_out <= rom_array(1704);
		when "0000011010101001" => data_out <= rom_array(1705);
		when "0000011010101010" => data_out <= rom_array(1706);
		when "0000011010101011" => data_out <= rom_array(1707);
		when "0000011010101100" => data_out <= rom_array(1708);
		when "0000011010101101" => data_out <= rom_array(1709);
		when "0000011010101110" => data_out <= rom_array(1710);
		when "0000011010101111" => data_out <= rom_array(1711);
		when "0000011010110000" => data_out <= rom_array(1712);
		when "0000011010110001" => data_out <= rom_array(1713);
		when "0000011010110010" => data_out <= rom_array(1714);
		when "0000011010110011" => data_out <= rom_array(1715);
		when "0000011010110100" => data_out <= rom_array(1716);
		when "0000011010110101" => data_out <= rom_array(1717);
		when "0000011010110110" => data_out <= rom_array(1718);
		when "0000011010110111" => data_out <= rom_array(1719);
		when "0000011010111000" => data_out <= rom_array(1720);
		when "0000011010111001" => data_out <= rom_array(1721);
		when "0000011010111010" => data_out <= rom_array(1722);
		when "0000011010111011" => data_out <= rom_array(1723);
		when "0000011010111100" => data_out <= rom_array(1724);
		when "0000011010111101" => data_out <= rom_array(1725);
		when "0000011010111110" => data_out <= rom_array(1726);
		when "0000011010111111" => data_out <= rom_array(1727);
		when "0000011011000000" => data_out <= rom_array(1728);
		when "0000011011000001" => data_out <= rom_array(1729);
		when "0000011011000010" => data_out <= rom_array(1730);
		when "0000011011000011" => data_out <= rom_array(1731);
		when "0000011011000100" => data_out <= rom_array(1732);
		when "0000011011000101" => data_out <= rom_array(1733);
		when "0000011011000110" => data_out <= rom_array(1734);
		when "0000011011000111" => data_out <= rom_array(1735);
		when "0000011011001000" => data_out <= rom_array(1736);
		when "0000011011001001" => data_out <= rom_array(1737);
		when "0000011011001010" => data_out <= rom_array(1738);
		when "0000011011001011" => data_out <= rom_array(1739);
		when "0000011011001100" => data_out <= rom_array(1740);
		when "0000011011001101" => data_out <= rom_array(1741);
		when "0000011011001110" => data_out <= rom_array(1742);
		when "0000011011001111" => data_out <= rom_array(1743);
		when "0000011011010000" => data_out <= rom_array(1744);
		when "0000011011010001" => data_out <= rom_array(1745);
		when "0000011011010010" => data_out <= rom_array(1746);
		when "0000011011010011" => data_out <= rom_array(1747);
		when "0000011011010100" => data_out <= rom_array(1748);
		when "0000011011010101" => data_out <= rom_array(1749);
		when "0000011011010110" => data_out <= rom_array(1750);
		when "0000011011010111" => data_out <= rom_array(1751);
		when "0000011011011000" => data_out <= rom_array(1752);
		when "0000011011011001" => data_out <= rom_array(1753);
		when "0000011011011010" => data_out <= rom_array(1754);
		when "0000011011011011" => data_out <= rom_array(1755);
		when "0000011011011100" => data_out <= rom_array(1756);
		when "0000011011011101" => data_out <= rom_array(1757);
		when "0000011011011110" => data_out <= rom_array(1758);
		when "0000011011011111" => data_out <= rom_array(1759);
		when "0000011011100000" => data_out <= rom_array(1760);
		when "0000011011100001" => data_out <= rom_array(1761);
		when "0000011011100010" => data_out <= rom_array(1762);
		when "0000011011100011" => data_out <= rom_array(1763);
		when "0000011011100100" => data_out <= rom_array(1764);
		when "0000011011100101" => data_out <= rom_array(1765);
		when "0000011011100110" => data_out <= rom_array(1766);
		when "0000011011100111" => data_out <= rom_array(1767);
		when "0000011011101000" => data_out <= rom_array(1768);
		when "0000011011101001" => data_out <= rom_array(1769);
		when "0000011011101010" => data_out <= rom_array(1770);
		when "0000011011101011" => data_out <= rom_array(1771);
		when "0000011011101100" => data_out <= rom_array(1772);
		when "0000011011101101" => data_out <= rom_array(1773);
		when "0000011011101110" => data_out <= rom_array(1774);
		when "0000011011101111" => data_out <= rom_array(1775);
		when "0000011011110000" => data_out <= rom_array(1776);
		when "0000011011110001" => data_out <= rom_array(1777);
		when "0000011011110010" => data_out <= rom_array(1778);
		when "0000011011110011" => data_out <= rom_array(1779);
		when "0000011011110100" => data_out <= rom_array(1780);
		when "0000011011110101" => data_out <= rom_array(1781);
		when "0000011011110110" => data_out <= rom_array(1782);
		when "0000011011110111" => data_out <= rom_array(1783);
		when "0000011011111000" => data_out <= rom_array(1784);
		when "0000011011111001" => data_out <= rom_array(1785);
		when "0000011011111010" => data_out <= rom_array(1786);
		when "0000011011111011" => data_out <= rom_array(1787);
		when "0000011011111100" => data_out <= rom_array(1788);
		when "0000011011111101" => data_out <= rom_array(1789);
		when "0000011011111110" => data_out <= rom_array(1790);
		when "0000011011111111" => data_out <= rom_array(1791);
		when "0000011100000000" => data_out <= rom_array(1792);
		when "0000011100000001" => data_out <= rom_array(1793);
		when "0000011100000010" => data_out <= rom_array(1794);
		when "0000011100000011" => data_out <= rom_array(1795);
		when "0000011100000100" => data_out <= rom_array(1796);
		when "0000011100000101" => data_out <= rom_array(1797);
		when "0000011100000110" => data_out <= rom_array(1798);
		when "0000011100000111" => data_out <= rom_array(1799);
		when "0000011100001000" => data_out <= rom_array(1800);
		when "0000011100001001" => data_out <= rom_array(1801);
		when "0000011100001010" => data_out <= rom_array(1802);
		when "0000011100001011" => data_out <= rom_array(1803);
		when "0000011100001100" => data_out <= rom_array(1804);
		when "0000011100001101" => data_out <= rom_array(1805);
		when "0000011100001110" => data_out <= rom_array(1806);
		when "0000011100001111" => data_out <= rom_array(1807);
		when "0000011100010000" => data_out <= rom_array(1808);
		when "0000011100010001" => data_out <= rom_array(1809);
		when "0000011100010010" => data_out <= rom_array(1810);
		when "0000011100010011" => data_out <= rom_array(1811);
		when "0000011100010100" => data_out <= rom_array(1812);
		when "0000011100010101" => data_out <= rom_array(1813);
		when "0000011100010110" => data_out <= rom_array(1814);
		when "0000011100010111" => data_out <= rom_array(1815);
		when "0000011100011000" => data_out <= rom_array(1816);
		when "0000011100011001" => data_out <= rom_array(1817);
		when "0000011100011010" => data_out <= rom_array(1818);
		when "0000011100011011" => data_out <= rom_array(1819);
		when "0000011100011100" => data_out <= rom_array(1820);
		when "0000011100011101" => data_out <= rom_array(1821);
		when "0000011100011110" => data_out <= rom_array(1822);
		when "0000011100011111" => data_out <= rom_array(1823);
		when "0000011100100000" => data_out <= rom_array(1824);
		when "0000011100100001" => data_out <= rom_array(1825);
		when "0000011100100010" => data_out <= rom_array(1826);
		when "0000011100100011" => data_out <= rom_array(1827);
		when "0000011100100100" => data_out <= rom_array(1828);
		when "0000011100100101" => data_out <= rom_array(1829);
		when "0000011100100110" => data_out <= rom_array(1830);
		when "0000011100100111" => data_out <= rom_array(1831);
		when "0000011100101000" => data_out <= rom_array(1832);
		when "0000011100101001" => data_out <= rom_array(1833);
		when "0000011100101010" => data_out <= rom_array(1834);
		when "0000011100101011" => data_out <= rom_array(1835);
		when "0000011100101100" => data_out <= rom_array(1836);
		when "0000011100101101" => data_out <= rom_array(1837);
		when "0000011100101110" => data_out <= rom_array(1838);
		when "0000011100101111" => data_out <= rom_array(1839);
		when "0000011100110000" => data_out <= rom_array(1840);
		when "0000011100110001" => data_out <= rom_array(1841);
		when "0000011100110010" => data_out <= rom_array(1842);
		when "0000011100110011" => data_out <= rom_array(1843);
		when "0000011100110100" => data_out <= rom_array(1844);
		when "0000011100110101" => data_out <= rom_array(1845);
		when "0000011100110110" => data_out <= rom_array(1846);
		when "0000011100110111" => data_out <= rom_array(1847);
		when "0000011100111000" => data_out <= rom_array(1848);
		when "0000011100111001" => data_out <= rom_array(1849);
		when "0000011100111010" => data_out <= rom_array(1850);
		when "0000011100111011" => data_out <= rom_array(1851);
		when "0000011100111100" => data_out <= rom_array(1852);
		when "0000011100111101" => data_out <= rom_array(1853);
		when "0000011100111110" => data_out <= rom_array(1854);
		when "0000011100111111" => data_out <= rom_array(1855);
		when "0000011101000000" => data_out <= rom_array(1856);
		when "0000011101000001" => data_out <= rom_array(1857);
		when "0000011101000010" => data_out <= rom_array(1858);
		when "0000011101000011" => data_out <= rom_array(1859);
		when "0000011101000100" => data_out <= rom_array(1860);
		when "0000011101000101" => data_out <= rom_array(1861);
		when "0000011101000110" => data_out <= rom_array(1862);
		when "0000011101000111" => data_out <= rom_array(1863);
		when "0000011101001000" => data_out <= rom_array(1864);
		when "0000011101001001" => data_out <= rom_array(1865);
		when "0000011101001010" => data_out <= rom_array(1866);
		when "0000011101001011" => data_out <= rom_array(1867);
		when "0000011101001100" => data_out <= rom_array(1868);
		when "0000011101001101" => data_out <= rom_array(1869);
		when "0000011101001110" => data_out <= rom_array(1870);
		when "0000011101001111" => data_out <= rom_array(1871);
		when "0000011101010000" => data_out <= rom_array(1872);
		when "0000011101010001" => data_out <= rom_array(1873);
		when "0000011101010010" => data_out <= rom_array(1874);
		when "0000011101010011" => data_out <= rom_array(1875);
		when "0000011101010100" => data_out <= rom_array(1876);
		when "0000011101010101" => data_out <= rom_array(1877);
		when "0000011101010110" => data_out <= rom_array(1878);
		when "0000011101010111" => data_out <= rom_array(1879);
		when "0000011101011000" => data_out <= rom_array(1880);
		when "0000011101011001" => data_out <= rom_array(1881);
		when "0000011101011010" => data_out <= rom_array(1882);
		when "0000011101011011" => data_out <= rom_array(1883);
		when "0000011101011100" => data_out <= rom_array(1884);
		when "0000011101011101" => data_out <= rom_array(1885);
		when "0000011101011110" => data_out <= rom_array(1886);
		when "0000011101011111" => data_out <= rom_array(1887);
		when "0000011101100000" => data_out <= rom_array(1888);
		when "0000011101100001" => data_out <= rom_array(1889);
		when "0000011101100010" => data_out <= rom_array(1890);
		when "0000011101100011" => data_out <= rom_array(1891);
		when "0000011101100100" => data_out <= rom_array(1892);
		when "0000011101100101" => data_out <= rom_array(1893);
		when "0000011101100110" => data_out <= rom_array(1894);
		when "0000011101100111" => data_out <= rom_array(1895);
		when "0000011101101000" => data_out <= rom_array(1896);
		when "0000011101101001" => data_out <= rom_array(1897);
		when "0000011101101010" => data_out <= rom_array(1898);
		when "0000011101101011" => data_out <= rom_array(1899);
		when "0000011101101100" => data_out <= rom_array(1900);
		when "0000011101101101" => data_out <= rom_array(1901);
		when "0000011101101110" => data_out <= rom_array(1902);
		when "0000011101101111" => data_out <= rom_array(1903);
		when "0000011101110000" => data_out <= rom_array(1904);
		when "0000011101110001" => data_out <= rom_array(1905);
		when "0000011101110010" => data_out <= rom_array(1906);
		when "0000011101110011" => data_out <= rom_array(1907);
		when "0000011101110100" => data_out <= rom_array(1908);
		when "0000011101110101" => data_out <= rom_array(1909);
		when "0000011101110110" => data_out <= rom_array(1910);
		when "0000011101110111" => data_out <= rom_array(1911);
		when "0000011101111000" => data_out <= rom_array(1912);
		when "0000011101111001" => data_out <= rom_array(1913);
		when "0000011101111010" => data_out <= rom_array(1914);
		when "0000011101111011" => data_out <= rom_array(1915);
		when "0000011101111100" => data_out <= rom_array(1916);
		when "0000011101111101" => data_out <= rom_array(1917);
		when "0000011101111110" => data_out <= rom_array(1918);
		when "0000011101111111" => data_out <= rom_array(1919);
		when "0000011110000000" => data_out <= rom_array(1920);
		when "0000011110000001" => data_out <= rom_array(1921);
		when "0000011110000010" => data_out <= rom_array(1922);
		when "0000011110000011" => data_out <= rom_array(1923);
		when "0000011110000100" => data_out <= rom_array(1924);
		when "0000011110000101" => data_out <= rom_array(1925);
		when "0000011110000110" => data_out <= rom_array(1926);
		when "0000011110000111" => data_out <= rom_array(1927);
		when "0000011110001000" => data_out <= rom_array(1928);
		when "0000011110001001" => data_out <= rom_array(1929);
		when "0000011110001010" => data_out <= rom_array(1930);
		when "0000011110001011" => data_out <= rom_array(1931);
		when "0000011110001100" => data_out <= rom_array(1932);
		when "0000011110001101" => data_out <= rom_array(1933);
		when "0000011110001110" => data_out <= rom_array(1934);
		when "0000011110001111" => data_out <= rom_array(1935);
		when "0000011110010000" => data_out <= rom_array(1936);
		when "0000011110010001" => data_out <= rom_array(1937);
		when "0000011110010010" => data_out <= rom_array(1938);
		when "0000011110010011" => data_out <= rom_array(1939);
		when "0000011110010100" => data_out <= rom_array(1940);
		when "0000011110010101" => data_out <= rom_array(1941);
		when "0000011110010110" => data_out <= rom_array(1942);
		when "0000011110010111" => data_out <= rom_array(1943);
		when "0000011110011000" => data_out <= rom_array(1944);
		when "0000011110011001" => data_out <= rom_array(1945);
		when "0000011110011010" => data_out <= rom_array(1946);
		when "0000011110011011" => data_out <= rom_array(1947);
		when "0000011110011100" => data_out <= rom_array(1948);
		when "0000011110011101" => data_out <= rom_array(1949);
		when "0000011110011110" => data_out <= rom_array(1950);
		when "0000011110011111" => data_out <= rom_array(1951);
		when "0000011110100000" => data_out <= rom_array(1952);
		when "0000011110100001" => data_out <= rom_array(1953);
		when "0000011110100010" => data_out <= rom_array(1954);
		when "0000011110100011" => data_out <= rom_array(1955);
		when "0000011110100100" => data_out <= rom_array(1956);
		when "0000011110100101" => data_out <= rom_array(1957);
		when "0000011110100110" => data_out <= rom_array(1958);
		when "0000011110100111" => data_out <= rom_array(1959);
		when "0000011110101000" => data_out <= rom_array(1960);
		when "0000011110101001" => data_out <= rom_array(1961);
		when "0000011110101010" => data_out <= rom_array(1962);
		when "0000011110101011" => data_out <= rom_array(1963);
		when "0000011110101100" => data_out <= rom_array(1964);
		when "0000011110101101" => data_out <= rom_array(1965);
		when "0000011110101110" => data_out <= rom_array(1966);
		when "0000011110101111" => data_out <= rom_array(1967);
		when "0000011110110000" => data_out <= rom_array(1968);
		when "0000011110110001" => data_out <= rom_array(1969);
		when "0000011110110010" => data_out <= rom_array(1970);
		when "0000011110110011" => data_out <= rom_array(1971);
		when "0000011110110100" => data_out <= rom_array(1972);
		when "0000011110110101" => data_out <= rom_array(1973);
		when "0000011110110110" => data_out <= rom_array(1974);
		when "0000011110110111" => data_out <= rom_array(1975);
		when "0000011110111000" => data_out <= rom_array(1976);
		when "0000011110111001" => data_out <= rom_array(1977);
		when "0000011110111010" => data_out <= rom_array(1978);
		when "0000011110111011" => data_out <= rom_array(1979);
		when "0000011110111100" => data_out <= rom_array(1980);
		when "0000011110111101" => data_out <= rom_array(1981);
		when "0000011110111110" => data_out <= rom_array(1982);
		when "0000011110111111" => data_out <= rom_array(1983);
		when "0000011111000000" => data_out <= rom_array(1984);
		when "0000011111000001" => data_out <= rom_array(1985);
		when "0000011111000010" => data_out <= rom_array(1986);
		when "0000011111000011" => data_out <= rom_array(1987);
		when "0000011111000100" => data_out <= rom_array(1988);
		when "0000011111000101" => data_out <= rom_array(1989);
		when "0000011111000110" => data_out <= rom_array(1990);
		when "0000011111000111" => data_out <= rom_array(1991);
		when "0000011111001000" => data_out <= rom_array(1992);
		when "0000011111001001" => data_out <= rom_array(1993);
		when "0000011111001010" => data_out <= rom_array(1994);
		when "0000011111001011" => data_out <= rom_array(1995);
		when "0000011111001100" => data_out <= rom_array(1996);
		when "0000011111001101" => data_out <= rom_array(1997);
		when "0000011111001110" => data_out <= rom_array(1998);
		when "0000011111001111" => data_out <= rom_array(1999);
		when "0000011111010000" => data_out <= rom_array(2000);
		when "0000011111010001" => data_out <= rom_array(2001);
		when "0000011111010010" => data_out <= rom_array(2002);
		when "0000011111010011" => data_out <= rom_array(2003);
		when "0000011111010100" => data_out <= rom_array(2004);
		when "0000011111010101" => data_out <= rom_array(2005);
		when "0000011111010110" => data_out <= rom_array(2006);
		when "0000011111010111" => data_out <= rom_array(2007);
		when "0000011111011000" => data_out <= rom_array(2008);
		when "0000011111011001" => data_out <= rom_array(2009);
		when "0000011111011010" => data_out <= rom_array(2010);
		when "0000011111011011" => data_out <= rom_array(2011);
		when "0000011111011100" => data_out <= rom_array(2012);
		when "0000011111011101" => data_out <= rom_array(2013);
		when "0000011111011110" => data_out <= rom_array(2014);
		when "0000011111011111" => data_out <= rom_array(2015);
		when "0000011111100000" => data_out <= rom_array(2016);
		when "0000011111100001" => data_out <= rom_array(2017);
		when "0000011111100010" => data_out <= rom_array(2018);
		when "0000011111100011" => data_out <= rom_array(2019);
		when "0000011111100100" => data_out <= rom_array(2020);
		when "0000011111100101" => data_out <= rom_array(2021);
		when "0000011111100110" => data_out <= rom_array(2022);
		when "0000011111100111" => data_out <= rom_array(2023);
		when "0000011111101000" => data_out <= rom_array(2024);
		when "0000011111101001" => data_out <= rom_array(2025);
		when "0000011111101010" => data_out <= rom_array(2026);
		when "0000011111101011" => data_out <= rom_array(2027);
		when "0000011111101100" => data_out <= rom_array(2028);
		when "0000011111101101" => data_out <= rom_array(2029);
		when "0000011111101110" => data_out <= rom_array(2030);
		when "0000011111101111" => data_out <= rom_array(2031);
		when "0000011111110000" => data_out <= rom_array(2032);
		when "0000011111110001" => data_out <= rom_array(2033);
		when "0000011111110010" => data_out <= rom_array(2034);
		when "0000011111110011" => data_out <= rom_array(2035);
		when "0000011111110100" => data_out <= rom_array(2036);
		when "0000011111110101" => data_out <= rom_array(2037);
		when "0000011111110110" => data_out <= rom_array(2038);
		when "0000011111110111" => data_out <= rom_array(2039);
		when "0000011111111000" => data_out <= rom_array(2040);
		when "0000011111111001" => data_out <= rom_array(2041);
		when "0000011111111010" => data_out <= rom_array(2042);
		when "0000011111111011" => data_out <= rom_array(2043);
		when "0000011111111100" => data_out <= rom_array(2044);
		when "0000011111111101" => data_out <= rom_array(2045);
		when "0000011111111110" => data_out <= rom_array(2046);
		when "0000011111111111" => data_out <= rom_array(2047);
		when "0000100000000000" => data_out <= rom_array(2048);
		when "0000100000000001" => data_out <= rom_array(2049);
		when "0000100000000010" => data_out <= rom_array(2050);
		when "0000100000000011" => data_out <= rom_array(2051);
		when "0000100000000100" => data_out <= rom_array(2052);
		when "0000100000000101" => data_out <= rom_array(2053);
		when "0000100000000110" => data_out <= rom_array(2054);
		when "0000100000000111" => data_out <= rom_array(2055);
		when "0000100000001000" => data_out <= rom_array(2056);
		when "0000100000001001" => data_out <= rom_array(2057);
		when "0000100000001010" => data_out <= rom_array(2058);
		when "0000100000001011" => data_out <= rom_array(2059);
		when "0000100000001100" => data_out <= rom_array(2060);
		when "0000100000001101" => data_out <= rom_array(2061);
		when "0000100000001110" => data_out <= rom_array(2062);
		when "0000100000001111" => data_out <= rom_array(2063);
		when "0000100000010000" => data_out <= rom_array(2064);
		when "0000100000010001" => data_out <= rom_array(2065);
		when "0000100000010010" => data_out <= rom_array(2066);
		when "0000100000010011" => data_out <= rom_array(2067);
		when "0000100000010100" => data_out <= rom_array(2068);
		when "0000100000010101" => data_out <= rom_array(2069);
		when "0000100000010110" => data_out <= rom_array(2070);
		when "0000100000010111" => data_out <= rom_array(2071);
		when "0000100000011000" => data_out <= rom_array(2072);
		when "0000100000011001" => data_out <= rom_array(2073);
		when "0000100000011010" => data_out <= rom_array(2074);
		when "0000100000011011" => data_out <= rom_array(2075);
		when "0000100000011100" => data_out <= rom_array(2076);
		when "0000100000011101" => data_out <= rom_array(2077);
		when "0000100000011110" => data_out <= rom_array(2078);
		when "0000100000011111" => data_out <= rom_array(2079);
		when "0000100000100000" => data_out <= rom_array(2080);
		when "0000100000100001" => data_out <= rom_array(2081);
		when "0000100000100010" => data_out <= rom_array(2082);
		when "0000100000100011" => data_out <= rom_array(2083);
		when "0000100000100100" => data_out <= rom_array(2084);
		when "0000100000100101" => data_out <= rom_array(2085);
		when "0000100000100110" => data_out <= rom_array(2086);
		when "0000100000100111" => data_out <= rom_array(2087);
		when "0000100000101000" => data_out <= rom_array(2088);
		when "0000100000101001" => data_out <= rom_array(2089);
		when "0000100000101010" => data_out <= rom_array(2090);
		when "0000100000101011" => data_out <= rom_array(2091);
		when "0000100000101100" => data_out <= rom_array(2092);
		when "0000100000101101" => data_out <= rom_array(2093);
		when "0000100000101110" => data_out <= rom_array(2094);
		when "0000100000101111" => data_out <= rom_array(2095);
		when "0000100000110000" => data_out <= rom_array(2096);
		when "0000100000110001" => data_out <= rom_array(2097);
		when "0000100000110010" => data_out <= rom_array(2098);
		when "0000100000110011" => data_out <= rom_array(2099);
		when "0000100000110100" => data_out <= rom_array(2100);
		when "0000100000110101" => data_out <= rom_array(2101);
		when "0000100000110110" => data_out <= rom_array(2102);
		when "0000100000110111" => data_out <= rom_array(2103);
		when "0000100000111000" => data_out <= rom_array(2104);
		when "0000100000111001" => data_out <= rom_array(2105);
		when "0000100000111010" => data_out <= rom_array(2106);
		when "0000100000111011" => data_out <= rom_array(2107);
		when "0000100000111100" => data_out <= rom_array(2108);
		when "0000100000111101" => data_out <= rom_array(2109);
		when "0000100000111110" => data_out <= rom_array(2110);
		when "0000100000111111" => data_out <= rom_array(2111);
		when "0000100001000000" => data_out <= rom_array(2112);
		when "0000100001000001" => data_out <= rom_array(2113);
		when "0000100001000010" => data_out <= rom_array(2114);
		when "0000100001000011" => data_out <= rom_array(2115);
		when "0000100001000100" => data_out <= rom_array(2116);
		when "0000100001000101" => data_out <= rom_array(2117);
		when "0000100001000110" => data_out <= rom_array(2118);
		when "0000100001000111" => data_out <= rom_array(2119);
		when "0000100001001000" => data_out <= rom_array(2120);
		when "0000100001001001" => data_out <= rom_array(2121);
		when "0000100001001010" => data_out <= rom_array(2122);
		when "0000100001001011" => data_out <= rom_array(2123);
		when "0000100001001100" => data_out <= rom_array(2124);
		when "0000100001001101" => data_out <= rom_array(2125);
		when "0000100001001110" => data_out <= rom_array(2126);
		when "0000100001001111" => data_out <= rom_array(2127);
		when "0000100001010000" => data_out <= rom_array(2128);
		when "0000100001010001" => data_out <= rom_array(2129);
		when "0000100001010010" => data_out <= rom_array(2130);
		when "0000100001010011" => data_out <= rom_array(2131);
		when "0000100001010100" => data_out <= rom_array(2132);
		when "0000100001010101" => data_out <= rom_array(2133);
		when "0000100001010110" => data_out <= rom_array(2134);
		when "0000100001010111" => data_out <= rom_array(2135);
		when "0000100001011000" => data_out <= rom_array(2136);
		when "0000100001011001" => data_out <= rom_array(2137);
		when "0000100001011010" => data_out <= rom_array(2138);
		when "0000100001011011" => data_out <= rom_array(2139);
		when "0000100001011100" => data_out <= rom_array(2140);
		when "0000100001011101" => data_out <= rom_array(2141);
		when "0000100001011110" => data_out <= rom_array(2142);
		when "0000100001011111" => data_out <= rom_array(2143);
		when "0000100001100000" => data_out <= rom_array(2144);
		when "0000100001100001" => data_out <= rom_array(2145);
		when "0000100001100010" => data_out <= rom_array(2146);
		when "0000100001100011" => data_out <= rom_array(2147);
		when "0000100001100100" => data_out <= rom_array(2148);
		when "0000100001100101" => data_out <= rom_array(2149);
		when "0000100001100110" => data_out <= rom_array(2150);
		when "0000100001100111" => data_out <= rom_array(2151);
		when "0000100001101000" => data_out <= rom_array(2152);
		when "0000100001101001" => data_out <= rom_array(2153);
		when "0000100001101010" => data_out <= rom_array(2154);
		when "0000100001101011" => data_out <= rom_array(2155);
		when "0000100001101100" => data_out <= rom_array(2156);
		when "0000100001101101" => data_out <= rom_array(2157);
		when "0000100001101110" => data_out <= rom_array(2158);
		when "0000100001101111" => data_out <= rom_array(2159);
		when "0000100001110000" => data_out <= rom_array(2160);
		when "0000100001110001" => data_out <= rom_array(2161);
		when "0000100001110010" => data_out <= rom_array(2162);
		when "0000100001110011" => data_out <= rom_array(2163);
		when "0000100001110100" => data_out <= rom_array(2164);
		when "0000100001110101" => data_out <= rom_array(2165);
		when "0000100001110110" => data_out <= rom_array(2166);
		when "0000100001110111" => data_out <= rom_array(2167);
		when "0000100001111000" => data_out <= rom_array(2168);
		when "0000100001111001" => data_out <= rom_array(2169);
		when "0000100001111010" => data_out <= rom_array(2170);
		when "0000100001111011" => data_out <= rom_array(2171);
		when "0000100001111100" => data_out <= rom_array(2172);
		when "0000100001111101" => data_out <= rom_array(2173);
		when "0000100001111110" => data_out <= rom_array(2174);
		when "0000100001111111" => data_out <= rom_array(2175);
		when "0000100010000000" => data_out <= rom_array(2176);
		when "0000100010000001" => data_out <= rom_array(2177);
		when "0000100010000010" => data_out <= rom_array(2178);
		when "0000100010000011" => data_out <= rom_array(2179);
		when "0000100010000100" => data_out <= rom_array(2180);
		when "0000100010000101" => data_out <= rom_array(2181);
		when "0000100010000110" => data_out <= rom_array(2182);
		when "0000100010000111" => data_out <= rom_array(2183);
		when "0000100010001000" => data_out <= rom_array(2184);
		when "0000100010001001" => data_out <= rom_array(2185);
		when "0000100010001010" => data_out <= rom_array(2186);
		when "0000100010001011" => data_out <= rom_array(2187);
		when "0000100010001100" => data_out <= rom_array(2188);
		when "0000100010001101" => data_out <= rom_array(2189);
		when "0000100010001110" => data_out <= rom_array(2190);
		when "0000100010001111" => data_out <= rom_array(2191);
		when "0000100010010000" => data_out <= rom_array(2192);
		when "0000100010010001" => data_out <= rom_array(2193);
		when "0000100010010010" => data_out <= rom_array(2194);
		when "0000100010010011" => data_out <= rom_array(2195);
		when "0000100010010100" => data_out <= rom_array(2196);
		when "0000100010010101" => data_out <= rom_array(2197);
		when "0000100010010110" => data_out <= rom_array(2198);
		when "0000100010010111" => data_out <= rom_array(2199);
		when "0000100010011000" => data_out <= rom_array(2200);
		when "0000100010011001" => data_out <= rom_array(2201);
		when "0000100010011010" => data_out <= rom_array(2202);
		when "0000100010011011" => data_out <= rom_array(2203);
		when "0000100010011100" => data_out <= rom_array(2204);
		when "0000100010011101" => data_out <= rom_array(2205);
		when "0000100010011110" => data_out <= rom_array(2206);
		when "0000100010011111" => data_out <= rom_array(2207);
		when "0000100010100000" => data_out <= rom_array(2208);
		when "0000100010100001" => data_out <= rom_array(2209);
		when "0000100010100010" => data_out <= rom_array(2210);
		when "0000100010100011" => data_out <= rom_array(2211);
		when "0000100010100100" => data_out <= rom_array(2212);
		when "0000100010100101" => data_out <= rom_array(2213);
		when "0000100010100110" => data_out <= rom_array(2214);
		when "0000100010100111" => data_out <= rom_array(2215);
		when "0000100010101000" => data_out <= rom_array(2216);
		when "0000100010101001" => data_out <= rom_array(2217);
		when "0000100010101010" => data_out <= rom_array(2218);
		when "0000100010101011" => data_out <= rom_array(2219);
		when "0000100010101100" => data_out <= rom_array(2220);
		when "0000100010101101" => data_out <= rom_array(2221);
		when "0000100010101110" => data_out <= rom_array(2222);
		when "0000100010101111" => data_out <= rom_array(2223);
		when "0000100010110000" => data_out <= rom_array(2224);
		when "0000100010110001" => data_out <= rom_array(2225);
		when "0000100010110010" => data_out <= rom_array(2226);
		when "0000100010110011" => data_out <= rom_array(2227);
		when "0000100010110100" => data_out <= rom_array(2228);
		when "0000100010110101" => data_out <= rom_array(2229);
		when "0000100010110110" => data_out <= rom_array(2230);
		when "0000100010110111" => data_out <= rom_array(2231);
		when "0000100010111000" => data_out <= rom_array(2232);
		when "0000100010111001" => data_out <= rom_array(2233);
		when "0000100010111010" => data_out <= rom_array(2234);
		when "0000100010111011" => data_out <= rom_array(2235);
		when "0000100010111100" => data_out <= rom_array(2236);
		when "0000100010111101" => data_out <= rom_array(2237);
		when "0000100010111110" => data_out <= rom_array(2238);
		when "0000100010111111" => data_out <= rom_array(2239);
		when "0000100011000000" => data_out <= rom_array(2240);
		when "0000100011000001" => data_out <= rom_array(2241);
		when "0000100011000010" => data_out <= rom_array(2242);
		when "0000100011000011" => data_out <= rom_array(2243);
		when "0000100011000100" => data_out <= rom_array(2244);
		when "0000100011000101" => data_out <= rom_array(2245);
		when "0000100011000110" => data_out <= rom_array(2246);
		when "0000100011000111" => data_out <= rom_array(2247);
		when "0000100011001000" => data_out <= rom_array(2248);
		when "0000100011001001" => data_out <= rom_array(2249);
		when "0000100011001010" => data_out <= rom_array(2250);
		when "0000100011001011" => data_out <= rom_array(2251);
		when "0000100011001100" => data_out <= rom_array(2252);
		when "0000100011001101" => data_out <= rom_array(2253);
		when "0000100011001110" => data_out <= rom_array(2254);
		when "0000100011001111" => data_out <= rom_array(2255);
		when "0000100011010000" => data_out <= rom_array(2256);
		when "0000100011010001" => data_out <= rom_array(2257);
		when "0000100011010010" => data_out <= rom_array(2258);
		when "0000100011010011" => data_out <= rom_array(2259);
		when "0000100011010100" => data_out <= rom_array(2260);
		when "0000100011010101" => data_out <= rom_array(2261);
		when "0000100011010110" => data_out <= rom_array(2262);
		when "0000100011010111" => data_out <= rom_array(2263);
		when "0000100011011000" => data_out <= rom_array(2264);
		when "0000100011011001" => data_out <= rom_array(2265);
		when "0000100011011010" => data_out <= rom_array(2266);
		when "0000100011011011" => data_out <= rom_array(2267);
		when "0000100011011100" => data_out <= rom_array(2268);
		when "0000100011011101" => data_out <= rom_array(2269);
		when "0000100011011110" => data_out <= rom_array(2270);
		when "0000100011011111" => data_out <= rom_array(2271);
		when "0000100011100000" => data_out <= rom_array(2272);
		when "0000100011100001" => data_out <= rom_array(2273);
		when "0000100011100010" => data_out <= rom_array(2274);
		when "0000100011100011" => data_out <= rom_array(2275);
		when "0000100011100100" => data_out <= rom_array(2276);
		when "0000100011100101" => data_out <= rom_array(2277);
		when "0000100011100110" => data_out <= rom_array(2278);
		when "0000100011100111" => data_out <= rom_array(2279);
		when "0000100011101000" => data_out <= rom_array(2280);
		when "0000100011101001" => data_out <= rom_array(2281);
		when "0000100011101010" => data_out <= rom_array(2282);
		when "0000100011101011" => data_out <= rom_array(2283);
		when "0000100011101100" => data_out <= rom_array(2284);
		when "0000100011101101" => data_out <= rom_array(2285);
		when "0000100011101110" => data_out <= rom_array(2286);
		when "0000100011101111" => data_out <= rom_array(2287);
		when "0000100011110000" => data_out <= rom_array(2288);
		when "0000100011110001" => data_out <= rom_array(2289);
		when "0000100011110010" => data_out <= rom_array(2290);
		when "0000100011110011" => data_out <= rom_array(2291);
		when "0000100011110100" => data_out <= rom_array(2292);
		when "0000100011110101" => data_out <= rom_array(2293);
		when "0000100011110110" => data_out <= rom_array(2294);
		when "0000100011110111" => data_out <= rom_array(2295);
		when "0000100011111000" => data_out <= rom_array(2296);
		when "0000100011111001" => data_out <= rom_array(2297);
		when "0000100011111010" => data_out <= rom_array(2298);
		when "0000100011111011" => data_out <= rom_array(2299);
		when "0000100011111100" => data_out <= rom_array(2300);
		when "0000100011111101" => data_out <= rom_array(2301);
		when "0000100011111110" => data_out <= rom_array(2302);
		when "0000100011111111" => data_out <= rom_array(2303);
		when "0000100100000000" => data_out <= rom_array(2304);
		when "0000100100000001" => data_out <= rom_array(2305);
		when "0000100100000010" => data_out <= rom_array(2306);
		when "0000100100000011" => data_out <= rom_array(2307);
		when "0000100100000100" => data_out <= rom_array(2308);
		when "0000100100000101" => data_out <= rom_array(2309);
		when "0000100100000110" => data_out <= rom_array(2310);
		when "0000100100000111" => data_out <= rom_array(2311);
		when "0000100100001000" => data_out <= rom_array(2312);
		when "0000100100001001" => data_out <= rom_array(2313);
		when "0000100100001010" => data_out <= rom_array(2314);
		when "0000100100001011" => data_out <= rom_array(2315);
		when "0000100100001100" => data_out <= rom_array(2316);
		when "0000100100001101" => data_out <= rom_array(2317);
		when "0000100100001110" => data_out <= rom_array(2318);
		when "0000100100001111" => data_out <= rom_array(2319);
		when "0000100100010000" => data_out <= rom_array(2320);
		when "0000100100010001" => data_out <= rom_array(2321);
		when "0000100100010010" => data_out <= rom_array(2322);
		when "0000100100010011" => data_out <= rom_array(2323);
		when "0000100100010100" => data_out <= rom_array(2324);
		when "0000100100010101" => data_out <= rom_array(2325);
		when "0000100100010110" => data_out <= rom_array(2326);
		when "0000100100010111" => data_out <= rom_array(2327);
		when "0000100100011000" => data_out <= rom_array(2328);
		when "0000100100011001" => data_out <= rom_array(2329);
		when "0000100100011010" => data_out <= rom_array(2330);
		when "0000100100011011" => data_out <= rom_array(2331);
		when "0000100100011100" => data_out <= rom_array(2332);
		when "0000100100011101" => data_out <= rom_array(2333);
		when "0000100100011110" => data_out <= rom_array(2334);
		when "0000100100011111" => data_out <= rom_array(2335);
		when "0000100100100000" => data_out <= rom_array(2336);
		when "0000100100100001" => data_out <= rom_array(2337);
		when "0000100100100010" => data_out <= rom_array(2338);
		when "0000100100100011" => data_out <= rom_array(2339);
		when "0000100100100100" => data_out <= rom_array(2340);
		when "0000100100100101" => data_out <= rom_array(2341);
		when "0000100100100110" => data_out <= rom_array(2342);
		when "0000100100100111" => data_out <= rom_array(2343);
		when "0000100100101000" => data_out <= rom_array(2344);
		when "0000100100101001" => data_out <= rom_array(2345);
		when "0000100100101010" => data_out <= rom_array(2346);
		when "0000100100101011" => data_out <= rom_array(2347);
		when "0000100100101100" => data_out <= rom_array(2348);
		when "0000100100101101" => data_out <= rom_array(2349);
		when "0000100100101110" => data_out <= rom_array(2350);
		when "0000100100101111" => data_out <= rom_array(2351);
		when "0000100100110000" => data_out <= rom_array(2352);
		when "0000100100110001" => data_out <= rom_array(2353);
		when "0000100100110010" => data_out <= rom_array(2354);
		when "0000100100110011" => data_out <= rom_array(2355);
		when "0000100100110100" => data_out <= rom_array(2356);
		when "0000100100110101" => data_out <= rom_array(2357);
		when "0000100100110110" => data_out <= rom_array(2358);
		when "0000100100110111" => data_out <= rom_array(2359);
		when "0000100100111000" => data_out <= rom_array(2360);
		when "0000100100111001" => data_out <= rom_array(2361);
		when "0000100100111010" => data_out <= rom_array(2362);
		when "0000100100111011" => data_out <= rom_array(2363);
		when "0000100100111100" => data_out <= rom_array(2364);
		when "0000100100111101" => data_out <= rom_array(2365);
		when "0000100100111110" => data_out <= rom_array(2366);
		when "0000100100111111" => data_out <= rom_array(2367);
		when "0000100101000000" => data_out <= rom_array(2368);
		when "0000100101000001" => data_out <= rom_array(2369);
		when "0000100101000010" => data_out <= rom_array(2370);
		when "0000100101000011" => data_out <= rom_array(2371);
		when "0000100101000100" => data_out <= rom_array(2372);
		when "0000100101000101" => data_out <= rom_array(2373);
		when "0000100101000110" => data_out <= rom_array(2374);
		when "0000100101000111" => data_out <= rom_array(2375);
		when "0000100101001000" => data_out <= rom_array(2376);
		when "0000100101001001" => data_out <= rom_array(2377);
		when "0000100101001010" => data_out <= rom_array(2378);
		when "0000100101001011" => data_out <= rom_array(2379);
		when "0000100101001100" => data_out <= rom_array(2380);
		when "0000100101001101" => data_out <= rom_array(2381);
		when "0000100101001110" => data_out <= rom_array(2382);
		when "0000100101001111" => data_out <= rom_array(2383);
		when "0000100101010000" => data_out <= rom_array(2384);
		when "0000100101010001" => data_out <= rom_array(2385);
		when "0000100101010010" => data_out <= rom_array(2386);
		when "0000100101010011" => data_out <= rom_array(2387);
		when "0000100101010100" => data_out <= rom_array(2388);
		when "0000100101010101" => data_out <= rom_array(2389);
		when "0000100101010110" => data_out <= rom_array(2390);
		when "0000100101010111" => data_out <= rom_array(2391);
		when "0000100101011000" => data_out <= rom_array(2392);
		when "0000100101011001" => data_out <= rom_array(2393);
		when "0000100101011010" => data_out <= rom_array(2394);
		when "0000100101011011" => data_out <= rom_array(2395);
		when "0000100101011100" => data_out <= rom_array(2396);
		when "0000100101011101" => data_out <= rom_array(2397);
		when "0000100101011110" => data_out <= rom_array(2398);
		when "0000100101011111" => data_out <= rom_array(2399);
		when "0000100101100000" => data_out <= rom_array(2400);
		when "0000100101100001" => data_out <= rom_array(2401);
		when "0000100101100010" => data_out <= rom_array(2402);
		when "0000100101100011" => data_out <= rom_array(2403);
		when "0000100101100100" => data_out <= rom_array(2404);
		when "0000100101100101" => data_out <= rom_array(2405);
		when "0000100101100110" => data_out <= rom_array(2406);
		when "0000100101100111" => data_out <= rom_array(2407);
		when "0000100101101000" => data_out <= rom_array(2408);
		when "0000100101101001" => data_out <= rom_array(2409);
		when "0000100101101010" => data_out <= rom_array(2410);
		when "0000100101101011" => data_out <= rom_array(2411);
		when "0000100101101100" => data_out <= rom_array(2412);
		when "0000100101101101" => data_out <= rom_array(2413);
		when "0000100101101110" => data_out <= rom_array(2414);
		when "0000100101101111" => data_out <= rom_array(2415);
		when "0000100101110000" => data_out <= rom_array(2416);
		when "0000100101110001" => data_out <= rom_array(2417);
		when "0000100101110010" => data_out <= rom_array(2418);
		when "0000100101110011" => data_out <= rom_array(2419);
		when "0000100101110100" => data_out <= rom_array(2420);
		when "0000100101110101" => data_out <= rom_array(2421);
		when "0000100101110110" => data_out <= rom_array(2422);
		when "0000100101110111" => data_out <= rom_array(2423);
		when "0000100101111000" => data_out <= rom_array(2424);
		when "0000100101111001" => data_out <= rom_array(2425);
		when "0000100101111010" => data_out <= rom_array(2426);
		when "0000100101111011" => data_out <= rom_array(2427);
		when "0000100101111100" => data_out <= rom_array(2428);
		when "0000100101111101" => data_out <= rom_array(2429);
		when "0000100101111110" => data_out <= rom_array(2430);
		when "0000100101111111" => data_out <= rom_array(2431);
		when "0000100110000000" => data_out <= rom_array(2432);
		when "0000100110000001" => data_out <= rom_array(2433);
		when "0000100110000010" => data_out <= rom_array(2434);
		when "0000100110000011" => data_out <= rom_array(2435);
		when "0000100110000100" => data_out <= rom_array(2436);
		when "0000100110000101" => data_out <= rom_array(2437);
		when "0000100110000110" => data_out <= rom_array(2438);
		when "0000100110000111" => data_out <= rom_array(2439);
		when "0000100110001000" => data_out <= rom_array(2440);
		when "0000100110001001" => data_out <= rom_array(2441);
		when "0000100110001010" => data_out <= rom_array(2442);
		when "0000100110001011" => data_out <= rom_array(2443);
		when "0000100110001100" => data_out <= rom_array(2444);
		when "0000100110001101" => data_out <= rom_array(2445);
		when "0000100110001110" => data_out <= rom_array(2446);
		when "0000100110001111" => data_out <= rom_array(2447);
		when "0000100110010000" => data_out <= rom_array(2448);
		when "0000100110010001" => data_out <= rom_array(2449);
		when "0000100110010010" => data_out <= rom_array(2450);
		when "0000100110010011" => data_out <= rom_array(2451);
		when "0000100110010100" => data_out <= rom_array(2452);
		when "0000100110010101" => data_out <= rom_array(2453);
		when "0000100110010110" => data_out <= rom_array(2454);
		when "0000100110010111" => data_out <= rom_array(2455);
		when "0000100110011000" => data_out <= rom_array(2456);
		when "0000100110011001" => data_out <= rom_array(2457);
		when "0000100110011010" => data_out <= rom_array(2458);
		when "0000100110011011" => data_out <= rom_array(2459);
		when "0000100110011100" => data_out <= rom_array(2460);
		when "0000100110011101" => data_out <= rom_array(2461);
		when "0000100110011110" => data_out <= rom_array(2462);
		when "0000100110011111" => data_out <= rom_array(2463);
		when "0000100110100000" => data_out <= rom_array(2464);
		when "0000100110100001" => data_out <= rom_array(2465);
		when "0000100110100010" => data_out <= rom_array(2466);
		when "0000100110100011" => data_out <= rom_array(2467);
		when "0000100110100100" => data_out <= rom_array(2468);
		when "0000100110100101" => data_out <= rom_array(2469);
		when "0000100110100110" => data_out <= rom_array(2470);
		when "0000100110100111" => data_out <= rom_array(2471);
		when "0000100110101000" => data_out <= rom_array(2472);
		when "0000100110101001" => data_out <= rom_array(2473);
		when "0000100110101010" => data_out <= rom_array(2474);
		when "0000100110101011" => data_out <= rom_array(2475);
		when "0000100110101100" => data_out <= rom_array(2476);
		when "0000100110101101" => data_out <= rom_array(2477);
		when "0000100110101110" => data_out <= rom_array(2478);
		when "0000100110101111" => data_out <= rom_array(2479);
		when "0000100110110000" => data_out <= rom_array(2480);
		when "0000100110110001" => data_out <= rom_array(2481);
		when "0000100110110010" => data_out <= rom_array(2482);
		when "0000100110110011" => data_out <= rom_array(2483);
		when "0000100110110100" => data_out <= rom_array(2484);
		when "0000100110110101" => data_out <= rom_array(2485);
		when "0000100110110110" => data_out <= rom_array(2486);
		when "0000100110110111" => data_out <= rom_array(2487);
		when "0000100110111000" => data_out <= rom_array(2488);
		when "0000100110111001" => data_out <= rom_array(2489);
		when "0000100110111010" => data_out <= rom_array(2490);
		when "0000100110111011" => data_out <= rom_array(2491);
		when "0000100110111100" => data_out <= rom_array(2492);
		when "0000100110111101" => data_out <= rom_array(2493);
		when "0000100110111110" => data_out <= rom_array(2494);
		when "0000100110111111" => data_out <= rom_array(2495);
		when "0000100111000000" => data_out <= rom_array(2496);
		when "0000100111000001" => data_out <= rom_array(2497);
		when "0000100111000010" => data_out <= rom_array(2498);
		when "0000100111000011" => data_out <= rom_array(2499);
		when "0000100111000100" => data_out <= rom_array(2500);
		when "0000100111000101" => data_out <= rom_array(2501);
		when "0000100111000110" => data_out <= rom_array(2502);
		when "0000100111000111" => data_out <= rom_array(2503);
		when "0000100111001000" => data_out <= rom_array(2504);
		when "0000100111001001" => data_out <= rom_array(2505);
		when "0000100111001010" => data_out <= rom_array(2506);
		when "0000100111001011" => data_out <= rom_array(2507);
		when "0000100111001100" => data_out <= rom_array(2508);
		when "0000100111001101" => data_out <= rom_array(2509);
		when "0000100111001110" => data_out <= rom_array(2510);
		when "0000100111001111" => data_out <= rom_array(2511);
		when "0000100111010000" => data_out <= rom_array(2512);
		when "0000100111010001" => data_out <= rom_array(2513);
		when "0000100111010010" => data_out <= rom_array(2514);
		when "0000100111010011" => data_out <= rom_array(2515);
		when "0000100111010100" => data_out <= rom_array(2516);
		when "0000100111010101" => data_out <= rom_array(2517);
		when "0000100111010110" => data_out <= rom_array(2518);
		when "0000100111010111" => data_out <= rom_array(2519);
		when "0000100111011000" => data_out <= rom_array(2520);
		when "0000100111011001" => data_out <= rom_array(2521);
		when "0000100111011010" => data_out <= rom_array(2522);
		when "0000100111011011" => data_out <= rom_array(2523);
		when "0000100111011100" => data_out <= rom_array(2524);
		when "0000100111011101" => data_out <= rom_array(2525);
		when "0000100111011110" => data_out <= rom_array(2526);
		when "0000100111011111" => data_out <= rom_array(2527);
		when "0000100111100000" => data_out <= rom_array(2528);
		when "0000100111100001" => data_out <= rom_array(2529);
		when "0000100111100010" => data_out <= rom_array(2530);
		when "0000100111100011" => data_out <= rom_array(2531);
		when "0000100111100100" => data_out <= rom_array(2532);
		when "0000100111100101" => data_out <= rom_array(2533);
		when "0000100111100110" => data_out <= rom_array(2534);
		when "0000100111100111" => data_out <= rom_array(2535);
		when "0000100111101000" => data_out <= rom_array(2536);
		when "0000100111101001" => data_out <= rom_array(2537);
		when "0000100111101010" => data_out <= rom_array(2538);
		when "0000100111101011" => data_out <= rom_array(2539);
		when "0000100111101100" => data_out <= rom_array(2540);
		when "0000100111101101" => data_out <= rom_array(2541);
		when "0000100111101110" => data_out <= rom_array(2542);
		when "0000100111101111" => data_out <= rom_array(2543);
		when "0000100111110000" => data_out <= rom_array(2544);
		when "0000100111110001" => data_out <= rom_array(2545);
		when "0000100111110010" => data_out <= rom_array(2546);
		when "0000100111110011" => data_out <= rom_array(2547);
		when "0000100111110100" => data_out <= rom_array(2548);
		when "0000100111110101" => data_out <= rom_array(2549);
		when "0000100111110110" => data_out <= rom_array(2550);
		when "0000100111110111" => data_out <= rom_array(2551);
		when "0000100111111000" => data_out <= rom_array(2552);
		when "0000100111111001" => data_out <= rom_array(2553);
		when "0000100111111010" => data_out <= rom_array(2554);
		when "0000100111111011" => data_out <= rom_array(2555);
		when "0000100111111100" => data_out <= rom_array(2556);
		when "0000100111111101" => data_out <= rom_array(2557);
		when "0000100111111110" => data_out <= rom_array(2558);
		when "0000100111111111" => data_out <= rom_array(2559);
		when "0000101000000000" => data_out <= rom_array(2560);
		when "0000101000000001" => data_out <= rom_array(2561);
		when "0000101000000010" => data_out <= rom_array(2562);
		when "0000101000000011" => data_out <= rom_array(2563);
		when "0000101000000100" => data_out <= rom_array(2564);
		when "0000101000000101" => data_out <= rom_array(2565);
		when "0000101000000110" => data_out <= rom_array(2566);
		when "0000101000000111" => data_out <= rom_array(2567);
		when "0000101000001000" => data_out <= rom_array(2568);
		when "0000101000001001" => data_out <= rom_array(2569);
		when "0000101000001010" => data_out <= rom_array(2570);
		when "0000101000001011" => data_out <= rom_array(2571);
		when "0000101000001100" => data_out <= rom_array(2572);
		when "0000101000001101" => data_out <= rom_array(2573);
		when "0000101000001110" => data_out <= rom_array(2574);
		when "0000101000001111" => data_out <= rom_array(2575);
		when "0000101000010000" => data_out <= rom_array(2576);
		when "0000101000010001" => data_out <= rom_array(2577);
		when "0000101000010010" => data_out <= rom_array(2578);
		when "0000101000010011" => data_out <= rom_array(2579);
		when "0000101000010100" => data_out <= rom_array(2580);
		when "0000101000010101" => data_out <= rom_array(2581);
		when "0000101000010110" => data_out <= rom_array(2582);
		when "0000101000010111" => data_out <= rom_array(2583);
		when "0000101000011000" => data_out <= rom_array(2584);
		when "0000101000011001" => data_out <= rom_array(2585);
		when "0000101000011010" => data_out <= rom_array(2586);
		when "0000101000011011" => data_out <= rom_array(2587);
		when "0000101000011100" => data_out <= rom_array(2588);
		when "0000101000011101" => data_out <= rom_array(2589);
		when "0000101000011110" => data_out <= rom_array(2590);
		when "0000101000011111" => data_out <= rom_array(2591);
		when "0000101000100000" => data_out <= rom_array(2592);
		when "0000101000100001" => data_out <= rom_array(2593);
		when "0000101000100010" => data_out <= rom_array(2594);
		when "0000101000100011" => data_out <= rom_array(2595);
		when "0000101000100100" => data_out <= rom_array(2596);
		when "0000101000100101" => data_out <= rom_array(2597);
		when "0000101000100110" => data_out <= rom_array(2598);
		when "0000101000100111" => data_out <= rom_array(2599);
		when "0000101000101000" => data_out <= rom_array(2600);
		when "0000101000101001" => data_out <= rom_array(2601);
		when "0000101000101010" => data_out <= rom_array(2602);
		when "0000101000101011" => data_out <= rom_array(2603);
		when "0000101000101100" => data_out <= rom_array(2604);
		when "0000101000101101" => data_out <= rom_array(2605);
		when "0000101000101110" => data_out <= rom_array(2606);
		when "0000101000101111" => data_out <= rom_array(2607);
		when "0000101000110000" => data_out <= rom_array(2608);
		when "0000101000110001" => data_out <= rom_array(2609);
		when "0000101000110010" => data_out <= rom_array(2610);
		when "0000101000110011" => data_out <= rom_array(2611);
		when "0000101000110100" => data_out <= rom_array(2612);
		when "0000101000110101" => data_out <= rom_array(2613);
		when "0000101000110110" => data_out <= rom_array(2614);
		when "0000101000110111" => data_out <= rom_array(2615);
		when "0000101000111000" => data_out <= rom_array(2616);
		when "0000101000111001" => data_out <= rom_array(2617);
		when "0000101000111010" => data_out <= rom_array(2618);
		when "0000101000111011" => data_out <= rom_array(2619);
		when "0000101000111100" => data_out <= rom_array(2620);
		when "0000101000111101" => data_out <= rom_array(2621);
		when "0000101000111110" => data_out <= rom_array(2622);
		when "0000101000111111" => data_out <= rom_array(2623);
		when "0000101001000000" => data_out <= rom_array(2624);
		when "0000101001000001" => data_out <= rom_array(2625);
		when "0000101001000010" => data_out <= rom_array(2626);
		when "0000101001000011" => data_out <= rom_array(2627);
		when "0000101001000100" => data_out <= rom_array(2628);
		when "0000101001000101" => data_out <= rom_array(2629);
		when "0000101001000110" => data_out <= rom_array(2630);
		when "0000101001000111" => data_out <= rom_array(2631);
		when "0000101001001000" => data_out <= rom_array(2632);
		when "0000101001001001" => data_out <= rom_array(2633);
		when "0000101001001010" => data_out <= rom_array(2634);
		when "0000101001001011" => data_out <= rom_array(2635);
		when "0000101001001100" => data_out <= rom_array(2636);
		when "0000101001001101" => data_out <= rom_array(2637);
		when "0000101001001110" => data_out <= rom_array(2638);
		when "0000101001001111" => data_out <= rom_array(2639);
		when "0000101001010000" => data_out <= rom_array(2640);
		when "0000101001010001" => data_out <= rom_array(2641);
		when "0000101001010010" => data_out <= rom_array(2642);
		when "0000101001010011" => data_out <= rom_array(2643);
		when "0000101001010100" => data_out <= rom_array(2644);
		when "0000101001010101" => data_out <= rom_array(2645);
		when "0000101001010110" => data_out <= rom_array(2646);
		when "0000101001010111" => data_out <= rom_array(2647);
		when "0000101001011000" => data_out <= rom_array(2648);
		when "0000101001011001" => data_out <= rom_array(2649);
		when "0000101001011010" => data_out <= rom_array(2650);
		when "0000101001011011" => data_out <= rom_array(2651);
		when "0000101001011100" => data_out <= rom_array(2652);
		when "0000101001011101" => data_out <= rom_array(2653);
		when "0000101001011110" => data_out <= rom_array(2654);
		when "0000101001011111" => data_out <= rom_array(2655);
		when "0000101001100000" => data_out <= rom_array(2656);
		when "0000101001100001" => data_out <= rom_array(2657);
		when "0000101001100010" => data_out <= rom_array(2658);
		when "0000101001100011" => data_out <= rom_array(2659);
		when "0000101001100100" => data_out <= rom_array(2660);
		when "0000101001100101" => data_out <= rom_array(2661);
		when "0000101001100110" => data_out <= rom_array(2662);
		when "0000101001100111" => data_out <= rom_array(2663);
		when "0000101001101000" => data_out <= rom_array(2664);
		when "0000101001101001" => data_out <= rom_array(2665);
		when "0000101001101010" => data_out <= rom_array(2666);
		when "0000101001101011" => data_out <= rom_array(2667);
		when "0000101001101100" => data_out <= rom_array(2668);
		when "0000101001101101" => data_out <= rom_array(2669);
		when "0000101001101110" => data_out <= rom_array(2670);
		when "0000101001101111" => data_out <= rom_array(2671);
		when "0000101001110000" => data_out <= rom_array(2672);
		when "0000101001110001" => data_out <= rom_array(2673);
		when "0000101001110010" => data_out <= rom_array(2674);
		when "0000101001110011" => data_out <= rom_array(2675);
		when "0000101001110100" => data_out <= rom_array(2676);
		when "0000101001110101" => data_out <= rom_array(2677);
		when "0000101001110110" => data_out <= rom_array(2678);
		when "0000101001110111" => data_out <= rom_array(2679);
		when "0000101001111000" => data_out <= rom_array(2680);
		when "0000101001111001" => data_out <= rom_array(2681);
		when "0000101001111010" => data_out <= rom_array(2682);
		when "0000101001111011" => data_out <= rom_array(2683);
		when "0000101001111100" => data_out <= rom_array(2684);
		when "0000101001111101" => data_out <= rom_array(2685);
		when "0000101001111110" => data_out <= rom_array(2686);
		when "0000101001111111" => data_out <= rom_array(2687);
		when "0000101010000000" => data_out <= rom_array(2688);
		when "0000101010000001" => data_out <= rom_array(2689);
		when "0000101010000010" => data_out <= rom_array(2690);
		when "0000101010000011" => data_out <= rom_array(2691);
		when "0000101010000100" => data_out <= rom_array(2692);
		when "0000101010000101" => data_out <= rom_array(2693);
		when "0000101010000110" => data_out <= rom_array(2694);
		when "0000101010000111" => data_out <= rom_array(2695);
		when "0000101010001000" => data_out <= rom_array(2696);
		when "0000101010001001" => data_out <= rom_array(2697);
		when "0000101010001010" => data_out <= rom_array(2698);
		when "0000101010001011" => data_out <= rom_array(2699);
		when "0000101010001100" => data_out <= rom_array(2700);
		when "0000101010001101" => data_out <= rom_array(2701);
		when "0000101010001110" => data_out <= rom_array(2702);
		when "0000101010001111" => data_out <= rom_array(2703);
		when "0000101010010000" => data_out <= rom_array(2704);
		when "0000101010010001" => data_out <= rom_array(2705);
		when "0000101010010010" => data_out <= rom_array(2706);
		when "0000101010010011" => data_out <= rom_array(2707);
		when "0000101010010100" => data_out <= rom_array(2708);
		when "0000101010010101" => data_out <= rom_array(2709);
		when "0000101010010110" => data_out <= rom_array(2710);
		when "0000101010010111" => data_out <= rom_array(2711);
		when "0000101010011000" => data_out <= rom_array(2712);
		when "0000101010011001" => data_out <= rom_array(2713);
		when "0000101010011010" => data_out <= rom_array(2714);
		when "0000101010011011" => data_out <= rom_array(2715);
		when "0000101010011100" => data_out <= rom_array(2716);
		when "0000101010011101" => data_out <= rom_array(2717);
		when "0000101010011110" => data_out <= rom_array(2718);
		when "0000101010011111" => data_out <= rom_array(2719);
		when "0000101010100000" => data_out <= rom_array(2720);
		when "0000101010100001" => data_out <= rom_array(2721);
		when "0000101010100010" => data_out <= rom_array(2722);
		when "0000101010100011" => data_out <= rom_array(2723);
		when "0000101010100100" => data_out <= rom_array(2724);
		when "0000101010100101" => data_out <= rom_array(2725);
		when "0000101010100110" => data_out <= rom_array(2726);
		when "0000101010100111" => data_out <= rom_array(2727);
		when "0000101010101000" => data_out <= rom_array(2728);
		when "0000101010101001" => data_out <= rom_array(2729);
		when "0000101010101010" => data_out <= rom_array(2730);
		when "0000101010101011" => data_out <= rom_array(2731);
		when "0000101010101100" => data_out <= rom_array(2732);
		when "0000101010101101" => data_out <= rom_array(2733);
		when "0000101010101110" => data_out <= rom_array(2734);
		when "0000101010101111" => data_out <= rom_array(2735);
		when "0000101010110000" => data_out <= rom_array(2736);
		when "0000101010110001" => data_out <= rom_array(2737);
		when "0000101010110010" => data_out <= rom_array(2738);
		when "0000101010110011" => data_out <= rom_array(2739);
		when "0000101010110100" => data_out <= rom_array(2740);
		when "0000101010110101" => data_out <= rom_array(2741);
		when "0000101010110110" => data_out <= rom_array(2742);
		when "0000101010110111" => data_out <= rom_array(2743);
		when "0000101010111000" => data_out <= rom_array(2744);
		when "0000101010111001" => data_out <= rom_array(2745);
		when "0000101010111010" => data_out <= rom_array(2746);
		when "0000101010111011" => data_out <= rom_array(2747);
		when "0000101010111100" => data_out <= rom_array(2748);
		when "0000101010111101" => data_out <= rom_array(2749);
		when "0000101010111110" => data_out <= rom_array(2750);
		when "0000101010111111" => data_out <= rom_array(2751);
		when "0000101011000000" => data_out <= rom_array(2752);
		when "0000101011000001" => data_out <= rom_array(2753);
		when "0000101011000010" => data_out <= rom_array(2754);
		when "0000101011000011" => data_out <= rom_array(2755);
		when "0000101011000100" => data_out <= rom_array(2756);
		when "0000101011000101" => data_out <= rom_array(2757);
		when "0000101011000110" => data_out <= rom_array(2758);
		when "0000101011000111" => data_out <= rom_array(2759);
		when "0000101011001000" => data_out <= rom_array(2760);
		when "0000101011001001" => data_out <= rom_array(2761);
		when "0000101011001010" => data_out <= rom_array(2762);
		when "0000101011001011" => data_out <= rom_array(2763);
		when "0000101011001100" => data_out <= rom_array(2764);
		when "0000101011001101" => data_out <= rom_array(2765);
		when "0000101011001110" => data_out <= rom_array(2766);
		when "0000101011001111" => data_out <= rom_array(2767);
		when "0000101011010000" => data_out <= rom_array(2768);
		when "0000101011010001" => data_out <= rom_array(2769);
		when "0000101011010010" => data_out <= rom_array(2770);
		when "0000101011010011" => data_out <= rom_array(2771);
		when "0000101011010100" => data_out <= rom_array(2772);
		when "0000101011010101" => data_out <= rom_array(2773);
		when "0000101011010110" => data_out <= rom_array(2774);
		when "0000101011010111" => data_out <= rom_array(2775);
		when "0000101011011000" => data_out <= rom_array(2776);
		when "0000101011011001" => data_out <= rom_array(2777);
		when "0000101011011010" => data_out <= rom_array(2778);
		when "0000101011011011" => data_out <= rom_array(2779);
		when "0000101011011100" => data_out <= rom_array(2780);
		when "0000101011011101" => data_out <= rom_array(2781);
		when "0000101011011110" => data_out <= rom_array(2782);
		when "0000101011011111" => data_out <= rom_array(2783);
		when "0000101011100000" => data_out <= rom_array(2784);
		when "0000101011100001" => data_out <= rom_array(2785);
		when "0000101011100010" => data_out <= rom_array(2786);
		when "0000101011100011" => data_out <= rom_array(2787);
		when "0000101011100100" => data_out <= rom_array(2788);
		when "0000101011100101" => data_out <= rom_array(2789);
		when "0000101011100110" => data_out <= rom_array(2790);
		when "0000101011100111" => data_out <= rom_array(2791);
		when "0000101011101000" => data_out <= rom_array(2792);
		when "0000101011101001" => data_out <= rom_array(2793);
		when "0000101011101010" => data_out <= rom_array(2794);
		when "0000101011101011" => data_out <= rom_array(2795);
		when "0000101011101100" => data_out <= rom_array(2796);
		when "0000101011101101" => data_out <= rom_array(2797);
		when "0000101011101110" => data_out <= rom_array(2798);
		when "0000101011101111" => data_out <= rom_array(2799);
		when "0000101011110000" => data_out <= rom_array(2800);
		when "0000101011110001" => data_out <= rom_array(2801);
		when "0000101011110010" => data_out <= rom_array(2802);
		when "0000101011110011" => data_out <= rom_array(2803);
		when "0000101011110100" => data_out <= rom_array(2804);
		when "0000101011110101" => data_out <= rom_array(2805);
		when "0000101011110110" => data_out <= rom_array(2806);
		when "0000101011110111" => data_out <= rom_array(2807);
		when "0000101011111000" => data_out <= rom_array(2808);
		when "0000101011111001" => data_out <= rom_array(2809);
		when "0000101011111010" => data_out <= rom_array(2810);
		when "0000101011111011" => data_out <= rom_array(2811);
		when "0000101011111100" => data_out <= rom_array(2812);
		when "0000101011111101" => data_out <= rom_array(2813);
		when "0000101011111110" => data_out <= rom_array(2814);
		when "0000101011111111" => data_out <= rom_array(2815);
		when "0000101100000000" => data_out <= rom_array(2816);
		when "0000101100000001" => data_out <= rom_array(2817);
		when "0000101100000010" => data_out <= rom_array(2818);
		when "0000101100000011" => data_out <= rom_array(2819);
		when "0000101100000100" => data_out <= rom_array(2820);
		when "0000101100000101" => data_out <= rom_array(2821);
		when "0000101100000110" => data_out <= rom_array(2822);
		when "0000101100000111" => data_out <= rom_array(2823);
		when "0000101100001000" => data_out <= rom_array(2824);
		when "0000101100001001" => data_out <= rom_array(2825);
		when "0000101100001010" => data_out <= rom_array(2826);
		when "0000101100001011" => data_out <= rom_array(2827);
		when "0000101100001100" => data_out <= rom_array(2828);
		when "0000101100001101" => data_out <= rom_array(2829);
		when "0000101100001110" => data_out <= rom_array(2830);
		when "0000101100001111" => data_out <= rom_array(2831);
		when "0000101100010000" => data_out <= rom_array(2832);
		when "0000101100010001" => data_out <= rom_array(2833);
		when "0000101100010010" => data_out <= rom_array(2834);
		when "0000101100010011" => data_out <= rom_array(2835);
		when "0000101100010100" => data_out <= rom_array(2836);
		when "0000101100010101" => data_out <= rom_array(2837);
		when "0000101100010110" => data_out <= rom_array(2838);
		when "0000101100010111" => data_out <= rom_array(2839);
		when "0000101100011000" => data_out <= rom_array(2840);
		when "0000101100011001" => data_out <= rom_array(2841);
		when "0000101100011010" => data_out <= rom_array(2842);
		when "0000101100011011" => data_out <= rom_array(2843);
		when "0000101100011100" => data_out <= rom_array(2844);
		when "0000101100011101" => data_out <= rom_array(2845);
		when "0000101100011110" => data_out <= rom_array(2846);
		when "0000101100011111" => data_out <= rom_array(2847);
		when "0000101100100000" => data_out <= rom_array(2848);
		when "0000101100100001" => data_out <= rom_array(2849);
		when "0000101100100010" => data_out <= rom_array(2850);
		when "0000101100100011" => data_out <= rom_array(2851);
		when "0000101100100100" => data_out <= rom_array(2852);
		when "0000101100100101" => data_out <= rom_array(2853);
		when "0000101100100110" => data_out <= rom_array(2854);
		when "0000101100100111" => data_out <= rom_array(2855);
		when "0000101100101000" => data_out <= rom_array(2856);
		when "0000101100101001" => data_out <= rom_array(2857);
		when "0000101100101010" => data_out <= rom_array(2858);
		when "0000101100101011" => data_out <= rom_array(2859);
		when "0000101100101100" => data_out <= rom_array(2860);
		when "0000101100101101" => data_out <= rom_array(2861);
		when "0000101100101110" => data_out <= rom_array(2862);
		when "0000101100101111" => data_out <= rom_array(2863);
		when "0000101100110000" => data_out <= rom_array(2864);
		when "0000101100110001" => data_out <= rom_array(2865);
		when "0000101100110010" => data_out <= rom_array(2866);
		when "0000101100110011" => data_out <= rom_array(2867);
		when "0000101100110100" => data_out <= rom_array(2868);
		when "0000101100110101" => data_out <= rom_array(2869);
		when "0000101100110110" => data_out <= rom_array(2870);
		when "0000101100110111" => data_out <= rom_array(2871);
		when "0000101100111000" => data_out <= rom_array(2872);
		when "0000101100111001" => data_out <= rom_array(2873);
		when "0000101100111010" => data_out <= rom_array(2874);
		when "0000101100111011" => data_out <= rom_array(2875);
		when "0000101100111100" => data_out <= rom_array(2876);
		when "0000101100111101" => data_out <= rom_array(2877);
		when "0000101100111110" => data_out <= rom_array(2878);
		when "0000101100111111" => data_out <= rom_array(2879);
		when "0000101101000000" => data_out <= rom_array(2880);
		when "0000101101000001" => data_out <= rom_array(2881);
		when "0000101101000010" => data_out <= rom_array(2882);
		when "0000101101000011" => data_out <= rom_array(2883);
		when "0000101101000100" => data_out <= rom_array(2884);
		when "0000101101000101" => data_out <= rom_array(2885);
		when "0000101101000110" => data_out <= rom_array(2886);
		when "0000101101000111" => data_out <= rom_array(2887);
		when "0000101101001000" => data_out <= rom_array(2888);
		when "0000101101001001" => data_out <= rom_array(2889);
		when "0000101101001010" => data_out <= rom_array(2890);
		when "0000101101001011" => data_out <= rom_array(2891);
		when "0000101101001100" => data_out <= rom_array(2892);
		when "0000101101001101" => data_out <= rom_array(2893);
		when "0000101101001110" => data_out <= rom_array(2894);
		when "0000101101001111" => data_out <= rom_array(2895);
		when "0000101101010000" => data_out <= rom_array(2896);
		when "0000101101010001" => data_out <= rom_array(2897);
		when "0000101101010010" => data_out <= rom_array(2898);
		when "0000101101010011" => data_out <= rom_array(2899);
		when "0000101101010100" => data_out <= rom_array(2900);
		when "0000101101010101" => data_out <= rom_array(2901);
		when "0000101101010110" => data_out <= rom_array(2902);
		when "0000101101010111" => data_out <= rom_array(2903);
		when "0000101101011000" => data_out <= rom_array(2904);
		when "0000101101011001" => data_out <= rom_array(2905);
		when "0000101101011010" => data_out <= rom_array(2906);
		when "0000101101011011" => data_out <= rom_array(2907);
		when "0000101101011100" => data_out <= rom_array(2908);
		when "0000101101011101" => data_out <= rom_array(2909);
		when "0000101101011110" => data_out <= rom_array(2910);
		when "0000101101011111" => data_out <= rom_array(2911);
		when "0000101101100000" => data_out <= rom_array(2912);
		when "0000101101100001" => data_out <= rom_array(2913);
		when "0000101101100010" => data_out <= rom_array(2914);
		when "0000101101100011" => data_out <= rom_array(2915);
		when "0000101101100100" => data_out <= rom_array(2916);
		when "0000101101100101" => data_out <= rom_array(2917);
		when "0000101101100110" => data_out <= rom_array(2918);
		when "0000101101100111" => data_out <= rom_array(2919);
		when "0000101101101000" => data_out <= rom_array(2920);
		when "0000101101101001" => data_out <= rom_array(2921);
		when "0000101101101010" => data_out <= rom_array(2922);
		when "0000101101101011" => data_out <= rom_array(2923);
		when "0000101101101100" => data_out <= rom_array(2924);
		when "0000101101101101" => data_out <= rom_array(2925);
		when "0000101101101110" => data_out <= rom_array(2926);
		when "0000101101101111" => data_out <= rom_array(2927);
		when "0000101101110000" => data_out <= rom_array(2928);
		when "0000101101110001" => data_out <= rom_array(2929);
		when "0000101101110010" => data_out <= rom_array(2930);
		when "0000101101110011" => data_out <= rom_array(2931);
		when "0000101101110100" => data_out <= rom_array(2932);
		when "0000101101110101" => data_out <= rom_array(2933);
		when "0000101101110110" => data_out <= rom_array(2934);
		when "0000101101110111" => data_out <= rom_array(2935);
		when "0000101101111000" => data_out <= rom_array(2936);
		when "0000101101111001" => data_out <= rom_array(2937);
		when "0000101101111010" => data_out <= rom_array(2938);
		when "0000101101111011" => data_out <= rom_array(2939);
		when "0000101101111100" => data_out <= rom_array(2940);
		when "0000101101111101" => data_out <= rom_array(2941);
		when "0000101101111110" => data_out <= rom_array(2942);
		when "0000101101111111" => data_out <= rom_array(2943);
		when "0000101110000000" => data_out <= rom_array(2944);
		when "0000101110000001" => data_out <= rom_array(2945);
		when "0000101110000010" => data_out <= rom_array(2946);
		when "0000101110000011" => data_out <= rom_array(2947);
		when "0000101110000100" => data_out <= rom_array(2948);
		when "0000101110000101" => data_out <= rom_array(2949);
		when "0000101110000110" => data_out <= rom_array(2950);
		when "0000101110000111" => data_out <= rom_array(2951);
		when "0000101110001000" => data_out <= rom_array(2952);
		when "0000101110001001" => data_out <= rom_array(2953);
		when "0000101110001010" => data_out <= rom_array(2954);
		when "0000101110001011" => data_out <= rom_array(2955);
		when "0000101110001100" => data_out <= rom_array(2956);
		when "0000101110001101" => data_out <= rom_array(2957);
		when "0000101110001110" => data_out <= rom_array(2958);
		when "0000101110001111" => data_out <= rom_array(2959);
		when "0000101110010000" => data_out <= rom_array(2960);
		when "0000101110010001" => data_out <= rom_array(2961);
		when "0000101110010010" => data_out <= rom_array(2962);
		when "0000101110010011" => data_out <= rom_array(2963);
		when "0000101110010100" => data_out <= rom_array(2964);
		when "0000101110010101" => data_out <= rom_array(2965);
		when "0000101110010110" => data_out <= rom_array(2966);
		when "0000101110010111" => data_out <= rom_array(2967);
		when "0000101110011000" => data_out <= rom_array(2968);
		when "0000101110011001" => data_out <= rom_array(2969);
		when "0000101110011010" => data_out <= rom_array(2970);
		when "0000101110011011" => data_out <= rom_array(2971);
		when "0000101110011100" => data_out <= rom_array(2972);
		when "0000101110011101" => data_out <= rom_array(2973);
		when "0000101110011110" => data_out <= rom_array(2974);
		when "0000101110011111" => data_out <= rom_array(2975);
		when "0000101110100000" => data_out <= rom_array(2976);
		when "0000101110100001" => data_out <= rom_array(2977);
		when "0000101110100010" => data_out <= rom_array(2978);
		when "0000101110100011" => data_out <= rom_array(2979);
		when "0000101110100100" => data_out <= rom_array(2980);
		when "0000101110100101" => data_out <= rom_array(2981);
		when "0000101110100110" => data_out <= rom_array(2982);
		when "0000101110100111" => data_out <= rom_array(2983);
		when "0000101110101000" => data_out <= rom_array(2984);
		when "0000101110101001" => data_out <= rom_array(2985);
		when "0000101110101010" => data_out <= rom_array(2986);
		when "0000101110101011" => data_out <= rom_array(2987);
		when "0000101110101100" => data_out <= rom_array(2988);
		when "0000101110101101" => data_out <= rom_array(2989);
		when "0000101110101110" => data_out <= rom_array(2990);
		when "0000101110101111" => data_out <= rom_array(2991);
		when "0000101110110000" => data_out <= rom_array(2992);
		when "0000101110110001" => data_out <= rom_array(2993);
		when "0000101110110010" => data_out <= rom_array(2994);
		when "0000101110110011" => data_out <= rom_array(2995);
		when "0000101110110100" => data_out <= rom_array(2996);
		when "0000101110110101" => data_out <= rom_array(2997);
		when "0000101110110110" => data_out <= rom_array(2998);
		when "0000101110110111" => data_out <= rom_array(2999);
		when "0000101110111000" => data_out <= rom_array(3000);
		when "0000101110111001" => data_out <= rom_array(3001);
		when "0000101110111010" => data_out <= rom_array(3002);
		when "0000101110111011" => data_out <= rom_array(3003);
		when "0000101110111100" => data_out <= rom_array(3004);
		when "0000101110111101" => data_out <= rom_array(3005);
		when "0000101110111110" => data_out <= rom_array(3006);
		when "0000101110111111" => data_out <= rom_array(3007);
		when "0000101111000000" => data_out <= rom_array(3008);
		when "0000101111000001" => data_out <= rom_array(3009);
		when "0000101111000010" => data_out <= rom_array(3010);
		when "0000101111000011" => data_out <= rom_array(3011);
		when "0000101111000100" => data_out <= rom_array(3012);
		when "0000101111000101" => data_out <= rom_array(3013);
		when "0000101111000110" => data_out <= rom_array(3014);
		when "0000101111000111" => data_out <= rom_array(3015);
		when "0000101111001000" => data_out <= rom_array(3016);
		when "0000101111001001" => data_out <= rom_array(3017);
		when "0000101111001010" => data_out <= rom_array(3018);
		when "0000101111001011" => data_out <= rom_array(3019);
		when "0000101111001100" => data_out <= rom_array(3020);
		when "0000101111001101" => data_out <= rom_array(3021);
		when "0000101111001110" => data_out <= rom_array(3022);
		when "0000101111001111" => data_out <= rom_array(3023);
		when "0000101111010000" => data_out <= rom_array(3024);
		when "0000101111010001" => data_out <= rom_array(3025);
		when "0000101111010010" => data_out <= rom_array(3026);
		when "0000101111010011" => data_out <= rom_array(3027);
		when "0000101111010100" => data_out <= rom_array(3028);
		when "0000101111010101" => data_out <= rom_array(3029);
		when "0000101111010110" => data_out <= rom_array(3030);
		when "0000101111010111" => data_out <= rom_array(3031);
		when "0000101111011000" => data_out <= rom_array(3032);
		when "0000101111011001" => data_out <= rom_array(3033);
		when "0000101111011010" => data_out <= rom_array(3034);
		when "0000101111011011" => data_out <= rom_array(3035);
		when "0000101111011100" => data_out <= rom_array(3036);
		when "0000101111011101" => data_out <= rom_array(3037);
		when "0000101111011110" => data_out <= rom_array(3038);
		when "0000101111011111" => data_out <= rom_array(3039);
		when "0000101111100000" => data_out <= rom_array(3040);
		when "0000101111100001" => data_out <= rom_array(3041);
		when "0000101111100010" => data_out <= rom_array(3042);
		when "0000101111100011" => data_out <= rom_array(3043);
		when "0000101111100100" => data_out <= rom_array(3044);
		when "0000101111100101" => data_out <= rom_array(3045);
		when "0000101111100110" => data_out <= rom_array(3046);
		when "0000101111100111" => data_out <= rom_array(3047);
		when "0000101111101000" => data_out <= rom_array(3048);
		when "0000101111101001" => data_out <= rom_array(3049);
		when "0000101111101010" => data_out <= rom_array(3050);
		when "0000101111101011" => data_out <= rom_array(3051);
		when "0000101111101100" => data_out <= rom_array(3052);
		when "0000101111101101" => data_out <= rom_array(3053);
		when "0000101111101110" => data_out <= rom_array(3054);
		when "0000101111101111" => data_out <= rom_array(3055);
		when "0000101111110000" => data_out <= rom_array(3056);
		when "0000101111110001" => data_out <= rom_array(3057);
		when "0000101111110010" => data_out <= rom_array(3058);
		when "0000101111110011" => data_out <= rom_array(3059);
		when "0000101111110100" => data_out <= rom_array(3060);
		when "0000101111110101" => data_out <= rom_array(3061);
		when "0000101111110110" => data_out <= rom_array(3062);
		when "0000101111110111" => data_out <= rom_array(3063);
		when "0000101111111000" => data_out <= rom_array(3064);
		when "0000101111111001" => data_out <= rom_array(3065);
		when "0000101111111010" => data_out <= rom_array(3066);
		when "0000101111111011" => data_out <= rom_array(3067);
		when "0000101111111100" => data_out <= rom_array(3068);
		when "0000101111111101" => data_out <= rom_array(3069);
		when "0000101111111110" => data_out <= rom_array(3070);
		when "0000101111111111" => data_out <= rom_array(3071);
		when "0000110000000000" => data_out <= rom_array(3072);
		when "0000110000000001" => data_out <= rom_array(3073);
		when "0000110000000010" => data_out <= rom_array(3074);
		when "0000110000000011" => data_out <= rom_array(3075);
		when "0000110000000100" => data_out <= rom_array(3076);
		when "0000110000000101" => data_out <= rom_array(3077);
		when "0000110000000110" => data_out <= rom_array(3078);
		when "0000110000000111" => data_out <= rom_array(3079);
		when "0000110000001000" => data_out <= rom_array(3080);
		when "0000110000001001" => data_out <= rom_array(3081);
		when "0000110000001010" => data_out <= rom_array(3082);
		when "0000110000001011" => data_out <= rom_array(3083);
		when "0000110000001100" => data_out <= rom_array(3084);
		when "0000110000001101" => data_out <= rom_array(3085);
		when "0000110000001110" => data_out <= rom_array(3086);
		when "0000110000001111" => data_out <= rom_array(3087);
		when "0000110000010000" => data_out <= rom_array(3088);
		when "0000110000010001" => data_out <= rom_array(3089);
		when "0000110000010010" => data_out <= rom_array(3090);
		when "0000110000010011" => data_out <= rom_array(3091);
		when "0000110000010100" => data_out <= rom_array(3092);
		when "0000110000010101" => data_out <= rom_array(3093);
		when "0000110000010110" => data_out <= rom_array(3094);
		when "0000110000010111" => data_out <= rom_array(3095);
		when "0000110000011000" => data_out <= rom_array(3096);
		when "0000110000011001" => data_out <= rom_array(3097);
		when "0000110000011010" => data_out <= rom_array(3098);
		when "0000110000011011" => data_out <= rom_array(3099);
		when "0000110000011100" => data_out <= rom_array(3100);
		when "0000110000011101" => data_out <= rom_array(3101);
		when "0000110000011110" => data_out <= rom_array(3102);
		when "0000110000011111" => data_out <= rom_array(3103);
		when "0000110000100000" => data_out <= rom_array(3104);
		when "0000110000100001" => data_out <= rom_array(3105);
		when "0000110000100010" => data_out <= rom_array(3106);
		when "0000110000100011" => data_out <= rom_array(3107);
		when "0000110000100100" => data_out <= rom_array(3108);
		when "0000110000100101" => data_out <= rom_array(3109);
		when "0000110000100110" => data_out <= rom_array(3110);
		when "0000110000100111" => data_out <= rom_array(3111);
		when "0000110000101000" => data_out <= rom_array(3112);
		when "0000110000101001" => data_out <= rom_array(3113);
		when "0000110000101010" => data_out <= rom_array(3114);
		when "0000110000101011" => data_out <= rom_array(3115);
		when "0000110000101100" => data_out <= rom_array(3116);
		when "0000110000101101" => data_out <= rom_array(3117);
		when "0000110000101110" => data_out <= rom_array(3118);
		when "0000110000101111" => data_out <= rom_array(3119);
		when "0000110000110000" => data_out <= rom_array(3120);
		when "0000110000110001" => data_out <= rom_array(3121);
		when "0000110000110010" => data_out <= rom_array(3122);
		when "0000110000110011" => data_out <= rom_array(3123);
		when "0000110000110100" => data_out <= rom_array(3124);
		when "0000110000110101" => data_out <= rom_array(3125);
		when "0000110000110110" => data_out <= rom_array(3126);
		when "0000110000110111" => data_out <= rom_array(3127);
		when "0000110000111000" => data_out <= rom_array(3128);
		when "0000110000111001" => data_out <= rom_array(3129);
		when "0000110000111010" => data_out <= rom_array(3130);
		when "0000110000111011" => data_out <= rom_array(3131);
		when "0000110000111100" => data_out <= rom_array(3132);
		when "0000110000111101" => data_out <= rom_array(3133);
		when "0000110000111110" => data_out <= rom_array(3134);
		when "0000110000111111" => data_out <= rom_array(3135);
		when "0000110001000000" => data_out <= rom_array(3136);
		when "0000110001000001" => data_out <= rom_array(3137);
		when "0000110001000010" => data_out <= rom_array(3138);
		when "0000110001000011" => data_out <= rom_array(3139);
		when "0000110001000100" => data_out <= rom_array(3140);
		when "0000110001000101" => data_out <= rom_array(3141);
		when "0000110001000110" => data_out <= rom_array(3142);
		when "0000110001000111" => data_out <= rom_array(3143);
		when "0000110001001000" => data_out <= rom_array(3144);
		when "0000110001001001" => data_out <= rom_array(3145);
		when "0000110001001010" => data_out <= rom_array(3146);
		when "0000110001001011" => data_out <= rom_array(3147);
		when "0000110001001100" => data_out <= rom_array(3148);
		when "0000110001001101" => data_out <= rom_array(3149);
		when "0000110001001110" => data_out <= rom_array(3150);
		when "0000110001001111" => data_out <= rom_array(3151);
		when "0000110001010000" => data_out <= rom_array(3152);
		when "0000110001010001" => data_out <= rom_array(3153);
		when "0000110001010010" => data_out <= rom_array(3154);
		when "0000110001010011" => data_out <= rom_array(3155);
		when "0000110001010100" => data_out <= rom_array(3156);
		when "0000110001010101" => data_out <= rom_array(3157);
		when "0000110001010110" => data_out <= rom_array(3158);
		when "0000110001010111" => data_out <= rom_array(3159);
		when "0000110001011000" => data_out <= rom_array(3160);
		when "0000110001011001" => data_out <= rom_array(3161);
		when "0000110001011010" => data_out <= rom_array(3162);
		when "0000110001011011" => data_out <= rom_array(3163);
		when "0000110001011100" => data_out <= rom_array(3164);
		when "0000110001011101" => data_out <= rom_array(3165);
		when "0000110001011110" => data_out <= rom_array(3166);
		when "0000110001011111" => data_out <= rom_array(3167);
		when "0000110001100000" => data_out <= rom_array(3168);
		when "0000110001100001" => data_out <= rom_array(3169);
		when "0000110001100010" => data_out <= rom_array(3170);
		when "0000110001100011" => data_out <= rom_array(3171);
		when "0000110001100100" => data_out <= rom_array(3172);
		when "0000110001100101" => data_out <= rom_array(3173);
		when "0000110001100110" => data_out <= rom_array(3174);
		when "0000110001100111" => data_out <= rom_array(3175);
		when "0000110001101000" => data_out <= rom_array(3176);
		when "0000110001101001" => data_out <= rom_array(3177);
		when "0000110001101010" => data_out <= rom_array(3178);
		when "0000110001101011" => data_out <= rom_array(3179);
		when "0000110001101100" => data_out <= rom_array(3180);
		when "0000110001101101" => data_out <= rom_array(3181);
		when "0000110001101110" => data_out <= rom_array(3182);
		when "0000110001101111" => data_out <= rom_array(3183);
		when "0000110001110000" => data_out <= rom_array(3184);
		when "0000110001110001" => data_out <= rom_array(3185);
		when "0000110001110010" => data_out <= rom_array(3186);
		when "0000110001110011" => data_out <= rom_array(3187);
		when "0000110001110100" => data_out <= rom_array(3188);
		when "0000110001110101" => data_out <= rom_array(3189);
		when "0000110001110110" => data_out <= rom_array(3190);
		when "0000110001110111" => data_out <= rom_array(3191);
		when "0000110001111000" => data_out <= rom_array(3192);
		when "0000110001111001" => data_out <= rom_array(3193);
		when "0000110001111010" => data_out <= rom_array(3194);
		when "0000110001111011" => data_out <= rom_array(3195);
		when "0000110001111100" => data_out <= rom_array(3196);
		when "0000110001111101" => data_out <= rom_array(3197);
		when "0000110001111110" => data_out <= rom_array(3198);
		when "0000110001111111" => data_out <= rom_array(3199);
		when "0000110010000000" => data_out <= rom_array(3200);
		when "0000110010000001" => data_out <= rom_array(3201);
		when "0000110010000010" => data_out <= rom_array(3202);
		when "0000110010000011" => data_out <= rom_array(3203);
		when "0000110010000100" => data_out <= rom_array(3204);
		when "0000110010000101" => data_out <= rom_array(3205);
		when "0000110010000110" => data_out <= rom_array(3206);
		when "0000110010000111" => data_out <= rom_array(3207);
		when "0000110010001000" => data_out <= rom_array(3208);
		when "0000110010001001" => data_out <= rom_array(3209);
		when "0000110010001010" => data_out <= rom_array(3210);
		when "0000110010001011" => data_out <= rom_array(3211);
		when "0000110010001100" => data_out <= rom_array(3212);
		when "0000110010001101" => data_out <= rom_array(3213);
		when "0000110010001110" => data_out <= rom_array(3214);
		when "0000110010001111" => data_out <= rom_array(3215);
		when "0000110010010000" => data_out <= rom_array(3216);
		when "0000110010010001" => data_out <= rom_array(3217);
		when "0000110010010010" => data_out <= rom_array(3218);
		when "0000110010010011" => data_out <= rom_array(3219);
		when "0000110010010100" => data_out <= rom_array(3220);
		when "0000110010010101" => data_out <= rom_array(3221);
		when "0000110010010110" => data_out <= rom_array(3222);
		when "0000110010010111" => data_out <= rom_array(3223);
		when "0000110010011000" => data_out <= rom_array(3224);
		when "0000110010011001" => data_out <= rom_array(3225);
		when "0000110010011010" => data_out <= rom_array(3226);
		when "0000110010011011" => data_out <= rom_array(3227);
		when "0000110010011100" => data_out <= rom_array(3228);
		when "0000110010011101" => data_out <= rom_array(3229);
		when "0000110010011110" => data_out <= rom_array(3230);
		when "0000110010011111" => data_out <= rom_array(3231);
		when "0000110010100000" => data_out <= rom_array(3232);
		when "0000110010100001" => data_out <= rom_array(3233);
		when "0000110010100010" => data_out <= rom_array(3234);
		when "0000110010100011" => data_out <= rom_array(3235);
		when "0000110010100100" => data_out <= rom_array(3236);
		when "0000110010100101" => data_out <= rom_array(3237);
		when "0000110010100110" => data_out <= rom_array(3238);
		when "0000110010100111" => data_out <= rom_array(3239);
		when "0000110010101000" => data_out <= rom_array(3240);
		when "0000110010101001" => data_out <= rom_array(3241);
		when "0000110010101010" => data_out <= rom_array(3242);
		when "0000110010101011" => data_out <= rom_array(3243);
		when "0000110010101100" => data_out <= rom_array(3244);
		when "0000110010101101" => data_out <= rom_array(3245);
		when "0000110010101110" => data_out <= rom_array(3246);
		when "0000110010101111" => data_out <= rom_array(3247);
		when "0000110010110000" => data_out <= rom_array(3248);
		when "0000110010110001" => data_out <= rom_array(3249);
		when "0000110010110010" => data_out <= rom_array(3250);
		when "0000110010110011" => data_out <= rom_array(3251);
		when "0000110010110100" => data_out <= rom_array(3252);
		when "0000110010110101" => data_out <= rom_array(3253);
		when "0000110010110110" => data_out <= rom_array(3254);
		when "0000110010110111" => data_out <= rom_array(3255);
		when "0000110010111000" => data_out <= rom_array(3256);
		when "0000110010111001" => data_out <= rom_array(3257);
		when "0000110010111010" => data_out <= rom_array(3258);
		when "0000110010111011" => data_out <= rom_array(3259);
		when "0000110010111100" => data_out <= rom_array(3260);
		when "0000110010111101" => data_out <= rom_array(3261);
		when "0000110010111110" => data_out <= rom_array(3262);
		when "0000110010111111" => data_out <= rom_array(3263);
		when "0000110011000000" => data_out <= rom_array(3264);
		when "0000110011000001" => data_out <= rom_array(3265);
		when "0000110011000010" => data_out <= rom_array(3266);
		when "0000110011000011" => data_out <= rom_array(3267);
		when "0000110011000100" => data_out <= rom_array(3268);
		when "0000110011000101" => data_out <= rom_array(3269);
		when "0000110011000110" => data_out <= rom_array(3270);
		when "0000110011000111" => data_out <= rom_array(3271);
		when "0000110011001000" => data_out <= rom_array(3272);
		when "0000110011001001" => data_out <= rom_array(3273);
		when "0000110011001010" => data_out <= rom_array(3274);
		when "0000110011001011" => data_out <= rom_array(3275);
		when "0000110011001100" => data_out <= rom_array(3276);
		when "0000110011001101" => data_out <= rom_array(3277);
		when "0000110011001110" => data_out <= rom_array(3278);
		when "0000110011001111" => data_out <= rom_array(3279);
		when "0000110011010000" => data_out <= rom_array(3280);
		when "0000110011010001" => data_out <= rom_array(3281);
		when "0000110011010010" => data_out <= rom_array(3282);
		when "0000110011010011" => data_out <= rom_array(3283);
		when "0000110011010100" => data_out <= rom_array(3284);
		when "0000110011010101" => data_out <= rom_array(3285);
		when "0000110011010110" => data_out <= rom_array(3286);
		when "0000110011010111" => data_out <= rom_array(3287);
		when "0000110011011000" => data_out <= rom_array(3288);
		when "0000110011011001" => data_out <= rom_array(3289);
		when "0000110011011010" => data_out <= rom_array(3290);
		when "0000110011011011" => data_out <= rom_array(3291);
		when "0000110011011100" => data_out <= rom_array(3292);
		when "0000110011011101" => data_out <= rom_array(3293);
		when "0000110011011110" => data_out <= rom_array(3294);
		when "0000110011011111" => data_out <= rom_array(3295);
		when "0000110011100000" => data_out <= rom_array(3296);
		when "0000110011100001" => data_out <= rom_array(3297);
		when "0000110011100010" => data_out <= rom_array(3298);
		when "0000110011100011" => data_out <= rom_array(3299);
		when "0000110011100100" => data_out <= rom_array(3300);
		when "0000110011100101" => data_out <= rom_array(3301);
		when "0000110011100110" => data_out <= rom_array(3302);
		when "0000110011100111" => data_out <= rom_array(3303);
		when "0000110011101000" => data_out <= rom_array(3304);
		when "0000110011101001" => data_out <= rom_array(3305);
		when "0000110011101010" => data_out <= rom_array(3306);
		when "0000110011101011" => data_out <= rom_array(3307);
		when "0000110011101100" => data_out <= rom_array(3308);
		when "0000110011101101" => data_out <= rom_array(3309);
		when "0000110011101110" => data_out <= rom_array(3310);
		when "0000110011101111" => data_out <= rom_array(3311);
		when "0000110011110000" => data_out <= rom_array(3312);
		when "0000110011110001" => data_out <= rom_array(3313);
		when "0000110011110010" => data_out <= rom_array(3314);
		when "0000110011110011" => data_out <= rom_array(3315);
		when "0000110011110100" => data_out <= rom_array(3316);
		when "0000110011110101" => data_out <= rom_array(3317);
		when "0000110011110110" => data_out <= rom_array(3318);
		when "0000110011110111" => data_out <= rom_array(3319);
		when "0000110011111000" => data_out <= rom_array(3320);
		when "0000110011111001" => data_out <= rom_array(3321);
		when "0000110011111010" => data_out <= rom_array(3322);
		when "0000110011111011" => data_out <= rom_array(3323);
		when "0000110011111100" => data_out <= rom_array(3324);
		when "0000110011111101" => data_out <= rom_array(3325);
		when "0000110011111110" => data_out <= rom_array(3326);
		when "0000110011111111" => data_out <= rom_array(3327);
		when "0000110100000000" => data_out <= rom_array(3328);
		when "0000110100000001" => data_out <= rom_array(3329);
		when "0000110100000010" => data_out <= rom_array(3330);
		when "0000110100000011" => data_out <= rom_array(3331);
		when "0000110100000100" => data_out <= rom_array(3332);
		when "0000110100000101" => data_out <= rom_array(3333);
		when "0000110100000110" => data_out <= rom_array(3334);
		when "0000110100000111" => data_out <= rom_array(3335);
		when "0000110100001000" => data_out <= rom_array(3336);
		when "0000110100001001" => data_out <= rom_array(3337);
		when "0000110100001010" => data_out <= rom_array(3338);
		when "0000110100001011" => data_out <= rom_array(3339);
		when "0000110100001100" => data_out <= rom_array(3340);
		when "0000110100001101" => data_out <= rom_array(3341);
		when "0000110100001110" => data_out <= rom_array(3342);
		when "0000110100001111" => data_out <= rom_array(3343);
		when "0000110100010000" => data_out <= rom_array(3344);
		when "0000110100010001" => data_out <= rom_array(3345);
		when "0000110100010010" => data_out <= rom_array(3346);
		when "0000110100010011" => data_out <= rom_array(3347);
		when "0000110100010100" => data_out <= rom_array(3348);
		when "0000110100010101" => data_out <= rom_array(3349);
		when "0000110100010110" => data_out <= rom_array(3350);
		when "0000110100010111" => data_out <= rom_array(3351);
		when "0000110100011000" => data_out <= rom_array(3352);
		when "0000110100011001" => data_out <= rom_array(3353);
		when "0000110100011010" => data_out <= rom_array(3354);
		when "0000110100011011" => data_out <= rom_array(3355);
		when "0000110100011100" => data_out <= rom_array(3356);
		when "0000110100011101" => data_out <= rom_array(3357);
		when "0000110100011110" => data_out <= rom_array(3358);
		when "0000110100011111" => data_out <= rom_array(3359);
		when "0000110100100000" => data_out <= rom_array(3360);
		when "0000110100100001" => data_out <= rom_array(3361);
		when "0000110100100010" => data_out <= rom_array(3362);
		when "0000110100100011" => data_out <= rom_array(3363);
		when "0000110100100100" => data_out <= rom_array(3364);
		when "0000110100100101" => data_out <= rom_array(3365);
		when "0000110100100110" => data_out <= rom_array(3366);
		when "0000110100100111" => data_out <= rom_array(3367);
		when "0000110100101000" => data_out <= rom_array(3368);
		when "0000110100101001" => data_out <= rom_array(3369);
		when "0000110100101010" => data_out <= rom_array(3370);
		when "0000110100101011" => data_out <= rom_array(3371);
		when "0000110100101100" => data_out <= rom_array(3372);
		when "0000110100101101" => data_out <= rom_array(3373);
		when "0000110100101110" => data_out <= rom_array(3374);
		when "0000110100101111" => data_out <= rom_array(3375);
		when "0000110100110000" => data_out <= rom_array(3376);
		when "0000110100110001" => data_out <= rom_array(3377);
		when "0000110100110010" => data_out <= rom_array(3378);
		when "0000110100110011" => data_out <= rom_array(3379);
		when "0000110100110100" => data_out <= rom_array(3380);
		when "0000110100110101" => data_out <= rom_array(3381);
		when "0000110100110110" => data_out <= rom_array(3382);
		when "0000110100110111" => data_out <= rom_array(3383);
		when "0000110100111000" => data_out <= rom_array(3384);
		when "0000110100111001" => data_out <= rom_array(3385);
		when "0000110100111010" => data_out <= rom_array(3386);
		when "0000110100111011" => data_out <= rom_array(3387);
		when "0000110100111100" => data_out <= rom_array(3388);
		when "0000110100111101" => data_out <= rom_array(3389);
		when "0000110100111110" => data_out <= rom_array(3390);
		when "0000110100111111" => data_out <= rom_array(3391);
		when "0000110101000000" => data_out <= rom_array(3392);
		when "0000110101000001" => data_out <= rom_array(3393);
		when "0000110101000010" => data_out <= rom_array(3394);
		when "0000110101000011" => data_out <= rom_array(3395);
		when "0000110101000100" => data_out <= rom_array(3396);
		when "0000110101000101" => data_out <= rom_array(3397);
		when "0000110101000110" => data_out <= rom_array(3398);
		when "0000110101000111" => data_out <= rom_array(3399);
		when "0000110101001000" => data_out <= rom_array(3400);
		when "0000110101001001" => data_out <= rom_array(3401);
		when "0000110101001010" => data_out <= rom_array(3402);
		when "0000110101001011" => data_out <= rom_array(3403);
		when "0000110101001100" => data_out <= rom_array(3404);
		when "0000110101001101" => data_out <= rom_array(3405);
		when "0000110101001110" => data_out <= rom_array(3406);
		when "0000110101001111" => data_out <= rom_array(3407);
		when "0000110101010000" => data_out <= rom_array(3408);
		when "0000110101010001" => data_out <= rom_array(3409);
		when "0000110101010010" => data_out <= rom_array(3410);
		when "0000110101010011" => data_out <= rom_array(3411);
		when "0000110101010100" => data_out <= rom_array(3412);
		when "0000110101010101" => data_out <= rom_array(3413);
		when "0000110101010110" => data_out <= rom_array(3414);
		when "0000110101010111" => data_out <= rom_array(3415);
		when "0000110101011000" => data_out <= rom_array(3416);
		when "0000110101011001" => data_out <= rom_array(3417);
		when "0000110101011010" => data_out <= rom_array(3418);
		when "0000110101011011" => data_out <= rom_array(3419);
		when "0000110101011100" => data_out <= rom_array(3420);
		when "0000110101011101" => data_out <= rom_array(3421);
		when "0000110101011110" => data_out <= rom_array(3422);
		when "0000110101011111" => data_out <= rom_array(3423);
		when "0000110101100000" => data_out <= rom_array(3424);
		when "0000110101100001" => data_out <= rom_array(3425);
		when "0000110101100010" => data_out <= rom_array(3426);
		when "0000110101100011" => data_out <= rom_array(3427);
		when "0000110101100100" => data_out <= rom_array(3428);
		when "0000110101100101" => data_out <= rom_array(3429);
		when "0000110101100110" => data_out <= rom_array(3430);
		when "0000110101100111" => data_out <= rom_array(3431);
		when "0000110101101000" => data_out <= rom_array(3432);
		when "0000110101101001" => data_out <= rom_array(3433);
		when "0000110101101010" => data_out <= rom_array(3434);
		when "0000110101101011" => data_out <= rom_array(3435);
		when "0000110101101100" => data_out <= rom_array(3436);
		when "0000110101101101" => data_out <= rom_array(3437);
		when "0000110101101110" => data_out <= rom_array(3438);
		when "0000110101101111" => data_out <= rom_array(3439);
		when "0000110101110000" => data_out <= rom_array(3440);
		when "0000110101110001" => data_out <= rom_array(3441);
		when "0000110101110010" => data_out <= rom_array(3442);
		when "0000110101110011" => data_out <= rom_array(3443);
		when "0000110101110100" => data_out <= rom_array(3444);
		when "0000110101110101" => data_out <= rom_array(3445);
		when "0000110101110110" => data_out <= rom_array(3446);
		when "0000110101110111" => data_out <= rom_array(3447);
		when "0000110101111000" => data_out <= rom_array(3448);
		when "0000110101111001" => data_out <= rom_array(3449);
		when "0000110101111010" => data_out <= rom_array(3450);
		when "0000110101111011" => data_out <= rom_array(3451);
		when "0000110101111100" => data_out <= rom_array(3452);
		when "0000110101111101" => data_out <= rom_array(3453);
		when "0000110101111110" => data_out <= rom_array(3454);
		when "0000110101111111" => data_out <= rom_array(3455);
		when "0000110110000000" => data_out <= rom_array(3456);
		when "0000110110000001" => data_out <= rom_array(3457);
		when "0000110110000010" => data_out <= rom_array(3458);
		when "0000110110000011" => data_out <= rom_array(3459);
		when "0000110110000100" => data_out <= rom_array(3460);
		when "0000110110000101" => data_out <= rom_array(3461);
		when "0000110110000110" => data_out <= rom_array(3462);
		when "0000110110000111" => data_out <= rom_array(3463);
		when "0000110110001000" => data_out <= rom_array(3464);
		when "0000110110001001" => data_out <= rom_array(3465);
		when "0000110110001010" => data_out <= rom_array(3466);
		when "0000110110001011" => data_out <= rom_array(3467);
		when "0000110110001100" => data_out <= rom_array(3468);
		when "0000110110001101" => data_out <= rom_array(3469);
		when "0000110110001110" => data_out <= rom_array(3470);
		when "0000110110001111" => data_out <= rom_array(3471);
		when "0000110110010000" => data_out <= rom_array(3472);
		when "0000110110010001" => data_out <= rom_array(3473);
		when "0000110110010010" => data_out <= rom_array(3474);
		when "0000110110010011" => data_out <= rom_array(3475);
		when "0000110110010100" => data_out <= rom_array(3476);
		when "0000110110010101" => data_out <= rom_array(3477);
		when "0000110110010110" => data_out <= rom_array(3478);
		when "0000110110010111" => data_out <= rom_array(3479);
		when "0000110110011000" => data_out <= rom_array(3480);
		when "0000110110011001" => data_out <= rom_array(3481);
		when "0000110110011010" => data_out <= rom_array(3482);
		when "0000110110011011" => data_out <= rom_array(3483);
		when "0000110110011100" => data_out <= rom_array(3484);
		when "0000110110011101" => data_out <= rom_array(3485);
		when "0000110110011110" => data_out <= rom_array(3486);
		when "0000110110011111" => data_out <= rom_array(3487);
		when "0000110110100000" => data_out <= rom_array(3488);
		when "0000110110100001" => data_out <= rom_array(3489);
		when "0000110110100010" => data_out <= rom_array(3490);
		when "0000110110100011" => data_out <= rom_array(3491);
		when "0000110110100100" => data_out <= rom_array(3492);
		when "0000110110100101" => data_out <= rom_array(3493);
		when "0000110110100110" => data_out <= rom_array(3494);
		when "0000110110100111" => data_out <= rom_array(3495);
		when "0000110110101000" => data_out <= rom_array(3496);
		when "0000110110101001" => data_out <= rom_array(3497);
		when "0000110110101010" => data_out <= rom_array(3498);
		when "0000110110101011" => data_out <= rom_array(3499);
		when "0000110110101100" => data_out <= rom_array(3500);
		when "0000110110101101" => data_out <= rom_array(3501);
		when "0000110110101110" => data_out <= rom_array(3502);
		when "0000110110101111" => data_out <= rom_array(3503);
		when "0000110110110000" => data_out <= rom_array(3504);
		when "0000110110110001" => data_out <= rom_array(3505);
		when "0000110110110010" => data_out <= rom_array(3506);
		when "0000110110110011" => data_out <= rom_array(3507);
		when "0000110110110100" => data_out <= rom_array(3508);
		when "0000110110110101" => data_out <= rom_array(3509);
		when "0000110110110110" => data_out <= rom_array(3510);
		when "0000110110110111" => data_out <= rom_array(3511);
		when "0000110110111000" => data_out <= rom_array(3512);
		when "0000110110111001" => data_out <= rom_array(3513);
		when "0000110110111010" => data_out <= rom_array(3514);
		when "0000110110111011" => data_out <= rom_array(3515);
		when "0000110110111100" => data_out <= rom_array(3516);
		when "0000110110111101" => data_out <= rom_array(3517);
		when "0000110110111110" => data_out <= rom_array(3518);
		when "0000110110111111" => data_out <= rom_array(3519);
		when "0000110111000000" => data_out <= rom_array(3520);
		when "0000110111000001" => data_out <= rom_array(3521);
		when "0000110111000010" => data_out <= rom_array(3522);
		when "0000110111000011" => data_out <= rom_array(3523);
		when "0000110111000100" => data_out <= rom_array(3524);
		when "0000110111000101" => data_out <= rom_array(3525);
		when "0000110111000110" => data_out <= rom_array(3526);
		when "0000110111000111" => data_out <= rom_array(3527);
		when "0000110111001000" => data_out <= rom_array(3528);
		when "0000110111001001" => data_out <= rom_array(3529);
		when "0000110111001010" => data_out <= rom_array(3530);
		when "0000110111001011" => data_out <= rom_array(3531);
		when "0000110111001100" => data_out <= rom_array(3532);
		when "0000110111001101" => data_out <= rom_array(3533);
		when "0000110111001110" => data_out <= rom_array(3534);
		when "0000110111001111" => data_out <= rom_array(3535);
		when "0000110111010000" => data_out <= rom_array(3536);
		when "0000110111010001" => data_out <= rom_array(3537);
		when "0000110111010010" => data_out <= rom_array(3538);
		when "0000110111010011" => data_out <= rom_array(3539);
		when "0000110111010100" => data_out <= rom_array(3540);
		when "0000110111010101" => data_out <= rom_array(3541);
		when "0000110111010110" => data_out <= rom_array(3542);
		when "0000110111010111" => data_out <= rom_array(3543);
		when "0000110111011000" => data_out <= rom_array(3544);
		when "0000110111011001" => data_out <= rom_array(3545);
		when "0000110111011010" => data_out <= rom_array(3546);
		when "0000110111011011" => data_out <= rom_array(3547);
		when "0000110111011100" => data_out <= rom_array(3548);
		when "0000110111011101" => data_out <= rom_array(3549);
		when "0000110111011110" => data_out <= rom_array(3550);
		when "0000110111011111" => data_out <= rom_array(3551);
		when "0000110111100000" => data_out <= rom_array(3552);
		when "0000110111100001" => data_out <= rom_array(3553);
		when "0000110111100010" => data_out <= rom_array(3554);
		when "0000110111100011" => data_out <= rom_array(3555);
		when "0000110111100100" => data_out <= rom_array(3556);
		when "0000110111100101" => data_out <= rom_array(3557);
		when "0000110111100110" => data_out <= rom_array(3558);
		when "0000110111100111" => data_out <= rom_array(3559);
		when "0000110111101000" => data_out <= rom_array(3560);
		when "0000110111101001" => data_out <= rom_array(3561);
		when "0000110111101010" => data_out <= rom_array(3562);
		when "0000110111101011" => data_out <= rom_array(3563);
		when "0000110111101100" => data_out <= rom_array(3564);
		when "0000110111101101" => data_out <= rom_array(3565);
		when "0000110111101110" => data_out <= rom_array(3566);
		when "0000110111101111" => data_out <= rom_array(3567);
		when "0000110111110000" => data_out <= rom_array(3568);
		when "0000110111110001" => data_out <= rom_array(3569);
		when "0000110111110010" => data_out <= rom_array(3570);
		when "0000110111110011" => data_out <= rom_array(3571);
		when "0000110111110100" => data_out <= rom_array(3572);
		when "0000110111110101" => data_out <= rom_array(3573);
		when "0000110111110110" => data_out <= rom_array(3574);
		when "0000110111110111" => data_out <= rom_array(3575);
		when "0000110111111000" => data_out <= rom_array(3576);
		when "0000110111111001" => data_out <= rom_array(3577);
		when "0000110111111010" => data_out <= rom_array(3578);
		when "0000110111111011" => data_out <= rom_array(3579);
		when "0000110111111100" => data_out <= rom_array(3580);
		when "0000110111111101" => data_out <= rom_array(3581);
		when "0000110111111110" => data_out <= rom_array(3582);
		when "0000110111111111" => data_out <= rom_array(3583);
		when "0000111000000000" => data_out <= rom_array(3584);
		when "0000111000000001" => data_out <= rom_array(3585);
		when "0000111000000010" => data_out <= rom_array(3586);
		when "0000111000000011" => data_out <= rom_array(3587);
		when "0000111000000100" => data_out <= rom_array(3588);
		when "0000111000000101" => data_out <= rom_array(3589);
		when "0000111000000110" => data_out <= rom_array(3590);
		when "0000111000000111" => data_out <= rom_array(3591);
		when "0000111000001000" => data_out <= rom_array(3592);
		when "0000111000001001" => data_out <= rom_array(3593);
		when "0000111000001010" => data_out <= rom_array(3594);
		when "0000111000001011" => data_out <= rom_array(3595);
		when "0000111000001100" => data_out <= rom_array(3596);
		when "0000111000001101" => data_out <= rom_array(3597);
		when "0000111000001110" => data_out <= rom_array(3598);
		when "0000111000001111" => data_out <= rom_array(3599);
		when "0000111000010000" => data_out <= rom_array(3600);
		when "0000111000010001" => data_out <= rom_array(3601);
		when "0000111000010010" => data_out <= rom_array(3602);
		when "0000111000010011" => data_out <= rom_array(3603);
		when "0000111000010100" => data_out <= rom_array(3604);
		when "0000111000010101" => data_out <= rom_array(3605);
		when "0000111000010110" => data_out <= rom_array(3606);
		when "0000111000010111" => data_out <= rom_array(3607);
		when "0000111000011000" => data_out <= rom_array(3608);
		when "0000111000011001" => data_out <= rom_array(3609);
		when "0000111000011010" => data_out <= rom_array(3610);
		when "0000111000011011" => data_out <= rom_array(3611);
		when "0000111000011100" => data_out <= rom_array(3612);
		when "0000111000011101" => data_out <= rom_array(3613);
		when "0000111000011110" => data_out <= rom_array(3614);
		when "0000111000011111" => data_out <= rom_array(3615);
		when "0000111000100000" => data_out <= rom_array(3616);
		when "0000111000100001" => data_out <= rom_array(3617);
		when "0000111000100010" => data_out <= rom_array(3618);
		when "0000111000100011" => data_out <= rom_array(3619);
		when "0000111000100100" => data_out <= rom_array(3620);
		when "0000111000100101" => data_out <= rom_array(3621);
		when "0000111000100110" => data_out <= rom_array(3622);
		when "0000111000100111" => data_out <= rom_array(3623);
		when "0000111000101000" => data_out <= rom_array(3624);
		when "0000111000101001" => data_out <= rom_array(3625);
		when "0000111000101010" => data_out <= rom_array(3626);
		when "0000111000101011" => data_out <= rom_array(3627);
		when "0000111000101100" => data_out <= rom_array(3628);
		when "0000111000101101" => data_out <= rom_array(3629);
		when "0000111000101110" => data_out <= rom_array(3630);
		when "0000111000101111" => data_out <= rom_array(3631);
		when "0000111000110000" => data_out <= rom_array(3632);
		when "0000111000110001" => data_out <= rom_array(3633);
		when "0000111000110010" => data_out <= rom_array(3634);
		when "0000111000110011" => data_out <= rom_array(3635);
		when "0000111000110100" => data_out <= rom_array(3636);
		when "0000111000110101" => data_out <= rom_array(3637);
		when "0000111000110110" => data_out <= rom_array(3638);
		when "0000111000110111" => data_out <= rom_array(3639);
		when "0000111000111000" => data_out <= rom_array(3640);
		when "0000111000111001" => data_out <= rom_array(3641);
		when "0000111000111010" => data_out <= rom_array(3642);
		when "0000111000111011" => data_out <= rom_array(3643);
		when "0000111000111100" => data_out <= rom_array(3644);
		when "0000111000111101" => data_out <= rom_array(3645);
		when "0000111000111110" => data_out <= rom_array(3646);
		when "0000111000111111" => data_out <= rom_array(3647);
		when "0000111001000000" => data_out <= rom_array(3648);
		when "0000111001000001" => data_out <= rom_array(3649);
		when "0000111001000010" => data_out <= rom_array(3650);
		when "0000111001000011" => data_out <= rom_array(3651);
		when "0000111001000100" => data_out <= rom_array(3652);
		when "0000111001000101" => data_out <= rom_array(3653);
		when "0000111001000110" => data_out <= rom_array(3654);
		when "0000111001000111" => data_out <= rom_array(3655);
		when "0000111001001000" => data_out <= rom_array(3656);
		when "0000111001001001" => data_out <= rom_array(3657);
		when "0000111001001010" => data_out <= rom_array(3658);
		when "0000111001001011" => data_out <= rom_array(3659);
		when "0000111001001100" => data_out <= rom_array(3660);
		when "0000111001001101" => data_out <= rom_array(3661);
		when "0000111001001110" => data_out <= rom_array(3662);
		when "0000111001001111" => data_out <= rom_array(3663);
		when "0000111001010000" => data_out <= rom_array(3664);
		when "0000111001010001" => data_out <= rom_array(3665);
		when "0000111001010010" => data_out <= rom_array(3666);
		when "0000111001010011" => data_out <= rom_array(3667);
		when "0000111001010100" => data_out <= rom_array(3668);
		when "0000111001010101" => data_out <= rom_array(3669);
		when "0000111001010110" => data_out <= rom_array(3670);
		when "0000111001010111" => data_out <= rom_array(3671);
		when "0000111001011000" => data_out <= rom_array(3672);
		when "0000111001011001" => data_out <= rom_array(3673);
		when "0000111001011010" => data_out <= rom_array(3674);
		when "0000111001011011" => data_out <= rom_array(3675);
		when "0000111001011100" => data_out <= rom_array(3676);
		when "0000111001011101" => data_out <= rom_array(3677);
		when "0000111001011110" => data_out <= rom_array(3678);
		when "0000111001011111" => data_out <= rom_array(3679);
		when "0000111001100000" => data_out <= rom_array(3680);
		when "0000111001100001" => data_out <= rom_array(3681);
		when "0000111001100010" => data_out <= rom_array(3682);
		when "0000111001100011" => data_out <= rom_array(3683);
		when "0000111001100100" => data_out <= rom_array(3684);
		when "0000111001100101" => data_out <= rom_array(3685);
		when "0000111001100110" => data_out <= rom_array(3686);
		when "0000111001100111" => data_out <= rom_array(3687);
		when "0000111001101000" => data_out <= rom_array(3688);
		when "0000111001101001" => data_out <= rom_array(3689);
		when "0000111001101010" => data_out <= rom_array(3690);
		when "0000111001101011" => data_out <= rom_array(3691);
		when "0000111001101100" => data_out <= rom_array(3692);
		when "0000111001101101" => data_out <= rom_array(3693);
		when "0000111001101110" => data_out <= rom_array(3694);
		when "0000111001101111" => data_out <= rom_array(3695);
		when "0000111001110000" => data_out <= rom_array(3696);
		when "0000111001110001" => data_out <= rom_array(3697);
		when "0000111001110010" => data_out <= rom_array(3698);
		when "0000111001110011" => data_out <= rom_array(3699);
		when "0000111001110100" => data_out <= rom_array(3700);
		when "0000111001110101" => data_out <= rom_array(3701);
		when "0000111001110110" => data_out <= rom_array(3702);
		when "0000111001110111" => data_out <= rom_array(3703);
		when "0000111001111000" => data_out <= rom_array(3704);
		when "0000111001111001" => data_out <= rom_array(3705);
		when "0000111001111010" => data_out <= rom_array(3706);
		when "0000111001111011" => data_out <= rom_array(3707);
		when "0000111001111100" => data_out <= rom_array(3708);
		when "0000111001111101" => data_out <= rom_array(3709);
		when "0000111001111110" => data_out <= rom_array(3710);
		when "0000111001111111" => data_out <= rom_array(3711);
		when "0000111010000000" => data_out <= rom_array(3712);
		when "0000111010000001" => data_out <= rom_array(3713);
		when "0000111010000010" => data_out <= rom_array(3714);
		when "0000111010000011" => data_out <= rom_array(3715);
		when "0000111010000100" => data_out <= rom_array(3716);
		when "0000111010000101" => data_out <= rom_array(3717);
		when "0000111010000110" => data_out <= rom_array(3718);
		when "0000111010000111" => data_out <= rom_array(3719);
		when "0000111010001000" => data_out <= rom_array(3720);
		when "0000111010001001" => data_out <= rom_array(3721);
		when "0000111010001010" => data_out <= rom_array(3722);
		when "0000111010001011" => data_out <= rom_array(3723);
		when "0000111010001100" => data_out <= rom_array(3724);
		when "0000111010001101" => data_out <= rom_array(3725);
		when "0000111010001110" => data_out <= rom_array(3726);
		when "0000111010001111" => data_out <= rom_array(3727);
		when "0000111010010000" => data_out <= rom_array(3728);
		when "0000111010010001" => data_out <= rom_array(3729);
		when "0000111010010010" => data_out <= rom_array(3730);
		when "0000111010010011" => data_out <= rom_array(3731);
		when "0000111010010100" => data_out <= rom_array(3732);
		when "0000111010010101" => data_out <= rom_array(3733);
		when "0000111010010110" => data_out <= rom_array(3734);
		when "0000111010010111" => data_out <= rom_array(3735);
		when "0000111010011000" => data_out <= rom_array(3736);
		when "0000111010011001" => data_out <= rom_array(3737);
		when "0000111010011010" => data_out <= rom_array(3738);
		when "0000111010011011" => data_out <= rom_array(3739);
		when "0000111010011100" => data_out <= rom_array(3740);
		when "0000111010011101" => data_out <= rom_array(3741);
		when "0000111010011110" => data_out <= rom_array(3742);
		when "0000111010011111" => data_out <= rom_array(3743);
		when "0000111010100000" => data_out <= rom_array(3744);
		when "0000111010100001" => data_out <= rom_array(3745);
		when "0000111010100010" => data_out <= rom_array(3746);
		when "0000111010100011" => data_out <= rom_array(3747);
		when "0000111010100100" => data_out <= rom_array(3748);
		when "0000111010100101" => data_out <= rom_array(3749);
		when "0000111010100110" => data_out <= rom_array(3750);
		when "0000111010100111" => data_out <= rom_array(3751);
		when "0000111010101000" => data_out <= rom_array(3752);
		when "0000111010101001" => data_out <= rom_array(3753);
		when "0000111010101010" => data_out <= rom_array(3754);
		when "0000111010101011" => data_out <= rom_array(3755);
		when "0000111010101100" => data_out <= rom_array(3756);
		when "0000111010101101" => data_out <= rom_array(3757);
		when "0000111010101110" => data_out <= rom_array(3758);
		when "0000111010101111" => data_out <= rom_array(3759);
		when "0000111010110000" => data_out <= rom_array(3760);
		when "0000111010110001" => data_out <= rom_array(3761);
		when "0000111010110010" => data_out <= rom_array(3762);
		when "0000111010110011" => data_out <= rom_array(3763);
		when "0000111010110100" => data_out <= rom_array(3764);
		when "0000111010110101" => data_out <= rom_array(3765);
		when "0000111010110110" => data_out <= rom_array(3766);
		when "0000111010110111" => data_out <= rom_array(3767);
		when "0000111010111000" => data_out <= rom_array(3768);
		when "0000111010111001" => data_out <= rom_array(3769);
		when "0000111010111010" => data_out <= rom_array(3770);
		when "0000111010111011" => data_out <= rom_array(3771);
		when "0000111010111100" => data_out <= rom_array(3772);
		when "0000111010111101" => data_out <= rom_array(3773);
		when "0000111010111110" => data_out <= rom_array(3774);
		when "0000111010111111" => data_out <= rom_array(3775);
		when "0000111011000000" => data_out <= rom_array(3776);
		when "0000111011000001" => data_out <= rom_array(3777);
		when "0000111011000010" => data_out <= rom_array(3778);
		when "0000111011000011" => data_out <= rom_array(3779);
		when "0000111011000100" => data_out <= rom_array(3780);
		when "0000111011000101" => data_out <= rom_array(3781);
		when "0000111011000110" => data_out <= rom_array(3782);
		when "0000111011000111" => data_out <= rom_array(3783);
		when "0000111011001000" => data_out <= rom_array(3784);
		when "0000111011001001" => data_out <= rom_array(3785);
		when "0000111011001010" => data_out <= rom_array(3786);
		when "0000111011001011" => data_out <= rom_array(3787);
		when "0000111011001100" => data_out <= rom_array(3788);
		when "0000111011001101" => data_out <= rom_array(3789);
		when "0000111011001110" => data_out <= rom_array(3790);
		when "0000111011001111" => data_out <= rom_array(3791);
		when "0000111011010000" => data_out <= rom_array(3792);
		when "0000111011010001" => data_out <= rom_array(3793);
		when "0000111011010010" => data_out <= rom_array(3794);
		when "0000111011010011" => data_out <= rom_array(3795);
		when "0000111011010100" => data_out <= rom_array(3796);
		when "0000111011010101" => data_out <= rom_array(3797);
		when "0000111011010110" => data_out <= rom_array(3798);
		when "0000111011010111" => data_out <= rom_array(3799);
		when "0000111011011000" => data_out <= rom_array(3800);
		when "0000111011011001" => data_out <= rom_array(3801);
		when "0000111011011010" => data_out <= rom_array(3802);
		when "0000111011011011" => data_out <= rom_array(3803);
		when "0000111011011100" => data_out <= rom_array(3804);
		when "0000111011011101" => data_out <= rom_array(3805);
		when "0000111011011110" => data_out <= rom_array(3806);
		when "0000111011011111" => data_out <= rom_array(3807);
		when "0000111011100000" => data_out <= rom_array(3808);
		when "0000111011100001" => data_out <= rom_array(3809);
		when "0000111011100010" => data_out <= rom_array(3810);
		when "0000111011100011" => data_out <= rom_array(3811);
		when "0000111011100100" => data_out <= rom_array(3812);
		when "0000111011100101" => data_out <= rom_array(3813);
		when "0000111011100110" => data_out <= rom_array(3814);
		when "0000111011100111" => data_out <= rom_array(3815);
		when "0000111011101000" => data_out <= rom_array(3816);
		when "0000111011101001" => data_out <= rom_array(3817);
		when "0000111011101010" => data_out <= rom_array(3818);
		when "0000111011101011" => data_out <= rom_array(3819);
		when "0000111011101100" => data_out <= rom_array(3820);
		when "0000111011101101" => data_out <= rom_array(3821);
		when "0000111011101110" => data_out <= rom_array(3822);
		when "0000111011101111" => data_out <= rom_array(3823);
		when "0000111011110000" => data_out <= rom_array(3824);
		when "0000111011110001" => data_out <= rom_array(3825);
		when "0000111011110010" => data_out <= rom_array(3826);
		when "0000111011110011" => data_out <= rom_array(3827);
		when "0000111011110100" => data_out <= rom_array(3828);
		when "0000111011110101" => data_out <= rom_array(3829);
		when "0000111011110110" => data_out <= rom_array(3830);
		when "0000111011110111" => data_out <= rom_array(3831);
		when "0000111011111000" => data_out <= rom_array(3832);
		when "0000111011111001" => data_out <= rom_array(3833);
		when "0000111011111010" => data_out <= rom_array(3834);
		when "0000111011111011" => data_out <= rom_array(3835);
		when "0000111011111100" => data_out <= rom_array(3836);
		when "0000111011111101" => data_out <= rom_array(3837);
		when "0000111011111110" => data_out <= rom_array(3838);
		when "0000111011111111" => data_out <= rom_array(3839);
		when "0000111100000000" => data_out <= rom_array(3840);
		when "0000111100000001" => data_out <= rom_array(3841);
		when "0000111100000010" => data_out <= rom_array(3842);
		when "0000111100000011" => data_out <= rom_array(3843);
		when "0000111100000100" => data_out <= rom_array(3844);
		when "0000111100000101" => data_out <= rom_array(3845);
		when "0000111100000110" => data_out <= rom_array(3846);
		when "0000111100000111" => data_out <= rom_array(3847);
		when "0000111100001000" => data_out <= rom_array(3848);
		when "0000111100001001" => data_out <= rom_array(3849);
		when "0000111100001010" => data_out <= rom_array(3850);
		when "0000111100001011" => data_out <= rom_array(3851);
		when "0000111100001100" => data_out <= rom_array(3852);
		when "0000111100001101" => data_out <= rom_array(3853);
		when "0000111100001110" => data_out <= rom_array(3854);
		when "0000111100001111" => data_out <= rom_array(3855);
		when "0000111100010000" => data_out <= rom_array(3856);
		when "0000111100010001" => data_out <= rom_array(3857);
		when "0000111100010010" => data_out <= rom_array(3858);
		when "0000111100010011" => data_out <= rom_array(3859);
		when "0000111100010100" => data_out <= rom_array(3860);
		when "0000111100010101" => data_out <= rom_array(3861);
		when "0000111100010110" => data_out <= rom_array(3862);
		when "0000111100010111" => data_out <= rom_array(3863);
		when "0000111100011000" => data_out <= rom_array(3864);
		when "0000111100011001" => data_out <= rom_array(3865);
		when "0000111100011010" => data_out <= rom_array(3866);
		when "0000111100011011" => data_out <= rom_array(3867);
		when "0000111100011100" => data_out <= rom_array(3868);
		when "0000111100011101" => data_out <= rom_array(3869);
		when "0000111100011110" => data_out <= rom_array(3870);
		when "0000111100011111" => data_out <= rom_array(3871);
		when "0000111100100000" => data_out <= rom_array(3872);
		when "0000111100100001" => data_out <= rom_array(3873);
		when "0000111100100010" => data_out <= rom_array(3874);
		when "0000111100100011" => data_out <= rom_array(3875);
		when "0000111100100100" => data_out <= rom_array(3876);
		when "0000111100100101" => data_out <= rom_array(3877);
		when "0000111100100110" => data_out <= rom_array(3878);
		when "0000111100100111" => data_out <= rom_array(3879);
		when "0000111100101000" => data_out <= rom_array(3880);
		when "0000111100101001" => data_out <= rom_array(3881);
		when "0000111100101010" => data_out <= rom_array(3882);
		when "0000111100101011" => data_out <= rom_array(3883);
		when "0000111100101100" => data_out <= rom_array(3884);
		when "0000111100101101" => data_out <= rom_array(3885);
		when "0000111100101110" => data_out <= rom_array(3886);
		when "0000111100101111" => data_out <= rom_array(3887);
		when "0000111100110000" => data_out <= rom_array(3888);
		when "0000111100110001" => data_out <= rom_array(3889);
		when "0000111100110010" => data_out <= rom_array(3890);
		when "0000111100110011" => data_out <= rom_array(3891);
		when "0000111100110100" => data_out <= rom_array(3892);
		when "0000111100110101" => data_out <= rom_array(3893);
		when "0000111100110110" => data_out <= rom_array(3894);
		when "0000111100110111" => data_out <= rom_array(3895);
		when "0000111100111000" => data_out <= rom_array(3896);
		when "0000111100111001" => data_out <= rom_array(3897);
		when "0000111100111010" => data_out <= rom_array(3898);
		when "0000111100111011" => data_out <= rom_array(3899);
		when "0000111100111100" => data_out <= rom_array(3900);
		when "0000111100111101" => data_out <= rom_array(3901);
		when "0000111100111110" => data_out <= rom_array(3902);
		when "0000111100111111" => data_out <= rom_array(3903);
		when "0000111101000000" => data_out <= rom_array(3904);
		when "0000111101000001" => data_out <= rom_array(3905);
		when "0000111101000010" => data_out <= rom_array(3906);
		when "0000111101000011" => data_out <= rom_array(3907);
		when "0000111101000100" => data_out <= rom_array(3908);
		when "0000111101000101" => data_out <= rom_array(3909);
		when "0000111101000110" => data_out <= rom_array(3910);
		when "0000111101000111" => data_out <= rom_array(3911);
		when "0000111101001000" => data_out <= rom_array(3912);
		when "0000111101001001" => data_out <= rom_array(3913);
		when "0000111101001010" => data_out <= rom_array(3914);
		when "0000111101001011" => data_out <= rom_array(3915);
		when "0000111101001100" => data_out <= rom_array(3916);
		when "0000111101001101" => data_out <= rom_array(3917);
		when "0000111101001110" => data_out <= rom_array(3918);
		when "0000111101001111" => data_out <= rom_array(3919);
		when "0000111101010000" => data_out <= rom_array(3920);
		when "0000111101010001" => data_out <= rom_array(3921);
		when "0000111101010010" => data_out <= rom_array(3922);
		when "0000111101010011" => data_out <= rom_array(3923);
		when "0000111101010100" => data_out <= rom_array(3924);
		when "0000111101010101" => data_out <= rom_array(3925);
		when "0000111101010110" => data_out <= rom_array(3926);
		when "0000111101010111" => data_out <= rom_array(3927);
		when "0000111101011000" => data_out <= rom_array(3928);
		when "0000111101011001" => data_out <= rom_array(3929);
		when "0000111101011010" => data_out <= rom_array(3930);
		when "0000111101011011" => data_out <= rom_array(3931);
		when "0000111101011100" => data_out <= rom_array(3932);
		when "0000111101011101" => data_out <= rom_array(3933);
		when "0000111101011110" => data_out <= rom_array(3934);
		when "0000111101011111" => data_out <= rom_array(3935);
		when "0000111101100000" => data_out <= rom_array(3936);
		when "0000111101100001" => data_out <= rom_array(3937);
		when "0000111101100010" => data_out <= rom_array(3938);
		when "0000111101100011" => data_out <= rom_array(3939);
		when "0000111101100100" => data_out <= rom_array(3940);
		when "0000111101100101" => data_out <= rom_array(3941);
		when "0000111101100110" => data_out <= rom_array(3942);
		when "0000111101100111" => data_out <= rom_array(3943);
		when "0000111101101000" => data_out <= rom_array(3944);
		when "0000111101101001" => data_out <= rom_array(3945);
		when "0000111101101010" => data_out <= rom_array(3946);
		when "0000111101101011" => data_out <= rom_array(3947);
		when "0000111101101100" => data_out <= rom_array(3948);
		when "0000111101101101" => data_out <= rom_array(3949);
		when "0000111101101110" => data_out <= rom_array(3950);
		when "0000111101101111" => data_out <= rom_array(3951);
		when "0000111101110000" => data_out <= rom_array(3952);
		when "0000111101110001" => data_out <= rom_array(3953);
		when "0000111101110010" => data_out <= rom_array(3954);
		when "0000111101110011" => data_out <= rom_array(3955);
		when "0000111101110100" => data_out <= rom_array(3956);
		when "0000111101110101" => data_out <= rom_array(3957);
		when "0000111101110110" => data_out <= rom_array(3958);
		when "0000111101110111" => data_out <= rom_array(3959);
		when "0000111101111000" => data_out <= rom_array(3960);
		when "0000111101111001" => data_out <= rom_array(3961);
		when "0000111101111010" => data_out <= rom_array(3962);
		when "0000111101111011" => data_out <= rom_array(3963);
		when "0000111101111100" => data_out <= rom_array(3964);
		when "0000111101111101" => data_out <= rom_array(3965);
		when "0000111101111110" => data_out <= rom_array(3966);
		when "0000111101111111" => data_out <= rom_array(3967);
		when "0000111110000000" => data_out <= rom_array(3968);
		when "0000111110000001" => data_out <= rom_array(3969);
		when "0000111110000010" => data_out <= rom_array(3970);
		when "0000111110000011" => data_out <= rom_array(3971);
		when "0000111110000100" => data_out <= rom_array(3972);
		when "0000111110000101" => data_out <= rom_array(3973);
		when "0000111110000110" => data_out <= rom_array(3974);
		when "0000111110000111" => data_out <= rom_array(3975);
		when "0000111110001000" => data_out <= rom_array(3976);
		when "0000111110001001" => data_out <= rom_array(3977);
		when "0000111110001010" => data_out <= rom_array(3978);
		when "0000111110001011" => data_out <= rom_array(3979);
		when "0000111110001100" => data_out <= rom_array(3980);
		when "0000111110001101" => data_out <= rom_array(3981);
		when "0000111110001110" => data_out <= rom_array(3982);
		when "0000111110001111" => data_out <= rom_array(3983);
		when "0000111110010000" => data_out <= rom_array(3984);
		when "0000111110010001" => data_out <= rom_array(3985);
		when "0000111110010010" => data_out <= rom_array(3986);
		when "0000111110010011" => data_out <= rom_array(3987);
		when "0000111110010100" => data_out <= rom_array(3988);
		when "0000111110010101" => data_out <= rom_array(3989);
		when "0000111110010110" => data_out <= rom_array(3990);
		when "0000111110010111" => data_out <= rom_array(3991);
		when "0000111110011000" => data_out <= rom_array(3992);
		when "0000111110011001" => data_out <= rom_array(3993);
		when "0000111110011010" => data_out <= rom_array(3994);
		when "0000111110011011" => data_out <= rom_array(3995);
		when "0000111110011100" => data_out <= rom_array(3996);
		when "0000111110011101" => data_out <= rom_array(3997);
		when "0000111110011110" => data_out <= rom_array(3998);
		when "0000111110011111" => data_out <= rom_array(3999);
		when "0000111110100000" => data_out <= rom_array(4000);
		when "0000111110100001" => data_out <= rom_array(4001);
		when "0000111110100010" => data_out <= rom_array(4002);
		when "0000111110100011" => data_out <= rom_array(4003);
		when "0000111110100100" => data_out <= rom_array(4004);
		when "0000111110100101" => data_out <= rom_array(4005);
		when "0000111110100110" => data_out <= rom_array(4006);
		when "0000111110100111" => data_out <= rom_array(4007);
		when "0000111110101000" => data_out <= rom_array(4008);
		when "0000111110101001" => data_out <= rom_array(4009);
		when "0000111110101010" => data_out <= rom_array(4010);
		when "0000111110101011" => data_out <= rom_array(4011);
		when "0000111110101100" => data_out <= rom_array(4012);
		when "0000111110101101" => data_out <= rom_array(4013);
		when "0000111110101110" => data_out <= rom_array(4014);
		when "0000111110101111" => data_out <= rom_array(4015);
		when "0000111110110000" => data_out <= rom_array(4016);
		when "0000111110110001" => data_out <= rom_array(4017);
		when "0000111110110010" => data_out <= rom_array(4018);
		when "0000111110110011" => data_out <= rom_array(4019);
		when "0000111110110100" => data_out <= rom_array(4020);
		when "0000111110110101" => data_out <= rom_array(4021);
		when "0000111110110110" => data_out <= rom_array(4022);
		when "0000111110110111" => data_out <= rom_array(4023);
		when "0000111110111000" => data_out <= rom_array(4024);
		when "0000111110111001" => data_out <= rom_array(4025);
		when "0000111110111010" => data_out <= rom_array(4026);
		when "0000111110111011" => data_out <= rom_array(4027);
		when "0000111110111100" => data_out <= rom_array(4028);
		when "0000111110111101" => data_out <= rom_array(4029);
		when "0000111110111110" => data_out <= rom_array(4030);
		when "0000111110111111" => data_out <= rom_array(4031);
		when "0000111111000000" => data_out <= rom_array(4032);
		when "0000111111000001" => data_out <= rom_array(4033);
		when "0000111111000010" => data_out <= rom_array(4034);
		when "0000111111000011" => data_out <= rom_array(4035);
		when "0000111111000100" => data_out <= rom_array(4036);
		when "0000111111000101" => data_out <= rom_array(4037);
		when "0000111111000110" => data_out <= rom_array(4038);
		when "0000111111000111" => data_out <= rom_array(4039);
		when "0000111111001000" => data_out <= rom_array(4040);
		when "0000111111001001" => data_out <= rom_array(4041);
		when "0000111111001010" => data_out <= rom_array(4042);
		when "0000111111001011" => data_out <= rom_array(4043);
		when "0000111111001100" => data_out <= rom_array(4044);
		when "0000111111001101" => data_out <= rom_array(4045);
		when "0000111111001110" => data_out <= rom_array(4046);
		when "0000111111001111" => data_out <= rom_array(4047);
		when "0000111111010000" => data_out <= rom_array(4048);
		when "0000111111010001" => data_out <= rom_array(4049);
		when "0000111111010010" => data_out <= rom_array(4050);
		when "0000111111010011" => data_out <= rom_array(4051);
		when "0000111111010100" => data_out <= rom_array(4052);
		when "0000111111010101" => data_out <= rom_array(4053);
		when "0000111111010110" => data_out <= rom_array(4054);
		when "0000111111010111" => data_out <= rom_array(4055);
		when "0000111111011000" => data_out <= rom_array(4056);
		when "0000111111011001" => data_out <= rom_array(4057);
		when "0000111111011010" => data_out <= rom_array(4058);
		when "0000111111011011" => data_out <= rom_array(4059);
		when "0000111111011100" => data_out <= rom_array(4060);
		when "0000111111011101" => data_out <= rom_array(4061);
		when "0000111111011110" => data_out <= rom_array(4062);
		when "0000111111011111" => data_out <= rom_array(4063);
		when "0000111111100000" => data_out <= rom_array(4064);
		when "0000111111100001" => data_out <= rom_array(4065);
		when "0000111111100010" => data_out <= rom_array(4066);
		when "0000111111100011" => data_out <= rom_array(4067);
		when "0000111111100100" => data_out <= rom_array(4068);
		when "0000111111100101" => data_out <= rom_array(4069);
		when "0000111111100110" => data_out <= rom_array(4070);
		when "0000111111100111" => data_out <= rom_array(4071);
		when "0000111111101000" => data_out <= rom_array(4072);
		when "0000111111101001" => data_out <= rom_array(4073);
		when "0000111111101010" => data_out <= rom_array(4074);
		when "0000111111101011" => data_out <= rom_array(4075);
		when "0000111111101100" => data_out <= rom_array(4076);
		when "0000111111101101" => data_out <= rom_array(4077);
		when "0000111111101110" => data_out <= rom_array(4078);
		when "0000111111101111" => data_out <= rom_array(4079);
		when "0000111111110000" => data_out <= rom_array(4080);
		when "0000111111110001" => data_out <= rom_array(4081);
		when "0000111111110010" => data_out <= rom_array(4082);
		when "0000111111110011" => data_out <= rom_array(4083);
		when "0000111111110100" => data_out <= rom_array(4084);
		when "0000111111110101" => data_out <= rom_array(4085);
		when "0000111111110110" => data_out <= rom_array(4086);
		when "0000111111110111" => data_out <= rom_array(4087);
		when "0000111111111000" => data_out <= rom_array(4088);
		when "0000111111111001" => data_out <= rom_array(4089);
		when "0000111111111010" => data_out <= rom_array(4090);
		when "0000111111111011" => data_out <= rom_array(4091);
		when "0000111111111100" => data_out <= rom_array(4092);
		when "0000111111111101" => data_out <= rom_array(4093);
		when "0000111111111110" => data_out <= rom_array(4094);
		when "0000111111111111" => data_out <= rom_array(4095);
		when "0001000000000000" => data_out <= rom_array(4096);
		when "0001000000000001" => data_out <= rom_array(4097);
		when "0001000000000010" => data_out <= rom_array(4098);
		when "0001000000000011" => data_out <= rom_array(4099);
		when "0001000000000100" => data_out <= rom_array(4100);
		when "0001000000000101" => data_out <= rom_array(4101);
		when "0001000000000110" => data_out <= rom_array(4102);
		when "0001000000000111" => data_out <= rom_array(4103);
		when "0001000000001000" => data_out <= rom_array(4104);
		when "0001000000001001" => data_out <= rom_array(4105);
		when "0001000000001010" => data_out <= rom_array(4106);
		when "0001000000001011" => data_out <= rom_array(4107);
		when "0001000000001100" => data_out <= rom_array(4108);
		when "0001000000001101" => data_out <= rom_array(4109);
		when "0001000000001110" => data_out <= rom_array(4110);
		when "0001000000001111" => data_out <= rom_array(4111);
		when "0001000000010000" => data_out <= rom_array(4112);
		when "0001000000010001" => data_out <= rom_array(4113);
		when "0001000000010010" => data_out <= rom_array(4114);
		when "0001000000010011" => data_out <= rom_array(4115);
		when "0001000000010100" => data_out <= rom_array(4116);
		when "0001000000010101" => data_out <= rom_array(4117);
		when "0001000000010110" => data_out <= rom_array(4118);
		when "0001000000010111" => data_out <= rom_array(4119);
		when "0001000000011000" => data_out <= rom_array(4120);
		when "0001000000011001" => data_out <= rom_array(4121);
		when "0001000000011010" => data_out <= rom_array(4122);
		when "0001000000011011" => data_out <= rom_array(4123);
		when "0001000000011100" => data_out <= rom_array(4124);
		when "0001000000011101" => data_out <= rom_array(4125);
		when "0001000000011110" => data_out <= rom_array(4126);
		when "0001000000011111" => data_out <= rom_array(4127);
		when "0001000000100000" => data_out <= rom_array(4128);
		when "0001000000100001" => data_out <= rom_array(4129);
		when "0001000000100010" => data_out <= rom_array(4130);
		when "0001000000100011" => data_out <= rom_array(4131);
		when "0001000000100100" => data_out <= rom_array(4132);
		when "0001000000100101" => data_out <= rom_array(4133);
		when "0001000000100110" => data_out <= rom_array(4134);
		when "0001000000100111" => data_out <= rom_array(4135);
		when "0001000000101000" => data_out <= rom_array(4136);
		when "0001000000101001" => data_out <= rom_array(4137);
		when "0001000000101010" => data_out <= rom_array(4138);
		when "0001000000101011" => data_out <= rom_array(4139);
		when "0001000000101100" => data_out <= rom_array(4140);
		when "0001000000101101" => data_out <= rom_array(4141);
		when "0001000000101110" => data_out <= rom_array(4142);
		when "0001000000101111" => data_out <= rom_array(4143);
		when "0001000000110000" => data_out <= rom_array(4144);
		when "0001000000110001" => data_out <= rom_array(4145);
		when "0001000000110010" => data_out <= rom_array(4146);
		when "0001000000110011" => data_out <= rom_array(4147);
		when "0001000000110100" => data_out <= rom_array(4148);
		when "0001000000110101" => data_out <= rom_array(4149);
		when "0001000000110110" => data_out <= rom_array(4150);
		when "0001000000110111" => data_out <= rom_array(4151);
		when "0001000000111000" => data_out <= rom_array(4152);
		when "0001000000111001" => data_out <= rom_array(4153);
		when "0001000000111010" => data_out <= rom_array(4154);
		when "0001000000111011" => data_out <= rom_array(4155);
		when "0001000000111100" => data_out <= rom_array(4156);
		when "0001000000111101" => data_out <= rom_array(4157);
		when "0001000000111110" => data_out <= rom_array(4158);
		when "0001000000111111" => data_out <= rom_array(4159);
		when "0001000001000000" => data_out <= rom_array(4160);
		when "0001000001000001" => data_out <= rom_array(4161);
		when "0001000001000010" => data_out <= rom_array(4162);
		when "0001000001000011" => data_out <= rom_array(4163);
		when "0001000001000100" => data_out <= rom_array(4164);
		when "0001000001000101" => data_out <= rom_array(4165);
		when "0001000001000110" => data_out <= rom_array(4166);
		when "0001000001000111" => data_out <= rom_array(4167);
		when "0001000001001000" => data_out <= rom_array(4168);
		when "0001000001001001" => data_out <= rom_array(4169);
		when "0001000001001010" => data_out <= rom_array(4170);
		when "0001000001001011" => data_out <= rom_array(4171);
		when "0001000001001100" => data_out <= rom_array(4172);
		when "0001000001001101" => data_out <= rom_array(4173);
		when "0001000001001110" => data_out <= rom_array(4174);
		when "0001000001001111" => data_out <= rom_array(4175);
		when "0001000001010000" => data_out <= rom_array(4176);
		when "0001000001010001" => data_out <= rom_array(4177);
		when "0001000001010010" => data_out <= rom_array(4178);
		when "0001000001010011" => data_out <= rom_array(4179);
		when "0001000001010100" => data_out <= rom_array(4180);
		when "0001000001010101" => data_out <= rom_array(4181);
		when "0001000001010110" => data_out <= rom_array(4182);
		when "0001000001010111" => data_out <= rom_array(4183);
		when "0001000001011000" => data_out <= rom_array(4184);
		when "0001000001011001" => data_out <= rom_array(4185);
		when "0001000001011010" => data_out <= rom_array(4186);
		when "0001000001011011" => data_out <= rom_array(4187);
		when "0001000001011100" => data_out <= rom_array(4188);
		when "0001000001011101" => data_out <= rom_array(4189);
		when "0001000001011110" => data_out <= rom_array(4190);
		when "0001000001011111" => data_out <= rom_array(4191);
		when "0001000001100000" => data_out <= rom_array(4192);
		when "0001000001100001" => data_out <= rom_array(4193);
		when "0001000001100010" => data_out <= rom_array(4194);
		when "0001000001100011" => data_out <= rom_array(4195);
		when "0001000001100100" => data_out <= rom_array(4196);
		when "0001000001100101" => data_out <= rom_array(4197);
		when "0001000001100110" => data_out <= rom_array(4198);
		when "0001000001100111" => data_out <= rom_array(4199);
		when "0001000001101000" => data_out <= rom_array(4200);
		when "0001000001101001" => data_out <= rom_array(4201);
		when "0001000001101010" => data_out <= rom_array(4202);
		when "0001000001101011" => data_out <= rom_array(4203);
		when "0001000001101100" => data_out <= rom_array(4204);
		when "0001000001101101" => data_out <= rom_array(4205);
		when "0001000001101110" => data_out <= rom_array(4206);
		when "0001000001101111" => data_out <= rom_array(4207);
		when "0001000001110000" => data_out <= rom_array(4208);
		when "0001000001110001" => data_out <= rom_array(4209);
		when "0001000001110010" => data_out <= rom_array(4210);
		when "0001000001110011" => data_out <= rom_array(4211);
		when "0001000001110100" => data_out <= rom_array(4212);
		when "0001000001110101" => data_out <= rom_array(4213);
		when "0001000001110110" => data_out <= rom_array(4214);
		when "0001000001110111" => data_out <= rom_array(4215);
		when "0001000001111000" => data_out <= rom_array(4216);
		when "0001000001111001" => data_out <= rom_array(4217);
		when "0001000001111010" => data_out <= rom_array(4218);
		when "0001000001111011" => data_out <= rom_array(4219);
		when "0001000001111100" => data_out <= rom_array(4220);
		when "0001000001111101" => data_out <= rom_array(4221);
		when "0001000001111110" => data_out <= rom_array(4222);
		when "0001000001111111" => data_out <= rom_array(4223);
		when "0001000010000000" => data_out <= rom_array(4224);
		when "0001000010000001" => data_out <= rom_array(4225);
		when "0001000010000010" => data_out <= rom_array(4226);
		when "0001000010000011" => data_out <= rom_array(4227);
		when "0001000010000100" => data_out <= rom_array(4228);
		when "0001000010000101" => data_out <= rom_array(4229);
		when "0001000010000110" => data_out <= rom_array(4230);
		when "0001000010000111" => data_out <= rom_array(4231);
		when "0001000010001000" => data_out <= rom_array(4232);
		when "0001000010001001" => data_out <= rom_array(4233);
		when "0001000010001010" => data_out <= rom_array(4234);
		when "0001000010001011" => data_out <= rom_array(4235);
		when "0001000010001100" => data_out <= rom_array(4236);
		when "0001000010001101" => data_out <= rom_array(4237);
		when "0001000010001110" => data_out <= rom_array(4238);
		when "0001000010001111" => data_out <= rom_array(4239);
		when "0001000010010000" => data_out <= rom_array(4240);
		when "0001000010010001" => data_out <= rom_array(4241);
		when "0001000010010010" => data_out <= rom_array(4242);
		when "0001000010010011" => data_out <= rom_array(4243);
		when "0001000010010100" => data_out <= rom_array(4244);
		when "0001000010010101" => data_out <= rom_array(4245);
		when "0001000010010110" => data_out <= rom_array(4246);
		when "0001000010010111" => data_out <= rom_array(4247);
		when "0001000010011000" => data_out <= rom_array(4248);
		when "0001000010011001" => data_out <= rom_array(4249);
		when "0001000010011010" => data_out <= rom_array(4250);
		when "0001000010011011" => data_out <= rom_array(4251);
		when "0001000010011100" => data_out <= rom_array(4252);
		when "0001000010011101" => data_out <= rom_array(4253);
		when "0001000010011110" => data_out <= rom_array(4254);
		when "0001000010011111" => data_out <= rom_array(4255);
		when "0001000010100000" => data_out <= rom_array(4256);
		when "0001000010100001" => data_out <= rom_array(4257);
		when "0001000010100010" => data_out <= rom_array(4258);
		when "0001000010100011" => data_out <= rom_array(4259);
		when "0001000010100100" => data_out <= rom_array(4260);
		when "0001000010100101" => data_out <= rom_array(4261);
		when "0001000010100110" => data_out <= rom_array(4262);
		when "0001000010100111" => data_out <= rom_array(4263);
		when "0001000010101000" => data_out <= rom_array(4264);
		when "0001000010101001" => data_out <= rom_array(4265);
		when "0001000010101010" => data_out <= rom_array(4266);
		when "0001000010101011" => data_out <= rom_array(4267);
		when "0001000010101100" => data_out <= rom_array(4268);
		when "0001000010101101" => data_out <= rom_array(4269);
		when "0001000010101110" => data_out <= rom_array(4270);
		when "0001000010101111" => data_out <= rom_array(4271);
		when "0001000010110000" => data_out <= rom_array(4272);
		when "0001000010110001" => data_out <= rom_array(4273);
		when "0001000010110010" => data_out <= rom_array(4274);
		when "0001000010110011" => data_out <= rom_array(4275);
		when "0001000010110100" => data_out <= rom_array(4276);
		when "0001000010110101" => data_out <= rom_array(4277);
		when "0001000010110110" => data_out <= rom_array(4278);
		when "0001000010110111" => data_out <= rom_array(4279);
		when "0001000010111000" => data_out <= rom_array(4280);
		when "0001000010111001" => data_out <= rom_array(4281);
		when "0001000010111010" => data_out <= rom_array(4282);
		when "0001000010111011" => data_out <= rom_array(4283);
		when "0001000010111100" => data_out <= rom_array(4284);
		when "0001000010111101" => data_out <= rom_array(4285);
		when "0001000010111110" => data_out <= rom_array(4286);
		when "0001000010111111" => data_out <= rom_array(4287);
		when "0001000011000000" => data_out <= rom_array(4288);
		when "0001000011000001" => data_out <= rom_array(4289);
		when "0001000011000010" => data_out <= rom_array(4290);
		when "0001000011000011" => data_out <= rom_array(4291);
		when "0001000011000100" => data_out <= rom_array(4292);
		when "0001000011000101" => data_out <= rom_array(4293);
		when "0001000011000110" => data_out <= rom_array(4294);
		when "0001000011000111" => data_out <= rom_array(4295);
		when "0001000011001000" => data_out <= rom_array(4296);
		when "0001000011001001" => data_out <= rom_array(4297);
		when "0001000011001010" => data_out <= rom_array(4298);
		when "0001000011001011" => data_out <= rom_array(4299);
		when "0001000011001100" => data_out <= rom_array(4300);
		when "0001000011001101" => data_out <= rom_array(4301);
		when "0001000011001110" => data_out <= rom_array(4302);
		when "0001000011001111" => data_out <= rom_array(4303);
		when "0001000011010000" => data_out <= rom_array(4304);
		when "0001000011010001" => data_out <= rom_array(4305);
		when "0001000011010010" => data_out <= rom_array(4306);
		when "0001000011010011" => data_out <= rom_array(4307);
		when "0001000011010100" => data_out <= rom_array(4308);
		when "0001000011010101" => data_out <= rom_array(4309);
		when "0001000011010110" => data_out <= rom_array(4310);
		when "0001000011010111" => data_out <= rom_array(4311);
		when "0001000011011000" => data_out <= rom_array(4312);
		when "0001000011011001" => data_out <= rom_array(4313);
		when "0001000011011010" => data_out <= rom_array(4314);
		when "0001000011011011" => data_out <= rom_array(4315);
		when "0001000011011100" => data_out <= rom_array(4316);
		when "0001000011011101" => data_out <= rom_array(4317);
		when "0001000011011110" => data_out <= rom_array(4318);
		when "0001000011011111" => data_out <= rom_array(4319);
		when "0001000011100000" => data_out <= rom_array(4320);
		when "0001000011100001" => data_out <= rom_array(4321);
		when "0001000011100010" => data_out <= rom_array(4322);
		when "0001000011100011" => data_out <= rom_array(4323);
		when "0001000011100100" => data_out <= rom_array(4324);
		when "0001000011100101" => data_out <= rom_array(4325);
		when "0001000011100110" => data_out <= rom_array(4326);
		when "0001000011100111" => data_out <= rom_array(4327);
		when "0001000011101000" => data_out <= rom_array(4328);
		when "0001000011101001" => data_out <= rom_array(4329);
		when "0001000011101010" => data_out <= rom_array(4330);
		when "0001000011101011" => data_out <= rom_array(4331);
		when "0001000011101100" => data_out <= rom_array(4332);
		when "0001000011101101" => data_out <= rom_array(4333);
		when "0001000011101110" => data_out <= rom_array(4334);
		when "0001000011101111" => data_out <= rom_array(4335);
		when "0001000011110000" => data_out <= rom_array(4336);
		when "0001000011110001" => data_out <= rom_array(4337);
		when "0001000011110010" => data_out <= rom_array(4338);
		when "0001000011110011" => data_out <= rom_array(4339);
		when "0001000011110100" => data_out <= rom_array(4340);
		when "0001000011110101" => data_out <= rom_array(4341);
		when "0001000011110110" => data_out <= rom_array(4342);
		when "0001000011110111" => data_out <= rom_array(4343);
		when "0001000011111000" => data_out <= rom_array(4344);
		when "0001000011111001" => data_out <= rom_array(4345);
		when "0001000011111010" => data_out <= rom_array(4346);
		when "0001000011111011" => data_out <= rom_array(4347);
		when "0001000011111100" => data_out <= rom_array(4348);
		when "0001000011111101" => data_out <= rom_array(4349);
		when "0001000011111110" => data_out <= rom_array(4350);
		when "0001000011111111" => data_out <= rom_array(4351);
		when "0001000100000000" => data_out <= rom_array(4352);
		when "0001000100000001" => data_out <= rom_array(4353);
		when "0001000100000010" => data_out <= rom_array(4354);
		when "0001000100000011" => data_out <= rom_array(4355);
		when "0001000100000100" => data_out <= rom_array(4356);
		when "0001000100000101" => data_out <= rom_array(4357);
		when "0001000100000110" => data_out <= rom_array(4358);
		when "0001000100000111" => data_out <= rom_array(4359);
		when "0001000100001000" => data_out <= rom_array(4360);
		when "0001000100001001" => data_out <= rom_array(4361);
		when "0001000100001010" => data_out <= rom_array(4362);
		when "0001000100001011" => data_out <= rom_array(4363);
		when "0001000100001100" => data_out <= rom_array(4364);
		when "0001000100001101" => data_out <= rom_array(4365);
		when "0001000100001110" => data_out <= rom_array(4366);
		when "0001000100001111" => data_out <= rom_array(4367);
		when "0001000100010000" => data_out <= rom_array(4368);
		when "0001000100010001" => data_out <= rom_array(4369);
		when "0001000100010010" => data_out <= rom_array(4370);
		when "0001000100010011" => data_out <= rom_array(4371);
		when "0001000100010100" => data_out <= rom_array(4372);
		when "0001000100010101" => data_out <= rom_array(4373);
		when "0001000100010110" => data_out <= rom_array(4374);
		when "0001000100010111" => data_out <= rom_array(4375);
		when "0001000100011000" => data_out <= rom_array(4376);
		when "0001000100011001" => data_out <= rom_array(4377);
		when "0001000100011010" => data_out <= rom_array(4378);
		when "0001000100011011" => data_out <= rom_array(4379);
		when "0001000100011100" => data_out <= rom_array(4380);
		when "0001000100011101" => data_out <= rom_array(4381);
		when "0001000100011110" => data_out <= rom_array(4382);
		when "0001000100011111" => data_out <= rom_array(4383);
		when "0001000100100000" => data_out <= rom_array(4384);
		when "0001000100100001" => data_out <= rom_array(4385);
		when "0001000100100010" => data_out <= rom_array(4386);
		when "0001000100100011" => data_out <= rom_array(4387);
		when "0001000100100100" => data_out <= rom_array(4388);
		when "0001000100100101" => data_out <= rom_array(4389);
		when "0001000100100110" => data_out <= rom_array(4390);
		when "0001000100100111" => data_out <= rom_array(4391);
		when "0001000100101000" => data_out <= rom_array(4392);
		when "0001000100101001" => data_out <= rom_array(4393);
		when "0001000100101010" => data_out <= rom_array(4394);
		when "0001000100101011" => data_out <= rom_array(4395);
		when "0001000100101100" => data_out <= rom_array(4396);
		when "0001000100101101" => data_out <= rom_array(4397);
		when "0001000100101110" => data_out <= rom_array(4398);
		when "0001000100101111" => data_out <= rom_array(4399);
		when "0001000100110000" => data_out <= rom_array(4400);
		when "0001000100110001" => data_out <= rom_array(4401);
		when "0001000100110010" => data_out <= rom_array(4402);
		when "0001000100110011" => data_out <= rom_array(4403);
		when "0001000100110100" => data_out <= rom_array(4404);
		when "0001000100110101" => data_out <= rom_array(4405);
		when "0001000100110110" => data_out <= rom_array(4406);
		when "0001000100110111" => data_out <= rom_array(4407);
		when "0001000100111000" => data_out <= rom_array(4408);
		when "0001000100111001" => data_out <= rom_array(4409);
		when "0001000100111010" => data_out <= rom_array(4410);
		when "0001000100111011" => data_out <= rom_array(4411);
		when "0001000100111100" => data_out <= rom_array(4412);
		when "0001000100111101" => data_out <= rom_array(4413);
		when "0001000100111110" => data_out <= rom_array(4414);
		when "0001000100111111" => data_out <= rom_array(4415);
		when "0001000101000000" => data_out <= rom_array(4416);
		when "0001000101000001" => data_out <= rom_array(4417);
		when "0001000101000010" => data_out <= rom_array(4418);
		when "0001000101000011" => data_out <= rom_array(4419);
		when "0001000101000100" => data_out <= rom_array(4420);
		when "0001000101000101" => data_out <= rom_array(4421);
		when "0001000101000110" => data_out <= rom_array(4422);
		when "0001000101000111" => data_out <= rom_array(4423);
		when "0001000101001000" => data_out <= rom_array(4424);
		when "0001000101001001" => data_out <= rom_array(4425);
		when "0001000101001010" => data_out <= rom_array(4426);
		when "0001000101001011" => data_out <= rom_array(4427);
		when "0001000101001100" => data_out <= rom_array(4428);
		when "0001000101001101" => data_out <= rom_array(4429);
		when "0001000101001110" => data_out <= rom_array(4430);
		when "0001000101001111" => data_out <= rom_array(4431);
		when "0001000101010000" => data_out <= rom_array(4432);
		when "0001000101010001" => data_out <= rom_array(4433);
		when "0001000101010010" => data_out <= rom_array(4434);
		when "0001000101010011" => data_out <= rom_array(4435);
		when "0001000101010100" => data_out <= rom_array(4436);
		when "0001000101010101" => data_out <= rom_array(4437);
		when "0001000101010110" => data_out <= rom_array(4438);
		when "0001000101010111" => data_out <= rom_array(4439);
		when "0001000101011000" => data_out <= rom_array(4440);
		when "0001000101011001" => data_out <= rom_array(4441);
		when "0001000101011010" => data_out <= rom_array(4442);
		when "0001000101011011" => data_out <= rom_array(4443);
		when "0001000101011100" => data_out <= rom_array(4444);
		when "0001000101011101" => data_out <= rom_array(4445);
		when "0001000101011110" => data_out <= rom_array(4446);
		when "0001000101011111" => data_out <= rom_array(4447);
		when "0001000101100000" => data_out <= rom_array(4448);
		when "0001000101100001" => data_out <= rom_array(4449);
		when "0001000101100010" => data_out <= rom_array(4450);
		when "0001000101100011" => data_out <= rom_array(4451);
		when "0001000101100100" => data_out <= rom_array(4452);
		when "0001000101100101" => data_out <= rom_array(4453);
		when "0001000101100110" => data_out <= rom_array(4454);
		when "0001000101100111" => data_out <= rom_array(4455);
		when "0001000101101000" => data_out <= rom_array(4456);
		when "0001000101101001" => data_out <= rom_array(4457);
		when "0001000101101010" => data_out <= rom_array(4458);
		when "0001000101101011" => data_out <= rom_array(4459);
		when "0001000101101100" => data_out <= rom_array(4460);
		when "0001000101101101" => data_out <= rom_array(4461);
		when "0001000101101110" => data_out <= rom_array(4462);
		when "0001000101101111" => data_out <= rom_array(4463);
		when "0001000101110000" => data_out <= rom_array(4464);
		when "0001000101110001" => data_out <= rom_array(4465);
		when "0001000101110010" => data_out <= rom_array(4466);
		when "0001000101110011" => data_out <= rom_array(4467);
		when "0001000101110100" => data_out <= rom_array(4468);
		when "0001000101110101" => data_out <= rom_array(4469);
		when "0001000101110110" => data_out <= rom_array(4470);
		when "0001000101110111" => data_out <= rom_array(4471);
		when "0001000101111000" => data_out <= rom_array(4472);
		when "0001000101111001" => data_out <= rom_array(4473);
		when "0001000101111010" => data_out <= rom_array(4474);
		when "0001000101111011" => data_out <= rom_array(4475);
		when "0001000101111100" => data_out <= rom_array(4476);
		when "0001000101111101" => data_out <= rom_array(4477);
		when "0001000101111110" => data_out <= rom_array(4478);
		when "0001000101111111" => data_out <= rom_array(4479);
		when "0001000110000000" => data_out <= rom_array(4480);
		when "0001000110000001" => data_out <= rom_array(4481);
		when "0001000110000010" => data_out <= rom_array(4482);
		when "0001000110000011" => data_out <= rom_array(4483);
		when "0001000110000100" => data_out <= rom_array(4484);
		when "0001000110000101" => data_out <= rom_array(4485);
		when "0001000110000110" => data_out <= rom_array(4486);
		when "0001000110000111" => data_out <= rom_array(4487);
		when "0001000110001000" => data_out <= rom_array(4488);
		when "0001000110001001" => data_out <= rom_array(4489);
		when "0001000110001010" => data_out <= rom_array(4490);
		when "0001000110001011" => data_out <= rom_array(4491);
		when "0001000110001100" => data_out <= rom_array(4492);
		when "0001000110001101" => data_out <= rom_array(4493);
		when "0001000110001110" => data_out <= rom_array(4494);
		when "0001000110001111" => data_out <= rom_array(4495);
		when "0001000110010000" => data_out <= rom_array(4496);
		when "0001000110010001" => data_out <= rom_array(4497);
		when "0001000110010010" => data_out <= rom_array(4498);
		when "0001000110010011" => data_out <= rom_array(4499);
		when "0001000110010100" => data_out <= rom_array(4500);
		when "0001000110010101" => data_out <= rom_array(4501);
		when "0001000110010110" => data_out <= rom_array(4502);
		when "0001000110010111" => data_out <= rom_array(4503);
		when "0001000110011000" => data_out <= rom_array(4504);
		when "0001000110011001" => data_out <= rom_array(4505);
		when "0001000110011010" => data_out <= rom_array(4506);
		when "0001000110011011" => data_out <= rom_array(4507);
		when "0001000110011100" => data_out <= rom_array(4508);
		when "0001000110011101" => data_out <= rom_array(4509);
		when "0001000110011110" => data_out <= rom_array(4510);
		when "0001000110011111" => data_out <= rom_array(4511);
		when "0001000110100000" => data_out <= rom_array(4512);
		when "0001000110100001" => data_out <= rom_array(4513);
		when "0001000110100010" => data_out <= rom_array(4514);
		when "0001000110100011" => data_out <= rom_array(4515);
		when "0001000110100100" => data_out <= rom_array(4516);
		when "0001000110100101" => data_out <= rom_array(4517);
		when "0001000110100110" => data_out <= rom_array(4518);
		when "0001000110100111" => data_out <= rom_array(4519);
		when "0001000110101000" => data_out <= rom_array(4520);
		when "0001000110101001" => data_out <= rom_array(4521);
		when "0001000110101010" => data_out <= rom_array(4522);
		when "0001000110101011" => data_out <= rom_array(4523);
		when "0001000110101100" => data_out <= rom_array(4524);
		when "0001000110101101" => data_out <= rom_array(4525);
		when "0001000110101110" => data_out <= rom_array(4526);
		when "0001000110101111" => data_out <= rom_array(4527);
		when "0001000110110000" => data_out <= rom_array(4528);
		when "0001000110110001" => data_out <= rom_array(4529);
		when "0001000110110010" => data_out <= rom_array(4530);
		when "0001000110110011" => data_out <= rom_array(4531);
		when "0001000110110100" => data_out <= rom_array(4532);
		when "0001000110110101" => data_out <= rom_array(4533);
		when "0001000110110110" => data_out <= rom_array(4534);
		when "0001000110110111" => data_out <= rom_array(4535);
		when "0001000110111000" => data_out <= rom_array(4536);
		when "0001000110111001" => data_out <= rom_array(4537);
		when "0001000110111010" => data_out <= rom_array(4538);
		when "0001000110111011" => data_out <= rom_array(4539);
		when "0001000110111100" => data_out <= rom_array(4540);
		when "0001000110111101" => data_out <= rom_array(4541);
		when "0001000110111110" => data_out <= rom_array(4542);
		when "0001000110111111" => data_out <= rom_array(4543);
		when "0001000111000000" => data_out <= rom_array(4544);
		when "0001000111000001" => data_out <= rom_array(4545);
		when "0001000111000010" => data_out <= rom_array(4546);
		when "0001000111000011" => data_out <= rom_array(4547);
		when "0001000111000100" => data_out <= rom_array(4548);
		when "0001000111000101" => data_out <= rom_array(4549);
		when "0001000111000110" => data_out <= rom_array(4550);
		when "0001000111000111" => data_out <= rom_array(4551);
		when "0001000111001000" => data_out <= rom_array(4552);
		when "0001000111001001" => data_out <= rom_array(4553);
		when "0001000111001010" => data_out <= rom_array(4554);
		when "0001000111001011" => data_out <= rom_array(4555);
		when "0001000111001100" => data_out <= rom_array(4556);
		when "0001000111001101" => data_out <= rom_array(4557);
		when "0001000111001110" => data_out <= rom_array(4558);
		when "0001000111001111" => data_out <= rom_array(4559);
		when "0001000111010000" => data_out <= rom_array(4560);
		when "0001000111010001" => data_out <= rom_array(4561);
		when "0001000111010010" => data_out <= rom_array(4562);
		when "0001000111010011" => data_out <= rom_array(4563);
		when "0001000111010100" => data_out <= rom_array(4564);
		when "0001000111010101" => data_out <= rom_array(4565);
		when "0001000111010110" => data_out <= rom_array(4566);
		when "0001000111010111" => data_out <= rom_array(4567);
		when "0001000111011000" => data_out <= rom_array(4568);
		when "0001000111011001" => data_out <= rom_array(4569);
		when "0001000111011010" => data_out <= rom_array(4570);
		when "0001000111011011" => data_out <= rom_array(4571);
		when "0001000111011100" => data_out <= rom_array(4572);
		when "0001000111011101" => data_out <= rom_array(4573);
		when "0001000111011110" => data_out <= rom_array(4574);
		when "0001000111011111" => data_out <= rom_array(4575);
		when "0001000111100000" => data_out <= rom_array(4576);
		when "0001000111100001" => data_out <= rom_array(4577);
		when "0001000111100010" => data_out <= rom_array(4578);
		when "0001000111100011" => data_out <= rom_array(4579);
		when "0001000111100100" => data_out <= rom_array(4580);
		when "0001000111100101" => data_out <= rom_array(4581);
		when "0001000111100110" => data_out <= rom_array(4582);
		when "0001000111100111" => data_out <= rom_array(4583);
		when "0001000111101000" => data_out <= rom_array(4584);
		when "0001000111101001" => data_out <= rom_array(4585);
		when "0001000111101010" => data_out <= rom_array(4586);
		when "0001000111101011" => data_out <= rom_array(4587);
		when "0001000111101100" => data_out <= rom_array(4588);
		when "0001000111101101" => data_out <= rom_array(4589);
		when "0001000111101110" => data_out <= rom_array(4590);
		when "0001000111101111" => data_out <= rom_array(4591);
		when "0001000111110000" => data_out <= rom_array(4592);
		when "0001000111110001" => data_out <= rom_array(4593);
		when "0001000111110010" => data_out <= rom_array(4594);
		when "0001000111110011" => data_out <= rom_array(4595);
		when "0001000111110100" => data_out <= rom_array(4596);
		when "0001000111110101" => data_out <= rom_array(4597);
		when "0001000111110110" => data_out <= rom_array(4598);
		when "0001000111110111" => data_out <= rom_array(4599);
		when "0001000111111000" => data_out <= rom_array(4600);
		when "0001000111111001" => data_out <= rom_array(4601);
		when "0001000111111010" => data_out <= rom_array(4602);
		when "0001000111111011" => data_out <= rom_array(4603);
		when "0001000111111100" => data_out <= rom_array(4604);
		when "0001000111111101" => data_out <= rom_array(4605);
		when "0001000111111110" => data_out <= rom_array(4606);
		when "0001000111111111" => data_out <= rom_array(4607);
		when "0001001000000000" => data_out <= rom_array(4608);
		when "0001001000000001" => data_out <= rom_array(4609);
		when "0001001000000010" => data_out <= rom_array(4610);
		when "0001001000000011" => data_out <= rom_array(4611);
		when "0001001000000100" => data_out <= rom_array(4612);
		when "0001001000000101" => data_out <= rom_array(4613);
		when "0001001000000110" => data_out <= rom_array(4614);
		when "0001001000000111" => data_out <= rom_array(4615);
		when "0001001000001000" => data_out <= rom_array(4616);
		when "0001001000001001" => data_out <= rom_array(4617);
		when "0001001000001010" => data_out <= rom_array(4618);
		when "0001001000001011" => data_out <= rom_array(4619);
		when "0001001000001100" => data_out <= rom_array(4620);
		when "0001001000001101" => data_out <= rom_array(4621);
		when "0001001000001110" => data_out <= rom_array(4622);
		when "0001001000001111" => data_out <= rom_array(4623);
		when "0001001000010000" => data_out <= rom_array(4624);
		when "0001001000010001" => data_out <= rom_array(4625);
		when "0001001000010010" => data_out <= rom_array(4626);
		when "0001001000010011" => data_out <= rom_array(4627);
		when "0001001000010100" => data_out <= rom_array(4628);
		when "0001001000010101" => data_out <= rom_array(4629);
		when "0001001000010110" => data_out <= rom_array(4630);
		when "0001001000010111" => data_out <= rom_array(4631);
		when "0001001000011000" => data_out <= rom_array(4632);
		when "0001001000011001" => data_out <= rom_array(4633);
		when "0001001000011010" => data_out <= rom_array(4634);
		when "0001001000011011" => data_out <= rom_array(4635);
		when "0001001000011100" => data_out <= rom_array(4636);
		when "0001001000011101" => data_out <= rom_array(4637);
		when "0001001000011110" => data_out <= rom_array(4638);
		when "0001001000011111" => data_out <= rom_array(4639);
		when "0001001000100000" => data_out <= rom_array(4640);
		when "0001001000100001" => data_out <= rom_array(4641);
		when "0001001000100010" => data_out <= rom_array(4642);
		when "0001001000100011" => data_out <= rom_array(4643);
		when "0001001000100100" => data_out <= rom_array(4644);
		when "0001001000100101" => data_out <= rom_array(4645);
		when "0001001000100110" => data_out <= rom_array(4646);
		when "0001001000100111" => data_out <= rom_array(4647);
		when "0001001000101000" => data_out <= rom_array(4648);
		when "0001001000101001" => data_out <= rom_array(4649);
		when "0001001000101010" => data_out <= rom_array(4650);
		when "0001001000101011" => data_out <= rom_array(4651);
		when "0001001000101100" => data_out <= rom_array(4652);
		when "0001001000101101" => data_out <= rom_array(4653);
		when "0001001000101110" => data_out <= rom_array(4654);
		when "0001001000101111" => data_out <= rom_array(4655);
		when "0001001000110000" => data_out <= rom_array(4656);
		when "0001001000110001" => data_out <= rom_array(4657);
		when "0001001000110010" => data_out <= rom_array(4658);
		when "0001001000110011" => data_out <= rom_array(4659);
		when "0001001000110100" => data_out <= rom_array(4660);
		when "0001001000110101" => data_out <= rom_array(4661);
		when "0001001000110110" => data_out <= rom_array(4662);
		when "0001001000110111" => data_out <= rom_array(4663);
		when "0001001000111000" => data_out <= rom_array(4664);
		when "0001001000111001" => data_out <= rom_array(4665);
		when "0001001000111010" => data_out <= rom_array(4666);
		when "0001001000111011" => data_out <= rom_array(4667);
		when "0001001000111100" => data_out <= rom_array(4668);
		when "0001001000111101" => data_out <= rom_array(4669);
		when "0001001000111110" => data_out <= rom_array(4670);
		when "0001001000111111" => data_out <= rom_array(4671);
		when "0001001001000000" => data_out <= rom_array(4672);
		when "0001001001000001" => data_out <= rom_array(4673);
		when "0001001001000010" => data_out <= rom_array(4674);
		when "0001001001000011" => data_out <= rom_array(4675);
		when "0001001001000100" => data_out <= rom_array(4676);
		when "0001001001000101" => data_out <= rom_array(4677);
		when "0001001001000110" => data_out <= rom_array(4678);
		when "0001001001000111" => data_out <= rom_array(4679);
		when "0001001001001000" => data_out <= rom_array(4680);
		when "0001001001001001" => data_out <= rom_array(4681);
		when "0001001001001010" => data_out <= rom_array(4682);
		when "0001001001001011" => data_out <= rom_array(4683);
		when "0001001001001100" => data_out <= rom_array(4684);
		when "0001001001001101" => data_out <= rom_array(4685);
		when "0001001001001110" => data_out <= rom_array(4686);
		when "0001001001001111" => data_out <= rom_array(4687);
		when "0001001001010000" => data_out <= rom_array(4688);
		when "0001001001010001" => data_out <= rom_array(4689);
		when "0001001001010010" => data_out <= rom_array(4690);
		when "0001001001010011" => data_out <= rom_array(4691);
		when "0001001001010100" => data_out <= rom_array(4692);
		when "0001001001010101" => data_out <= rom_array(4693);
		when "0001001001010110" => data_out <= rom_array(4694);
		when "0001001001010111" => data_out <= rom_array(4695);
		when "0001001001011000" => data_out <= rom_array(4696);
		when "0001001001011001" => data_out <= rom_array(4697);
		when "0001001001011010" => data_out <= rom_array(4698);
		when "0001001001011011" => data_out <= rom_array(4699);
		when "0001001001011100" => data_out <= rom_array(4700);
		when "0001001001011101" => data_out <= rom_array(4701);
		when "0001001001011110" => data_out <= rom_array(4702);
		when "0001001001011111" => data_out <= rom_array(4703);
		when "0001001001100000" => data_out <= rom_array(4704);
		when "0001001001100001" => data_out <= rom_array(4705);
		when "0001001001100010" => data_out <= rom_array(4706);
		when "0001001001100011" => data_out <= rom_array(4707);
		when "0001001001100100" => data_out <= rom_array(4708);
		when "0001001001100101" => data_out <= rom_array(4709);
		when "0001001001100110" => data_out <= rom_array(4710);
		when "0001001001100111" => data_out <= rom_array(4711);
		when "0001001001101000" => data_out <= rom_array(4712);
		when "0001001001101001" => data_out <= rom_array(4713);
		when "0001001001101010" => data_out <= rom_array(4714);
		when "0001001001101011" => data_out <= rom_array(4715);
		when "0001001001101100" => data_out <= rom_array(4716);
		when "0001001001101101" => data_out <= rom_array(4717);
		when "0001001001101110" => data_out <= rom_array(4718);
		when "0001001001101111" => data_out <= rom_array(4719);
		when "0001001001110000" => data_out <= rom_array(4720);
		when "0001001001110001" => data_out <= rom_array(4721);
		when "0001001001110010" => data_out <= rom_array(4722);
		when "0001001001110011" => data_out <= rom_array(4723);
		when "0001001001110100" => data_out <= rom_array(4724);
		when "0001001001110101" => data_out <= rom_array(4725);
		when "0001001001110110" => data_out <= rom_array(4726);
		when "0001001001110111" => data_out <= rom_array(4727);
		when "0001001001111000" => data_out <= rom_array(4728);
		when "0001001001111001" => data_out <= rom_array(4729);
		when "0001001001111010" => data_out <= rom_array(4730);
		when "0001001001111011" => data_out <= rom_array(4731);
		when "0001001001111100" => data_out <= rom_array(4732);
		when "0001001001111101" => data_out <= rom_array(4733);
		when "0001001001111110" => data_out <= rom_array(4734);
		when "0001001001111111" => data_out <= rom_array(4735);
		when "0001001010000000" => data_out <= rom_array(4736);
		when "0001001010000001" => data_out <= rom_array(4737);
		when "0001001010000010" => data_out <= rom_array(4738);
		when "0001001010000011" => data_out <= rom_array(4739);
		when "0001001010000100" => data_out <= rom_array(4740);
		when "0001001010000101" => data_out <= rom_array(4741);
		when "0001001010000110" => data_out <= rom_array(4742);
		when "0001001010000111" => data_out <= rom_array(4743);
		when "0001001010001000" => data_out <= rom_array(4744);
		when "0001001010001001" => data_out <= rom_array(4745);
		when "0001001010001010" => data_out <= rom_array(4746);
		when "0001001010001011" => data_out <= rom_array(4747);
		when "0001001010001100" => data_out <= rom_array(4748);
		when "0001001010001101" => data_out <= rom_array(4749);
		when "0001001010001110" => data_out <= rom_array(4750);
		when "0001001010001111" => data_out <= rom_array(4751);
		when "0001001010010000" => data_out <= rom_array(4752);
		when "0001001010010001" => data_out <= rom_array(4753);
		when "0001001010010010" => data_out <= rom_array(4754);
		when "0001001010010011" => data_out <= rom_array(4755);
		when "0001001010010100" => data_out <= rom_array(4756);
		when "0001001010010101" => data_out <= rom_array(4757);
		when "0001001010010110" => data_out <= rom_array(4758);
		when "0001001010010111" => data_out <= rom_array(4759);
		when "0001001010011000" => data_out <= rom_array(4760);
		when "0001001010011001" => data_out <= rom_array(4761);
		when "0001001010011010" => data_out <= rom_array(4762);
		when "0001001010011011" => data_out <= rom_array(4763);
		when "0001001010011100" => data_out <= rom_array(4764);
		when "0001001010011101" => data_out <= rom_array(4765);
		when "0001001010011110" => data_out <= rom_array(4766);
		when "0001001010011111" => data_out <= rom_array(4767);
		when "0001001010100000" => data_out <= rom_array(4768);
		when "0001001010100001" => data_out <= rom_array(4769);
		when "0001001010100010" => data_out <= rom_array(4770);
		when "0001001010100011" => data_out <= rom_array(4771);
		when "0001001010100100" => data_out <= rom_array(4772);
		when "0001001010100101" => data_out <= rom_array(4773);
		when "0001001010100110" => data_out <= rom_array(4774);
		when "0001001010100111" => data_out <= rom_array(4775);
		when "0001001010101000" => data_out <= rom_array(4776);
		when "0001001010101001" => data_out <= rom_array(4777);
		when "0001001010101010" => data_out <= rom_array(4778);
		when "0001001010101011" => data_out <= rom_array(4779);
		when "0001001010101100" => data_out <= rom_array(4780);
		when "0001001010101101" => data_out <= rom_array(4781);
		when "0001001010101110" => data_out <= rom_array(4782);
		when "0001001010101111" => data_out <= rom_array(4783);
		when "0001001010110000" => data_out <= rom_array(4784);
		when "0001001010110001" => data_out <= rom_array(4785);
		when "0001001010110010" => data_out <= rom_array(4786);
		when "0001001010110011" => data_out <= rom_array(4787);
		when "0001001010110100" => data_out <= rom_array(4788);
		when "0001001010110101" => data_out <= rom_array(4789);
		when "0001001010110110" => data_out <= rom_array(4790);
		when "0001001010110111" => data_out <= rom_array(4791);
		when "0001001010111000" => data_out <= rom_array(4792);
		when "0001001010111001" => data_out <= rom_array(4793);
		when "0001001010111010" => data_out <= rom_array(4794);
		when "0001001010111011" => data_out <= rom_array(4795);
		when "0001001010111100" => data_out <= rom_array(4796);
		when "0001001010111101" => data_out <= rom_array(4797);
		when "0001001010111110" => data_out <= rom_array(4798);
		when "0001001010111111" => data_out <= rom_array(4799);
		when "0001001011000000" => data_out <= rom_array(4800);
		when "0001001011000001" => data_out <= rom_array(4801);
		when "0001001011000010" => data_out <= rom_array(4802);
		when "0001001011000011" => data_out <= rom_array(4803);
		when "0001001011000100" => data_out <= rom_array(4804);
		when "0001001011000101" => data_out <= rom_array(4805);
		when "0001001011000110" => data_out <= rom_array(4806);
		when "0001001011000111" => data_out <= rom_array(4807);
		when "0001001011001000" => data_out <= rom_array(4808);
		when "0001001011001001" => data_out <= rom_array(4809);
		when "0001001011001010" => data_out <= rom_array(4810);
		when "0001001011001011" => data_out <= rom_array(4811);
		when "0001001011001100" => data_out <= rom_array(4812);
		when "0001001011001101" => data_out <= rom_array(4813);
		when "0001001011001110" => data_out <= rom_array(4814);
		when "0001001011001111" => data_out <= rom_array(4815);
		when "0001001011010000" => data_out <= rom_array(4816);
		when "0001001011010001" => data_out <= rom_array(4817);
		when "0001001011010010" => data_out <= rom_array(4818);
		when "0001001011010011" => data_out <= rom_array(4819);
		when "0001001011010100" => data_out <= rom_array(4820);
		when "0001001011010101" => data_out <= rom_array(4821);
		when "0001001011010110" => data_out <= rom_array(4822);
		when "0001001011010111" => data_out <= rom_array(4823);
		when "0001001011011000" => data_out <= rom_array(4824);
		when "0001001011011001" => data_out <= rom_array(4825);
		when "0001001011011010" => data_out <= rom_array(4826);
		when "0001001011011011" => data_out <= rom_array(4827);
		when "0001001011011100" => data_out <= rom_array(4828);
		when "0001001011011101" => data_out <= rom_array(4829);
		when "0001001011011110" => data_out <= rom_array(4830);
		when "0001001011011111" => data_out <= rom_array(4831);
		when "0001001011100000" => data_out <= rom_array(4832);
		when "0001001011100001" => data_out <= rom_array(4833);
		when "0001001011100010" => data_out <= rom_array(4834);
		when "0001001011100011" => data_out <= rom_array(4835);
		when "0001001011100100" => data_out <= rom_array(4836);
		when "0001001011100101" => data_out <= rom_array(4837);
		when "0001001011100110" => data_out <= rom_array(4838);
		when "0001001011100111" => data_out <= rom_array(4839);
		when "0001001011101000" => data_out <= rom_array(4840);
		when "0001001011101001" => data_out <= rom_array(4841);
		when "0001001011101010" => data_out <= rom_array(4842);
		when "0001001011101011" => data_out <= rom_array(4843);
		when "0001001011101100" => data_out <= rom_array(4844);
		when "0001001011101101" => data_out <= rom_array(4845);
		when "0001001011101110" => data_out <= rom_array(4846);
		when "0001001011101111" => data_out <= rom_array(4847);
		when "0001001011110000" => data_out <= rom_array(4848);
		when "0001001011110001" => data_out <= rom_array(4849);
		when "0001001011110010" => data_out <= rom_array(4850);
		when "0001001011110011" => data_out <= rom_array(4851);
		when "0001001011110100" => data_out <= rom_array(4852);
		when "0001001011110101" => data_out <= rom_array(4853);
		when "0001001011110110" => data_out <= rom_array(4854);
		when "0001001011110111" => data_out <= rom_array(4855);
		when "0001001011111000" => data_out <= rom_array(4856);
		when "0001001011111001" => data_out <= rom_array(4857);
		when "0001001011111010" => data_out <= rom_array(4858);
		when "0001001011111011" => data_out <= rom_array(4859);
		when "0001001011111100" => data_out <= rom_array(4860);
		when "0001001011111101" => data_out <= rom_array(4861);
		when "0001001011111110" => data_out <= rom_array(4862);
		when "0001001011111111" => data_out <= rom_array(4863);
		when "0001001100000000" => data_out <= rom_array(4864);
		when "0001001100000001" => data_out <= rom_array(4865);
		when "0001001100000010" => data_out <= rom_array(4866);
		when "0001001100000011" => data_out <= rom_array(4867);
		when "0001001100000100" => data_out <= rom_array(4868);
		when "0001001100000101" => data_out <= rom_array(4869);
		when "0001001100000110" => data_out <= rom_array(4870);
		when "0001001100000111" => data_out <= rom_array(4871);
		when "0001001100001000" => data_out <= rom_array(4872);
		when "0001001100001001" => data_out <= rom_array(4873);
		when "0001001100001010" => data_out <= rom_array(4874);
		when "0001001100001011" => data_out <= rom_array(4875);
		when "0001001100001100" => data_out <= rom_array(4876);
		when "0001001100001101" => data_out <= rom_array(4877);
		when "0001001100001110" => data_out <= rom_array(4878);
		when "0001001100001111" => data_out <= rom_array(4879);
		when "0001001100010000" => data_out <= rom_array(4880);
		when "0001001100010001" => data_out <= rom_array(4881);
		when "0001001100010010" => data_out <= rom_array(4882);
		when "0001001100010011" => data_out <= rom_array(4883);
		when "0001001100010100" => data_out <= rom_array(4884);
		when "0001001100010101" => data_out <= rom_array(4885);
		when "0001001100010110" => data_out <= rom_array(4886);
		when "0001001100010111" => data_out <= rom_array(4887);
		when "0001001100011000" => data_out <= rom_array(4888);
		when "0001001100011001" => data_out <= rom_array(4889);
		when "0001001100011010" => data_out <= rom_array(4890);
		when "0001001100011011" => data_out <= rom_array(4891);
		when "0001001100011100" => data_out <= rom_array(4892);
		when "0001001100011101" => data_out <= rom_array(4893);
		when "0001001100011110" => data_out <= rom_array(4894);
		when "0001001100011111" => data_out <= rom_array(4895);
		when "0001001100100000" => data_out <= rom_array(4896);
		when "0001001100100001" => data_out <= rom_array(4897);
		when "0001001100100010" => data_out <= rom_array(4898);
		when "0001001100100011" => data_out <= rom_array(4899);
		when "0001001100100100" => data_out <= rom_array(4900);
		when "0001001100100101" => data_out <= rom_array(4901);
		when "0001001100100110" => data_out <= rom_array(4902);
		when "0001001100100111" => data_out <= rom_array(4903);
		when "0001001100101000" => data_out <= rom_array(4904);
		when "0001001100101001" => data_out <= rom_array(4905);
		when "0001001100101010" => data_out <= rom_array(4906);
		when "0001001100101011" => data_out <= rom_array(4907);
		when "0001001100101100" => data_out <= rom_array(4908);
		when "0001001100101101" => data_out <= rom_array(4909);
		when "0001001100101110" => data_out <= rom_array(4910);
		when "0001001100101111" => data_out <= rom_array(4911);
		when "0001001100110000" => data_out <= rom_array(4912);
		when "0001001100110001" => data_out <= rom_array(4913);
		when "0001001100110010" => data_out <= rom_array(4914);
		when "0001001100110011" => data_out <= rom_array(4915);
		when "0001001100110100" => data_out <= rom_array(4916);
		when "0001001100110101" => data_out <= rom_array(4917);
		when "0001001100110110" => data_out <= rom_array(4918);
		when "0001001100110111" => data_out <= rom_array(4919);
		when "0001001100111000" => data_out <= rom_array(4920);
		when "0001001100111001" => data_out <= rom_array(4921);
		when "0001001100111010" => data_out <= rom_array(4922);
		when "0001001100111011" => data_out <= rom_array(4923);
		when "0001001100111100" => data_out <= rom_array(4924);
		when "0001001100111101" => data_out <= rom_array(4925);
		when "0001001100111110" => data_out <= rom_array(4926);
		when "0001001100111111" => data_out <= rom_array(4927);
		when "0001001101000000" => data_out <= rom_array(4928);
		when "0001001101000001" => data_out <= rom_array(4929);
		when "0001001101000010" => data_out <= rom_array(4930);
		when "0001001101000011" => data_out <= rom_array(4931);
		when "0001001101000100" => data_out <= rom_array(4932);
		when "0001001101000101" => data_out <= rom_array(4933);
		when "0001001101000110" => data_out <= rom_array(4934);
		when "0001001101000111" => data_out <= rom_array(4935);
		when "0001001101001000" => data_out <= rom_array(4936);
		when "0001001101001001" => data_out <= rom_array(4937);
		when "0001001101001010" => data_out <= rom_array(4938);
		when "0001001101001011" => data_out <= rom_array(4939);
		when "0001001101001100" => data_out <= rom_array(4940);
		when "0001001101001101" => data_out <= rom_array(4941);
		when "0001001101001110" => data_out <= rom_array(4942);
		when "0001001101001111" => data_out <= rom_array(4943);
		when "0001001101010000" => data_out <= rom_array(4944);
		when "0001001101010001" => data_out <= rom_array(4945);
		when "0001001101010010" => data_out <= rom_array(4946);
		when "0001001101010011" => data_out <= rom_array(4947);
		when "0001001101010100" => data_out <= rom_array(4948);
		when "0001001101010101" => data_out <= rom_array(4949);
		when "0001001101010110" => data_out <= rom_array(4950);
		when "0001001101010111" => data_out <= rom_array(4951);
		when "0001001101011000" => data_out <= rom_array(4952);
		when "0001001101011001" => data_out <= rom_array(4953);
		when "0001001101011010" => data_out <= rom_array(4954);
		when "0001001101011011" => data_out <= rom_array(4955);
		when "0001001101011100" => data_out <= rom_array(4956);
		when "0001001101011101" => data_out <= rom_array(4957);
		when "0001001101011110" => data_out <= rom_array(4958);
		when "0001001101011111" => data_out <= rom_array(4959);
		when "0001001101100000" => data_out <= rom_array(4960);
		when "0001001101100001" => data_out <= rom_array(4961);
		when "0001001101100010" => data_out <= rom_array(4962);
		when "0001001101100011" => data_out <= rom_array(4963);
		when "0001001101100100" => data_out <= rom_array(4964);
		when "0001001101100101" => data_out <= rom_array(4965);
		when "0001001101100110" => data_out <= rom_array(4966);
		when "0001001101100111" => data_out <= rom_array(4967);
		when "0001001101101000" => data_out <= rom_array(4968);
		when "0001001101101001" => data_out <= rom_array(4969);
		when "0001001101101010" => data_out <= rom_array(4970);
		when "0001001101101011" => data_out <= rom_array(4971);
		when "0001001101101100" => data_out <= rom_array(4972);
		when "0001001101101101" => data_out <= rom_array(4973);
		when "0001001101101110" => data_out <= rom_array(4974);
		when "0001001101101111" => data_out <= rom_array(4975);
		when "0001001101110000" => data_out <= rom_array(4976);
		when "0001001101110001" => data_out <= rom_array(4977);
		when "0001001101110010" => data_out <= rom_array(4978);
		when "0001001101110011" => data_out <= rom_array(4979);
		when "0001001101110100" => data_out <= rom_array(4980);
		when "0001001101110101" => data_out <= rom_array(4981);
		when "0001001101110110" => data_out <= rom_array(4982);
		when "0001001101110111" => data_out <= rom_array(4983);
		when "0001001101111000" => data_out <= rom_array(4984);
		when "0001001101111001" => data_out <= rom_array(4985);
		when "0001001101111010" => data_out <= rom_array(4986);
		when "0001001101111011" => data_out <= rom_array(4987);
		when "0001001101111100" => data_out <= rom_array(4988);
		when "0001001101111101" => data_out <= rom_array(4989);
		when "0001001101111110" => data_out <= rom_array(4990);
		when "0001001101111111" => data_out <= rom_array(4991);
		when "0001001110000000" => data_out <= rom_array(4992);
		when "0001001110000001" => data_out <= rom_array(4993);
		when "0001001110000010" => data_out <= rom_array(4994);
		when "0001001110000011" => data_out <= rom_array(4995);
		when "0001001110000100" => data_out <= rom_array(4996);
		when "0001001110000101" => data_out <= rom_array(4997);
		when "0001001110000110" => data_out <= rom_array(4998);
		when "0001001110000111" => data_out <= rom_array(4999);
		when "0001001110001000" => data_out <= rom_array(5000);
		when "0001001110001001" => data_out <= rom_array(5001);
		when "0001001110001010" => data_out <= rom_array(5002);
		when "0001001110001011" => data_out <= rom_array(5003);
		when "0001001110001100" => data_out <= rom_array(5004);
		when "0001001110001101" => data_out <= rom_array(5005);
		when "0001001110001110" => data_out <= rom_array(5006);
		when "0001001110001111" => data_out <= rom_array(5007);
		when "0001001110010000" => data_out <= rom_array(5008);
		when "0001001110010001" => data_out <= rom_array(5009);
		when "0001001110010010" => data_out <= rom_array(5010);
		when "0001001110010011" => data_out <= rom_array(5011);
		when "0001001110010100" => data_out <= rom_array(5012);
		when "0001001110010101" => data_out <= rom_array(5013);
		when "0001001110010110" => data_out <= rom_array(5014);
		when "0001001110010111" => data_out <= rom_array(5015);
		when "0001001110011000" => data_out <= rom_array(5016);
		when "0001001110011001" => data_out <= rom_array(5017);
		when "0001001110011010" => data_out <= rom_array(5018);
		when "0001001110011011" => data_out <= rom_array(5019);
		when "0001001110011100" => data_out <= rom_array(5020);
		when "0001001110011101" => data_out <= rom_array(5021);
		when "0001001110011110" => data_out <= rom_array(5022);
		when "0001001110011111" => data_out <= rom_array(5023);
		when "0001001110100000" => data_out <= rom_array(5024);
		when "0001001110100001" => data_out <= rom_array(5025);
		when "0001001110100010" => data_out <= rom_array(5026);
		when "0001001110100011" => data_out <= rom_array(5027);
		when "0001001110100100" => data_out <= rom_array(5028);
		when "0001001110100101" => data_out <= rom_array(5029);
		when "0001001110100110" => data_out <= rom_array(5030);
		when "0001001110100111" => data_out <= rom_array(5031);
		when "0001001110101000" => data_out <= rom_array(5032);
		when "0001001110101001" => data_out <= rom_array(5033);
		when "0001001110101010" => data_out <= rom_array(5034);
		when "0001001110101011" => data_out <= rom_array(5035);
		when "0001001110101100" => data_out <= rom_array(5036);
		when "0001001110101101" => data_out <= rom_array(5037);
		when "0001001110101110" => data_out <= rom_array(5038);
		when "0001001110101111" => data_out <= rom_array(5039);
		when "0001001110110000" => data_out <= rom_array(5040);
		when "0001001110110001" => data_out <= rom_array(5041);
		when "0001001110110010" => data_out <= rom_array(5042);
		when "0001001110110011" => data_out <= rom_array(5043);
		when "0001001110110100" => data_out <= rom_array(5044);
		when "0001001110110101" => data_out <= rom_array(5045);
		when "0001001110110110" => data_out <= rom_array(5046);
		when "0001001110110111" => data_out <= rom_array(5047);
		when "0001001110111000" => data_out <= rom_array(5048);
		when "0001001110111001" => data_out <= rom_array(5049);
		when "0001001110111010" => data_out <= rom_array(5050);
		when "0001001110111011" => data_out <= rom_array(5051);
		when "0001001110111100" => data_out <= rom_array(5052);
		when "0001001110111101" => data_out <= rom_array(5053);
		when "0001001110111110" => data_out <= rom_array(5054);
		when "0001001110111111" => data_out <= rom_array(5055);
		when "0001001111000000" => data_out <= rom_array(5056);
		when "0001001111000001" => data_out <= rom_array(5057);
		when "0001001111000010" => data_out <= rom_array(5058);
		when "0001001111000011" => data_out <= rom_array(5059);
		when "0001001111000100" => data_out <= rom_array(5060);
		when "0001001111000101" => data_out <= rom_array(5061);
		when "0001001111000110" => data_out <= rom_array(5062);
		when "0001001111000111" => data_out <= rom_array(5063);
		when "0001001111001000" => data_out <= rom_array(5064);
		when "0001001111001001" => data_out <= rom_array(5065);
		when "0001001111001010" => data_out <= rom_array(5066);
		when "0001001111001011" => data_out <= rom_array(5067);
		when "0001001111001100" => data_out <= rom_array(5068);
		when "0001001111001101" => data_out <= rom_array(5069);
		when "0001001111001110" => data_out <= rom_array(5070);
		when "0001001111001111" => data_out <= rom_array(5071);
		when "0001001111010000" => data_out <= rom_array(5072);
		when "0001001111010001" => data_out <= rom_array(5073);
		when "0001001111010010" => data_out <= rom_array(5074);
		when "0001001111010011" => data_out <= rom_array(5075);
		when "0001001111010100" => data_out <= rom_array(5076);
		when "0001001111010101" => data_out <= rom_array(5077);
		when "0001001111010110" => data_out <= rom_array(5078);
		when "0001001111010111" => data_out <= rom_array(5079);
		when "0001001111011000" => data_out <= rom_array(5080);
		when "0001001111011001" => data_out <= rom_array(5081);
		when "0001001111011010" => data_out <= rom_array(5082);
		when "0001001111011011" => data_out <= rom_array(5083);
		when "0001001111011100" => data_out <= rom_array(5084);
		when "0001001111011101" => data_out <= rom_array(5085);
		when "0001001111011110" => data_out <= rom_array(5086);
		when "0001001111011111" => data_out <= rom_array(5087);
		when "0001001111100000" => data_out <= rom_array(5088);
		when "0001001111100001" => data_out <= rom_array(5089);
		when "0001001111100010" => data_out <= rom_array(5090);
		when "0001001111100011" => data_out <= rom_array(5091);
		when "0001001111100100" => data_out <= rom_array(5092);
		when "0001001111100101" => data_out <= rom_array(5093);
		when "0001001111100110" => data_out <= rom_array(5094);
		when "0001001111100111" => data_out <= rom_array(5095);
		when "0001001111101000" => data_out <= rom_array(5096);
		when "0001001111101001" => data_out <= rom_array(5097);
		when "0001001111101010" => data_out <= rom_array(5098);
		when "0001001111101011" => data_out <= rom_array(5099);
		when "0001001111101100" => data_out <= rom_array(5100);
		when "0001001111101101" => data_out <= rom_array(5101);
		when "0001001111101110" => data_out <= rom_array(5102);
		when "0001001111101111" => data_out <= rom_array(5103);
		when "0001001111110000" => data_out <= rom_array(5104);
		when "0001001111110001" => data_out <= rom_array(5105);
		when "0001001111110010" => data_out <= rom_array(5106);
		when "0001001111110011" => data_out <= rom_array(5107);
		when "0001001111110100" => data_out <= rom_array(5108);
		when "0001001111110101" => data_out <= rom_array(5109);
		when "0001001111110110" => data_out <= rom_array(5110);
		when "0001001111110111" => data_out <= rom_array(5111);
		when "0001001111111000" => data_out <= rom_array(5112);
		when "0001001111111001" => data_out <= rom_array(5113);
		when "0001001111111010" => data_out <= rom_array(5114);
		when "0001001111111011" => data_out <= rom_array(5115);
		when "0001001111111100" => data_out <= rom_array(5116);
		when "0001001111111101" => data_out <= rom_array(5117);
		when "0001001111111110" => data_out <= rom_array(5118);
		when "0001001111111111" => data_out <= rom_array(5119);
		when "0001010000000000" => data_out <= rom_array(5120);
		when "0001010000000001" => data_out <= rom_array(5121);
		when "0001010000000010" => data_out <= rom_array(5122);
		when "0001010000000011" => data_out <= rom_array(5123);
		when "0001010000000100" => data_out <= rom_array(5124);
		when "0001010000000101" => data_out <= rom_array(5125);
		when "0001010000000110" => data_out <= rom_array(5126);
		when "0001010000000111" => data_out <= rom_array(5127);
		when "0001010000001000" => data_out <= rom_array(5128);
		when "0001010000001001" => data_out <= rom_array(5129);
		when "0001010000001010" => data_out <= rom_array(5130);
		when "0001010000001011" => data_out <= rom_array(5131);
		when "0001010000001100" => data_out <= rom_array(5132);
		when "0001010000001101" => data_out <= rom_array(5133);
		when "0001010000001110" => data_out <= rom_array(5134);
		when "0001010000001111" => data_out <= rom_array(5135);
		when "0001010000010000" => data_out <= rom_array(5136);
		when "0001010000010001" => data_out <= rom_array(5137);
		when "0001010000010010" => data_out <= rom_array(5138);
		when "0001010000010011" => data_out <= rom_array(5139);
		when "0001010000010100" => data_out <= rom_array(5140);
		when "0001010000010101" => data_out <= rom_array(5141);
		when "0001010000010110" => data_out <= rom_array(5142);
		when "0001010000010111" => data_out <= rom_array(5143);
		when "0001010000011000" => data_out <= rom_array(5144);
		when "0001010000011001" => data_out <= rom_array(5145);
		when "0001010000011010" => data_out <= rom_array(5146);
		when "0001010000011011" => data_out <= rom_array(5147);
		when "0001010000011100" => data_out <= rom_array(5148);
		when "0001010000011101" => data_out <= rom_array(5149);
		when "0001010000011110" => data_out <= rom_array(5150);
		when "0001010000011111" => data_out <= rom_array(5151);
		when "0001010000100000" => data_out <= rom_array(5152);
		when "0001010000100001" => data_out <= rom_array(5153);
		when "0001010000100010" => data_out <= rom_array(5154);
		when "0001010000100011" => data_out <= rom_array(5155);
		when "0001010000100100" => data_out <= rom_array(5156);
		when "0001010000100101" => data_out <= rom_array(5157);
		when "0001010000100110" => data_out <= rom_array(5158);
		when "0001010000100111" => data_out <= rom_array(5159);
		when "0001010000101000" => data_out <= rom_array(5160);
		when "0001010000101001" => data_out <= rom_array(5161);
		when "0001010000101010" => data_out <= rom_array(5162);
		when "0001010000101011" => data_out <= rom_array(5163);
		when "0001010000101100" => data_out <= rom_array(5164);
		when "0001010000101101" => data_out <= rom_array(5165);
		when "0001010000101110" => data_out <= rom_array(5166);
		when "0001010000101111" => data_out <= rom_array(5167);
		when "0001010000110000" => data_out <= rom_array(5168);
		when "0001010000110001" => data_out <= rom_array(5169);
		when "0001010000110010" => data_out <= rom_array(5170);
		when "0001010000110011" => data_out <= rom_array(5171);
		when "0001010000110100" => data_out <= rom_array(5172);
		when "0001010000110101" => data_out <= rom_array(5173);
		when "0001010000110110" => data_out <= rom_array(5174);
		when "0001010000110111" => data_out <= rom_array(5175);
		when "0001010000111000" => data_out <= rom_array(5176);
		when "0001010000111001" => data_out <= rom_array(5177);
		when "0001010000111010" => data_out <= rom_array(5178);
		when "0001010000111011" => data_out <= rom_array(5179);
		when "0001010000111100" => data_out <= rom_array(5180);
		when "0001010000111101" => data_out <= rom_array(5181);
		when "0001010000111110" => data_out <= rom_array(5182);
		when "0001010000111111" => data_out <= rom_array(5183);
		when "0001010001000000" => data_out <= rom_array(5184);
		when "0001010001000001" => data_out <= rom_array(5185);
		when "0001010001000010" => data_out <= rom_array(5186);
		when "0001010001000011" => data_out <= rom_array(5187);
		when "0001010001000100" => data_out <= rom_array(5188);
		when "0001010001000101" => data_out <= rom_array(5189);
		when "0001010001000110" => data_out <= rom_array(5190);
		when "0001010001000111" => data_out <= rom_array(5191);
		when "0001010001001000" => data_out <= rom_array(5192);
		when "0001010001001001" => data_out <= rom_array(5193);
		when "0001010001001010" => data_out <= rom_array(5194);
		when "0001010001001011" => data_out <= rom_array(5195);
		when "0001010001001100" => data_out <= rom_array(5196);
		when "0001010001001101" => data_out <= rom_array(5197);
		when "0001010001001110" => data_out <= rom_array(5198);
		when "0001010001001111" => data_out <= rom_array(5199);
		when "0001010001010000" => data_out <= rom_array(5200);
		when "0001010001010001" => data_out <= rom_array(5201);
		when "0001010001010010" => data_out <= rom_array(5202);
		when "0001010001010011" => data_out <= rom_array(5203);
		when "0001010001010100" => data_out <= rom_array(5204);
		when "0001010001010101" => data_out <= rom_array(5205);
		when "0001010001010110" => data_out <= rom_array(5206);
		when "0001010001010111" => data_out <= rom_array(5207);
		when "0001010001011000" => data_out <= rom_array(5208);
		when "0001010001011001" => data_out <= rom_array(5209);
		when "0001010001011010" => data_out <= rom_array(5210);
		when "0001010001011011" => data_out <= rom_array(5211);
		when "0001010001011100" => data_out <= rom_array(5212);
		when "0001010001011101" => data_out <= rom_array(5213);
		when "0001010001011110" => data_out <= rom_array(5214);
		when "0001010001011111" => data_out <= rom_array(5215);
		when "0001010001100000" => data_out <= rom_array(5216);
		when "0001010001100001" => data_out <= rom_array(5217);
		when "0001010001100010" => data_out <= rom_array(5218);
		when "0001010001100011" => data_out <= rom_array(5219);
		when "0001010001100100" => data_out <= rom_array(5220);
		when "0001010001100101" => data_out <= rom_array(5221);
		when "0001010001100110" => data_out <= rom_array(5222);
		when "0001010001100111" => data_out <= rom_array(5223);
		when "0001010001101000" => data_out <= rom_array(5224);
		when "0001010001101001" => data_out <= rom_array(5225);
		when "0001010001101010" => data_out <= rom_array(5226);
		when "0001010001101011" => data_out <= rom_array(5227);
		when "0001010001101100" => data_out <= rom_array(5228);
		when "0001010001101101" => data_out <= rom_array(5229);
		when "0001010001101110" => data_out <= rom_array(5230);
		when "0001010001101111" => data_out <= rom_array(5231);
		when "0001010001110000" => data_out <= rom_array(5232);
		when "0001010001110001" => data_out <= rom_array(5233);
		when "0001010001110010" => data_out <= rom_array(5234);
		when "0001010001110011" => data_out <= rom_array(5235);
		when "0001010001110100" => data_out <= rom_array(5236);
		when "0001010001110101" => data_out <= rom_array(5237);
		when "0001010001110110" => data_out <= rom_array(5238);
		when "0001010001110111" => data_out <= rom_array(5239);
		when "0001010001111000" => data_out <= rom_array(5240);
		when "0001010001111001" => data_out <= rom_array(5241);
		when "0001010001111010" => data_out <= rom_array(5242);
		when "0001010001111011" => data_out <= rom_array(5243);
		when "0001010001111100" => data_out <= rom_array(5244);
		when "0001010001111101" => data_out <= rom_array(5245);
		when "0001010001111110" => data_out <= rom_array(5246);
		when "0001010001111111" => data_out <= rom_array(5247);
		when "0001010010000000" => data_out <= rom_array(5248);
		when "0001010010000001" => data_out <= rom_array(5249);
		when "0001010010000010" => data_out <= rom_array(5250);
		when "0001010010000011" => data_out <= rom_array(5251);
		when "0001010010000100" => data_out <= rom_array(5252);
		when "0001010010000101" => data_out <= rom_array(5253);
		when "0001010010000110" => data_out <= rom_array(5254);
		when "0001010010000111" => data_out <= rom_array(5255);
		when "0001010010001000" => data_out <= rom_array(5256);
		when "0001010010001001" => data_out <= rom_array(5257);
		when "0001010010001010" => data_out <= rom_array(5258);
		when "0001010010001011" => data_out <= rom_array(5259);
		when "0001010010001100" => data_out <= rom_array(5260);
		when "0001010010001101" => data_out <= rom_array(5261);
		when "0001010010001110" => data_out <= rom_array(5262);
		when "0001010010001111" => data_out <= rom_array(5263);
		when "0001010010010000" => data_out <= rom_array(5264);
		when "0001010010010001" => data_out <= rom_array(5265);
		when "0001010010010010" => data_out <= rom_array(5266);
		when "0001010010010011" => data_out <= rom_array(5267);
		when "0001010010010100" => data_out <= rom_array(5268);
		when "0001010010010101" => data_out <= rom_array(5269);
		when "0001010010010110" => data_out <= rom_array(5270);
		when "0001010010010111" => data_out <= rom_array(5271);
		when "0001010010011000" => data_out <= rom_array(5272);
		when "0001010010011001" => data_out <= rom_array(5273);
		when "0001010010011010" => data_out <= rom_array(5274);
		when "0001010010011011" => data_out <= rom_array(5275);
		when "0001010010011100" => data_out <= rom_array(5276);
		when "0001010010011101" => data_out <= rom_array(5277);
		when "0001010010011110" => data_out <= rom_array(5278);
		when "0001010010011111" => data_out <= rom_array(5279);
		when "0001010010100000" => data_out <= rom_array(5280);
		when "0001010010100001" => data_out <= rom_array(5281);
		when "0001010010100010" => data_out <= rom_array(5282);
		when "0001010010100011" => data_out <= rom_array(5283);
		when "0001010010100100" => data_out <= rom_array(5284);
		when "0001010010100101" => data_out <= rom_array(5285);
		when "0001010010100110" => data_out <= rom_array(5286);
		when "0001010010100111" => data_out <= rom_array(5287);
		when "0001010010101000" => data_out <= rom_array(5288);
		when "0001010010101001" => data_out <= rom_array(5289);
		when "0001010010101010" => data_out <= rom_array(5290);
		when "0001010010101011" => data_out <= rom_array(5291);
		when "0001010010101100" => data_out <= rom_array(5292);
		when "0001010010101101" => data_out <= rom_array(5293);
		when "0001010010101110" => data_out <= rom_array(5294);
		when "0001010010101111" => data_out <= rom_array(5295);
		when "0001010010110000" => data_out <= rom_array(5296);
		when "0001010010110001" => data_out <= rom_array(5297);
		when "0001010010110010" => data_out <= rom_array(5298);
		when "0001010010110011" => data_out <= rom_array(5299);
		when "0001010010110100" => data_out <= rom_array(5300);
		when "0001010010110101" => data_out <= rom_array(5301);
		when "0001010010110110" => data_out <= rom_array(5302);
		when "0001010010110111" => data_out <= rom_array(5303);
		when "0001010010111000" => data_out <= rom_array(5304);
		when "0001010010111001" => data_out <= rom_array(5305);
		when "0001010010111010" => data_out <= rom_array(5306);
		when "0001010010111011" => data_out <= rom_array(5307);
		when "0001010010111100" => data_out <= rom_array(5308);
		when "0001010010111101" => data_out <= rom_array(5309);
		when "0001010010111110" => data_out <= rom_array(5310);
		when "0001010010111111" => data_out <= rom_array(5311);
		when "0001010011000000" => data_out <= rom_array(5312);
		when "0001010011000001" => data_out <= rom_array(5313);
		when "0001010011000010" => data_out <= rom_array(5314);
		when "0001010011000011" => data_out <= rom_array(5315);
		when "0001010011000100" => data_out <= rom_array(5316);
		when "0001010011000101" => data_out <= rom_array(5317);
		when "0001010011000110" => data_out <= rom_array(5318);
		when "0001010011000111" => data_out <= rom_array(5319);
		when "0001010011001000" => data_out <= rom_array(5320);
		when "0001010011001001" => data_out <= rom_array(5321);
		when "0001010011001010" => data_out <= rom_array(5322);
		when "0001010011001011" => data_out <= rom_array(5323);
		when "0001010011001100" => data_out <= rom_array(5324);
		when "0001010011001101" => data_out <= rom_array(5325);
		when "0001010011001110" => data_out <= rom_array(5326);
		when "0001010011001111" => data_out <= rom_array(5327);
		when "0001010011010000" => data_out <= rom_array(5328);
		when "0001010011010001" => data_out <= rom_array(5329);
		when "0001010011010010" => data_out <= rom_array(5330);
		when "0001010011010011" => data_out <= rom_array(5331);
		when "0001010011010100" => data_out <= rom_array(5332);
		when "0001010011010101" => data_out <= rom_array(5333);
		when "0001010011010110" => data_out <= rom_array(5334);
		when "0001010011010111" => data_out <= rom_array(5335);
		when "0001010011011000" => data_out <= rom_array(5336);
		when "0001010011011001" => data_out <= rom_array(5337);
		when "0001010011011010" => data_out <= rom_array(5338);
		when "0001010011011011" => data_out <= rom_array(5339);
		when "0001010011011100" => data_out <= rom_array(5340);
		when "0001010011011101" => data_out <= rom_array(5341);
		when "0001010011011110" => data_out <= rom_array(5342);
		when "0001010011011111" => data_out <= rom_array(5343);
		when "0001010011100000" => data_out <= rom_array(5344);
		when "0001010011100001" => data_out <= rom_array(5345);
		when "0001010011100010" => data_out <= rom_array(5346);
		when "0001010011100011" => data_out <= rom_array(5347);
		when "0001010011100100" => data_out <= rom_array(5348);
		when "0001010011100101" => data_out <= rom_array(5349);
		when "0001010011100110" => data_out <= rom_array(5350);
		when "0001010011100111" => data_out <= rom_array(5351);
		when "0001010011101000" => data_out <= rom_array(5352);
		when "0001010011101001" => data_out <= rom_array(5353);
		when "0001010011101010" => data_out <= rom_array(5354);
		when "0001010011101011" => data_out <= rom_array(5355);
		when "0001010011101100" => data_out <= rom_array(5356);
		when "0001010011101101" => data_out <= rom_array(5357);
		when "0001010011101110" => data_out <= rom_array(5358);
		when "0001010011101111" => data_out <= rom_array(5359);
		when "0001010011110000" => data_out <= rom_array(5360);
		when "0001010011110001" => data_out <= rom_array(5361);
		when "0001010011110010" => data_out <= rom_array(5362);
		when "0001010011110011" => data_out <= rom_array(5363);
		when "0001010011110100" => data_out <= rom_array(5364);
		when "0001010011110101" => data_out <= rom_array(5365);
		when "0001010011110110" => data_out <= rom_array(5366);
		when "0001010011110111" => data_out <= rom_array(5367);
		when "0001010011111000" => data_out <= rom_array(5368);
		when "0001010011111001" => data_out <= rom_array(5369);
		when "0001010011111010" => data_out <= rom_array(5370);
		when "0001010011111011" => data_out <= rom_array(5371);
		when "0001010011111100" => data_out <= rom_array(5372);
		when "0001010011111101" => data_out <= rom_array(5373);
		when "0001010011111110" => data_out <= rom_array(5374);
		when "0001010011111111" => data_out <= rom_array(5375);
		when "0001010100000000" => data_out <= rom_array(5376);
		when "0001010100000001" => data_out <= rom_array(5377);
		when "0001010100000010" => data_out <= rom_array(5378);
		when "0001010100000011" => data_out <= rom_array(5379);
		when "0001010100000100" => data_out <= rom_array(5380);
		when "0001010100000101" => data_out <= rom_array(5381);
		when "0001010100000110" => data_out <= rom_array(5382);
		when "0001010100000111" => data_out <= rom_array(5383);
		when "0001010100001000" => data_out <= rom_array(5384);
		when "0001010100001001" => data_out <= rom_array(5385);
		when "0001010100001010" => data_out <= rom_array(5386);
		when "0001010100001011" => data_out <= rom_array(5387);
		when "0001010100001100" => data_out <= rom_array(5388);
		when "0001010100001101" => data_out <= rom_array(5389);
		when "0001010100001110" => data_out <= rom_array(5390);
		when "0001010100001111" => data_out <= rom_array(5391);
		when "0001010100010000" => data_out <= rom_array(5392);
		when "0001010100010001" => data_out <= rom_array(5393);
		when "0001010100010010" => data_out <= rom_array(5394);
		when "0001010100010011" => data_out <= rom_array(5395);
		when "0001010100010100" => data_out <= rom_array(5396);
		when "0001010100010101" => data_out <= rom_array(5397);
		when "0001010100010110" => data_out <= rom_array(5398);
		when "0001010100010111" => data_out <= rom_array(5399);
		when "0001010100011000" => data_out <= rom_array(5400);
		when "0001010100011001" => data_out <= rom_array(5401);
		when "0001010100011010" => data_out <= rom_array(5402);
		when "0001010100011011" => data_out <= rom_array(5403);
		when "0001010100011100" => data_out <= rom_array(5404);
		when "0001010100011101" => data_out <= rom_array(5405);
		when "0001010100011110" => data_out <= rom_array(5406);
		when "0001010100011111" => data_out <= rom_array(5407);
		when "0001010100100000" => data_out <= rom_array(5408);
		when "0001010100100001" => data_out <= rom_array(5409);
		when "0001010100100010" => data_out <= rom_array(5410);
		when "0001010100100011" => data_out <= rom_array(5411);
		when "0001010100100100" => data_out <= rom_array(5412);
		when "0001010100100101" => data_out <= rom_array(5413);
		when "0001010100100110" => data_out <= rom_array(5414);
		when "0001010100100111" => data_out <= rom_array(5415);
		when "0001010100101000" => data_out <= rom_array(5416);
		when "0001010100101001" => data_out <= rom_array(5417);
		when "0001010100101010" => data_out <= rom_array(5418);
		when "0001010100101011" => data_out <= rom_array(5419);
		when "0001010100101100" => data_out <= rom_array(5420);
		when "0001010100101101" => data_out <= rom_array(5421);
		when "0001010100101110" => data_out <= rom_array(5422);
		when "0001010100101111" => data_out <= rom_array(5423);
		when "0001010100110000" => data_out <= rom_array(5424);
		when "0001010100110001" => data_out <= rom_array(5425);
		when "0001010100110010" => data_out <= rom_array(5426);
		when "0001010100110011" => data_out <= rom_array(5427);
		when "0001010100110100" => data_out <= rom_array(5428);
		when "0001010100110101" => data_out <= rom_array(5429);
		when "0001010100110110" => data_out <= rom_array(5430);
		when "0001010100110111" => data_out <= rom_array(5431);
		when "0001010100111000" => data_out <= rom_array(5432);
		when "0001010100111001" => data_out <= rom_array(5433);
		when "0001010100111010" => data_out <= rom_array(5434);
		when "0001010100111011" => data_out <= rom_array(5435);
		when "0001010100111100" => data_out <= rom_array(5436);
		when "0001010100111101" => data_out <= rom_array(5437);
		when "0001010100111110" => data_out <= rom_array(5438);
		when "0001010100111111" => data_out <= rom_array(5439);
		when "0001010101000000" => data_out <= rom_array(5440);
		when "0001010101000001" => data_out <= rom_array(5441);
		when "0001010101000010" => data_out <= rom_array(5442);
		when "0001010101000011" => data_out <= rom_array(5443);
		when "0001010101000100" => data_out <= rom_array(5444);
		when "0001010101000101" => data_out <= rom_array(5445);
		when "0001010101000110" => data_out <= rom_array(5446);
		when "0001010101000111" => data_out <= rom_array(5447);
		when "0001010101001000" => data_out <= rom_array(5448);
		when "0001010101001001" => data_out <= rom_array(5449);
		when "0001010101001010" => data_out <= rom_array(5450);
		when "0001010101001011" => data_out <= rom_array(5451);
		when "0001010101001100" => data_out <= rom_array(5452);
		when "0001010101001101" => data_out <= rom_array(5453);
		when "0001010101001110" => data_out <= rom_array(5454);
		when "0001010101001111" => data_out <= rom_array(5455);
		when "0001010101010000" => data_out <= rom_array(5456);
		when "0001010101010001" => data_out <= rom_array(5457);
		when "0001010101010010" => data_out <= rom_array(5458);
		when "0001010101010011" => data_out <= rom_array(5459);
		when "0001010101010100" => data_out <= rom_array(5460);
		when "0001010101010101" => data_out <= rom_array(5461);
		when "0001010101010110" => data_out <= rom_array(5462);
		when "0001010101010111" => data_out <= rom_array(5463);
		when "0001010101011000" => data_out <= rom_array(5464);
		when "0001010101011001" => data_out <= rom_array(5465);
		when "0001010101011010" => data_out <= rom_array(5466);
		when "0001010101011011" => data_out <= rom_array(5467);
		when "0001010101011100" => data_out <= rom_array(5468);
		when "0001010101011101" => data_out <= rom_array(5469);
		when "0001010101011110" => data_out <= rom_array(5470);
		when "0001010101011111" => data_out <= rom_array(5471);
		when "0001010101100000" => data_out <= rom_array(5472);
		when "0001010101100001" => data_out <= rom_array(5473);
		when "0001010101100010" => data_out <= rom_array(5474);
		when "0001010101100011" => data_out <= rom_array(5475);
		when "0001010101100100" => data_out <= rom_array(5476);
		when "0001010101100101" => data_out <= rom_array(5477);
		when "0001010101100110" => data_out <= rom_array(5478);
		when "0001010101100111" => data_out <= rom_array(5479);
		when "0001010101101000" => data_out <= rom_array(5480);
		when "0001010101101001" => data_out <= rom_array(5481);
		when "0001010101101010" => data_out <= rom_array(5482);
		when "0001010101101011" => data_out <= rom_array(5483);
		when "0001010101101100" => data_out <= rom_array(5484);
		when "0001010101101101" => data_out <= rom_array(5485);
		when "0001010101101110" => data_out <= rom_array(5486);
		when "0001010101101111" => data_out <= rom_array(5487);
		when "0001010101110000" => data_out <= rom_array(5488);
		when "0001010101110001" => data_out <= rom_array(5489);
		when "0001010101110010" => data_out <= rom_array(5490);
		when "0001010101110011" => data_out <= rom_array(5491);
		when "0001010101110100" => data_out <= rom_array(5492);
		when "0001010101110101" => data_out <= rom_array(5493);
		when "0001010101110110" => data_out <= rom_array(5494);
		when "0001010101110111" => data_out <= rom_array(5495);
		when "0001010101111000" => data_out <= rom_array(5496);
		when "0001010101111001" => data_out <= rom_array(5497);
		when "0001010101111010" => data_out <= rom_array(5498);
		when "0001010101111011" => data_out <= rom_array(5499);
		when "0001010101111100" => data_out <= rom_array(5500);
		when "0001010101111101" => data_out <= rom_array(5501);
		when "0001010101111110" => data_out <= rom_array(5502);
		when "0001010101111111" => data_out <= rom_array(5503);
		when "0001010110000000" => data_out <= rom_array(5504);
		when "0001010110000001" => data_out <= rom_array(5505);
		when "0001010110000010" => data_out <= rom_array(5506);
		when "0001010110000011" => data_out <= rom_array(5507);
		when "0001010110000100" => data_out <= rom_array(5508);
		when "0001010110000101" => data_out <= rom_array(5509);
		when "0001010110000110" => data_out <= rom_array(5510);
		when "0001010110000111" => data_out <= rom_array(5511);
		when "0001010110001000" => data_out <= rom_array(5512);
		when "0001010110001001" => data_out <= rom_array(5513);
		when "0001010110001010" => data_out <= rom_array(5514);
		when "0001010110001011" => data_out <= rom_array(5515);
		when "0001010110001100" => data_out <= rom_array(5516);
		when "0001010110001101" => data_out <= rom_array(5517);
		when "0001010110001110" => data_out <= rom_array(5518);
		when "0001010110001111" => data_out <= rom_array(5519);
		when "0001010110010000" => data_out <= rom_array(5520);
		when "0001010110010001" => data_out <= rom_array(5521);
		when "0001010110010010" => data_out <= rom_array(5522);
		when "0001010110010011" => data_out <= rom_array(5523);
		when "0001010110010100" => data_out <= rom_array(5524);
		when "0001010110010101" => data_out <= rom_array(5525);
		when "0001010110010110" => data_out <= rom_array(5526);
		when "0001010110010111" => data_out <= rom_array(5527);
		when "0001010110011000" => data_out <= rom_array(5528);
		when "0001010110011001" => data_out <= rom_array(5529);
		when "0001010110011010" => data_out <= rom_array(5530);
		when "0001010110011011" => data_out <= rom_array(5531);
		when "0001010110011100" => data_out <= rom_array(5532);
		when "0001010110011101" => data_out <= rom_array(5533);
		when "0001010110011110" => data_out <= rom_array(5534);
		when "0001010110011111" => data_out <= rom_array(5535);
		when "0001010110100000" => data_out <= rom_array(5536);
		when "0001010110100001" => data_out <= rom_array(5537);
		when "0001010110100010" => data_out <= rom_array(5538);
		when "0001010110100011" => data_out <= rom_array(5539);
		when "0001010110100100" => data_out <= rom_array(5540);
		when "0001010110100101" => data_out <= rom_array(5541);
		when "0001010110100110" => data_out <= rom_array(5542);
		when "0001010110100111" => data_out <= rom_array(5543);
		when "0001010110101000" => data_out <= rom_array(5544);
		when "0001010110101001" => data_out <= rom_array(5545);
		when "0001010110101010" => data_out <= rom_array(5546);
		when "0001010110101011" => data_out <= rom_array(5547);
		when "0001010110101100" => data_out <= rom_array(5548);
		when "0001010110101101" => data_out <= rom_array(5549);
		when "0001010110101110" => data_out <= rom_array(5550);
		when "0001010110101111" => data_out <= rom_array(5551);
		when "0001010110110000" => data_out <= rom_array(5552);
		when "0001010110110001" => data_out <= rom_array(5553);
		when "0001010110110010" => data_out <= rom_array(5554);
		when "0001010110110011" => data_out <= rom_array(5555);
		when "0001010110110100" => data_out <= rom_array(5556);
		when "0001010110110101" => data_out <= rom_array(5557);
		when "0001010110110110" => data_out <= rom_array(5558);
		when "0001010110110111" => data_out <= rom_array(5559);
		when "0001010110111000" => data_out <= rom_array(5560);
		when "0001010110111001" => data_out <= rom_array(5561);
		when "0001010110111010" => data_out <= rom_array(5562);
		when "0001010110111011" => data_out <= rom_array(5563);
		when "0001010110111100" => data_out <= rom_array(5564);
		when "0001010110111101" => data_out <= rom_array(5565);
		when "0001010110111110" => data_out <= rom_array(5566);
		when "0001010110111111" => data_out <= rom_array(5567);
		when "0001010111000000" => data_out <= rom_array(5568);
		when "0001010111000001" => data_out <= rom_array(5569);
		when "0001010111000010" => data_out <= rom_array(5570);
		when "0001010111000011" => data_out <= rom_array(5571);
		when "0001010111000100" => data_out <= rom_array(5572);
		when "0001010111000101" => data_out <= rom_array(5573);
		when "0001010111000110" => data_out <= rom_array(5574);
		when "0001010111000111" => data_out <= rom_array(5575);
		when "0001010111001000" => data_out <= rom_array(5576);
		when "0001010111001001" => data_out <= rom_array(5577);
		when "0001010111001010" => data_out <= rom_array(5578);
		when "0001010111001011" => data_out <= rom_array(5579);
		when "0001010111001100" => data_out <= rom_array(5580);
		when "0001010111001101" => data_out <= rom_array(5581);
		when "0001010111001110" => data_out <= rom_array(5582);
		when "0001010111001111" => data_out <= rom_array(5583);
		when "0001010111010000" => data_out <= rom_array(5584);
		when "0001010111010001" => data_out <= rom_array(5585);
		when "0001010111010010" => data_out <= rom_array(5586);
		when "0001010111010011" => data_out <= rom_array(5587);
		when "0001010111010100" => data_out <= rom_array(5588);
		when "0001010111010101" => data_out <= rom_array(5589);
		when "0001010111010110" => data_out <= rom_array(5590);
		when "0001010111010111" => data_out <= rom_array(5591);
		when "0001010111011000" => data_out <= rom_array(5592);
		when "0001010111011001" => data_out <= rom_array(5593);
		when "0001010111011010" => data_out <= rom_array(5594);
		when "0001010111011011" => data_out <= rom_array(5595);
		when "0001010111011100" => data_out <= rom_array(5596);
		when "0001010111011101" => data_out <= rom_array(5597);
		when "0001010111011110" => data_out <= rom_array(5598);
		when "0001010111011111" => data_out <= rom_array(5599);
		when "0001010111100000" => data_out <= rom_array(5600);
		when "0001010111100001" => data_out <= rom_array(5601);
		when "0001010111100010" => data_out <= rom_array(5602);
		when "0001010111100011" => data_out <= rom_array(5603);
		when "0001010111100100" => data_out <= rom_array(5604);
		when "0001010111100101" => data_out <= rom_array(5605);
		when "0001010111100110" => data_out <= rom_array(5606);
		when "0001010111100111" => data_out <= rom_array(5607);
		when "0001010111101000" => data_out <= rom_array(5608);
		when "0001010111101001" => data_out <= rom_array(5609);
		when "0001010111101010" => data_out <= rom_array(5610);
		when "0001010111101011" => data_out <= rom_array(5611);
		when "0001010111101100" => data_out <= rom_array(5612);
		when "0001010111101101" => data_out <= rom_array(5613);
		when "0001010111101110" => data_out <= rom_array(5614);
		when "0001010111101111" => data_out <= rom_array(5615);
		when "0001010111110000" => data_out <= rom_array(5616);
		when "0001010111110001" => data_out <= rom_array(5617);
		when "0001010111110010" => data_out <= rom_array(5618);
		when "0001010111110011" => data_out <= rom_array(5619);
		when "0001010111110100" => data_out <= rom_array(5620);
		when "0001010111110101" => data_out <= rom_array(5621);
		when "0001010111110110" => data_out <= rom_array(5622);
		when "0001010111110111" => data_out <= rom_array(5623);
		when "0001010111111000" => data_out <= rom_array(5624);
		when "0001010111111001" => data_out <= rom_array(5625);
		when "0001010111111010" => data_out <= rom_array(5626);
		when "0001010111111011" => data_out <= rom_array(5627);
		when "0001010111111100" => data_out <= rom_array(5628);
		when "0001010111111101" => data_out <= rom_array(5629);
		when "0001010111111110" => data_out <= rom_array(5630);
		when "0001010111111111" => data_out <= rom_array(5631);
		when "0001011000000000" => data_out <= rom_array(5632);
		when "0001011000000001" => data_out <= rom_array(5633);
		when "0001011000000010" => data_out <= rom_array(5634);
		when "0001011000000011" => data_out <= rom_array(5635);
		when "0001011000000100" => data_out <= rom_array(5636);
		when "0001011000000101" => data_out <= rom_array(5637);
		when "0001011000000110" => data_out <= rom_array(5638);
		when "0001011000000111" => data_out <= rom_array(5639);
		when "0001011000001000" => data_out <= rom_array(5640);
		when "0001011000001001" => data_out <= rom_array(5641);
		when "0001011000001010" => data_out <= rom_array(5642);
		when "0001011000001011" => data_out <= rom_array(5643);
		when "0001011000001100" => data_out <= rom_array(5644);
		when "0001011000001101" => data_out <= rom_array(5645);
		when "0001011000001110" => data_out <= rom_array(5646);
		when "0001011000001111" => data_out <= rom_array(5647);
		when "0001011000010000" => data_out <= rom_array(5648);
		when "0001011000010001" => data_out <= rom_array(5649);
		when "0001011000010010" => data_out <= rom_array(5650);
		when "0001011000010011" => data_out <= rom_array(5651);
		when "0001011000010100" => data_out <= rom_array(5652);
		when "0001011000010101" => data_out <= rom_array(5653);
		when "0001011000010110" => data_out <= rom_array(5654);
		when "0001011000010111" => data_out <= rom_array(5655);
		when "0001011000011000" => data_out <= rom_array(5656);
		when "0001011000011001" => data_out <= rom_array(5657);
		when "0001011000011010" => data_out <= rom_array(5658);
		when "0001011000011011" => data_out <= rom_array(5659);
		when "0001011000011100" => data_out <= rom_array(5660);
		when "0001011000011101" => data_out <= rom_array(5661);
		when "0001011000011110" => data_out <= rom_array(5662);
		when "0001011000011111" => data_out <= rom_array(5663);
		when "0001011000100000" => data_out <= rom_array(5664);
		when "0001011000100001" => data_out <= rom_array(5665);
		when "0001011000100010" => data_out <= rom_array(5666);
		when "0001011000100011" => data_out <= rom_array(5667);
		when "0001011000100100" => data_out <= rom_array(5668);
		when "0001011000100101" => data_out <= rom_array(5669);
		when "0001011000100110" => data_out <= rom_array(5670);
		when "0001011000100111" => data_out <= rom_array(5671);
		when "0001011000101000" => data_out <= rom_array(5672);
		when "0001011000101001" => data_out <= rom_array(5673);
		when "0001011000101010" => data_out <= rom_array(5674);
		when "0001011000101011" => data_out <= rom_array(5675);
		when "0001011000101100" => data_out <= rom_array(5676);
		when "0001011000101101" => data_out <= rom_array(5677);
		when "0001011000101110" => data_out <= rom_array(5678);
		when "0001011000101111" => data_out <= rom_array(5679);
		when "0001011000110000" => data_out <= rom_array(5680);
		when "0001011000110001" => data_out <= rom_array(5681);
		when "0001011000110010" => data_out <= rom_array(5682);
		when "0001011000110011" => data_out <= rom_array(5683);
		when "0001011000110100" => data_out <= rom_array(5684);
		when "0001011000110101" => data_out <= rom_array(5685);
		when "0001011000110110" => data_out <= rom_array(5686);
		when "0001011000110111" => data_out <= rom_array(5687);
		when "0001011000111000" => data_out <= rom_array(5688);
		when "0001011000111001" => data_out <= rom_array(5689);
		when "0001011000111010" => data_out <= rom_array(5690);
		when "0001011000111011" => data_out <= rom_array(5691);
		when "0001011000111100" => data_out <= rom_array(5692);
		when "0001011000111101" => data_out <= rom_array(5693);
		when "0001011000111110" => data_out <= rom_array(5694);
		when "0001011000111111" => data_out <= rom_array(5695);
		when "0001011001000000" => data_out <= rom_array(5696);
		when "0001011001000001" => data_out <= rom_array(5697);
		when "0001011001000010" => data_out <= rom_array(5698);
		when "0001011001000011" => data_out <= rom_array(5699);
		when "0001011001000100" => data_out <= rom_array(5700);
		when "0001011001000101" => data_out <= rom_array(5701);
		when "0001011001000110" => data_out <= rom_array(5702);
		when "0001011001000111" => data_out <= rom_array(5703);
		when "0001011001001000" => data_out <= rom_array(5704);
		when "0001011001001001" => data_out <= rom_array(5705);
		when "0001011001001010" => data_out <= rom_array(5706);
		when "0001011001001011" => data_out <= rom_array(5707);
		when "0001011001001100" => data_out <= rom_array(5708);
		when "0001011001001101" => data_out <= rom_array(5709);
		when "0001011001001110" => data_out <= rom_array(5710);
		when "0001011001001111" => data_out <= rom_array(5711);
		when "0001011001010000" => data_out <= rom_array(5712);
		when "0001011001010001" => data_out <= rom_array(5713);
		when "0001011001010010" => data_out <= rom_array(5714);
		when "0001011001010011" => data_out <= rom_array(5715);
		when "0001011001010100" => data_out <= rom_array(5716);
		when "0001011001010101" => data_out <= rom_array(5717);
		when "0001011001010110" => data_out <= rom_array(5718);
		when "0001011001010111" => data_out <= rom_array(5719);
		when "0001011001011000" => data_out <= rom_array(5720);
		when "0001011001011001" => data_out <= rom_array(5721);
		when "0001011001011010" => data_out <= rom_array(5722);
		when "0001011001011011" => data_out <= rom_array(5723);
		when "0001011001011100" => data_out <= rom_array(5724);
		when "0001011001011101" => data_out <= rom_array(5725);
		when "0001011001011110" => data_out <= rom_array(5726);
		when "0001011001011111" => data_out <= rom_array(5727);
		when "0001011001100000" => data_out <= rom_array(5728);
		when "0001011001100001" => data_out <= rom_array(5729);
		when "0001011001100010" => data_out <= rom_array(5730);
		when "0001011001100011" => data_out <= rom_array(5731);
		when "0001011001100100" => data_out <= rom_array(5732);
		when "0001011001100101" => data_out <= rom_array(5733);
		when "0001011001100110" => data_out <= rom_array(5734);
		when "0001011001100111" => data_out <= rom_array(5735);
		when "0001011001101000" => data_out <= rom_array(5736);
		when "0001011001101001" => data_out <= rom_array(5737);
		when "0001011001101010" => data_out <= rom_array(5738);
		when "0001011001101011" => data_out <= rom_array(5739);
		when "0001011001101100" => data_out <= rom_array(5740);
		when "0001011001101101" => data_out <= rom_array(5741);
		when "0001011001101110" => data_out <= rom_array(5742);
		when "0001011001101111" => data_out <= rom_array(5743);
		when "0001011001110000" => data_out <= rom_array(5744);
		when "0001011001110001" => data_out <= rom_array(5745);
		when "0001011001110010" => data_out <= rom_array(5746);
		when "0001011001110011" => data_out <= rom_array(5747);
		when "0001011001110100" => data_out <= rom_array(5748);
		when "0001011001110101" => data_out <= rom_array(5749);
		when "0001011001110110" => data_out <= rom_array(5750);
		when "0001011001110111" => data_out <= rom_array(5751);
		when "0001011001111000" => data_out <= rom_array(5752);
		when "0001011001111001" => data_out <= rom_array(5753);
		when "0001011001111010" => data_out <= rom_array(5754);
		when "0001011001111011" => data_out <= rom_array(5755);
		when "0001011001111100" => data_out <= rom_array(5756);
		when "0001011001111101" => data_out <= rom_array(5757);
		when "0001011001111110" => data_out <= rom_array(5758);
		when "0001011001111111" => data_out <= rom_array(5759);
		when "0001011010000000" => data_out <= rom_array(5760);
		when "0001011010000001" => data_out <= rom_array(5761);
		when "0001011010000010" => data_out <= rom_array(5762);
		when "0001011010000011" => data_out <= rom_array(5763);
		when "0001011010000100" => data_out <= rom_array(5764);
		when "0001011010000101" => data_out <= rom_array(5765);
		when "0001011010000110" => data_out <= rom_array(5766);
		when "0001011010000111" => data_out <= rom_array(5767);
		when "0001011010001000" => data_out <= rom_array(5768);
		when "0001011010001001" => data_out <= rom_array(5769);
		when "0001011010001010" => data_out <= rom_array(5770);
		when "0001011010001011" => data_out <= rom_array(5771);
		when "0001011010001100" => data_out <= rom_array(5772);
		when "0001011010001101" => data_out <= rom_array(5773);
		when "0001011010001110" => data_out <= rom_array(5774);
		when "0001011010001111" => data_out <= rom_array(5775);
		when "0001011010010000" => data_out <= rom_array(5776);
		when "0001011010010001" => data_out <= rom_array(5777);
		when "0001011010010010" => data_out <= rom_array(5778);
		when "0001011010010011" => data_out <= rom_array(5779);
		when "0001011010010100" => data_out <= rom_array(5780);
		when "0001011010010101" => data_out <= rom_array(5781);
		when "0001011010010110" => data_out <= rom_array(5782);
		when "0001011010010111" => data_out <= rom_array(5783);
		when "0001011010011000" => data_out <= rom_array(5784);
		when "0001011010011001" => data_out <= rom_array(5785);
		when "0001011010011010" => data_out <= rom_array(5786);
		when "0001011010011011" => data_out <= rom_array(5787);
		when "0001011010011100" => data_out <= rom_array(5788);
		when "0001011010011101" => data_out <= rom_array(5789);
		when "0001011010011110" => data_out <= rom_array(5790);
		when "0001011010011111" => data_out <= rom_array(5791);
		when "0001011010100000" => data_out <= rom_array(5792);
		when "0001011010100001" => data_out <= rom_array(5793);
		when "0001011010100010" => data_out <= rom_array(5794);
		when "0001011010100011" => data_out <= rom_array(5795);
		when "0001011010100100" => data_out <= rom_array(5796);
		when "0001011010100101" => data_out <= rom_array(5797);
		when "0001011010100110" => data_out <= rom_array(5798);
		when "0001011010100111" => data_out <= rom_array(5799);
		when "0001011010101000" => data_out <= rom_array(5800);
		when "0001011010101001" => data_out <= rom_array(5801);
		when "0001011010101010" => data_out <= rom_array(5802);
		when "0001011010101011" => data_out <= rom_array(5803);
		when "0001011010101100" => data_out <= rom_array(5804);
		when "0001011010101101" => data_out <= rom_array(5805);
		when "0001011010101110" => data_out <= rom_array(5806);
		when "0001011010101111" => data_out <= rom_array(5807);
		when "0001011010110000" => data_out <= rom_array(5808);
		when "0001011010110001" => data_out <= rom_array(5809);
		when "0001011010110010" => data_out <= rom_array(5810);
		when "0001011010110011" => data_out <= rom_array(5811);
		when "0001011010110100" => data_out <= rom_array(5812);
		when "0001011010110101" => data_out <= rom_array(5813);
		when "0001011010110110" => data_out <= rom_array(5814);
		when "0001011010110111" => data_out <= rom_array(5815);
		when "0001011010111000" => data_out <= rom_array(5816);
		when "0001011010111001" => data_out <= rom_array(5817);
		when "0001011010111010" => data_out <= rom_array(5818);
		when "0001011010111011" => data_out <= rom_array(5819);
		when "0001011010111100" => data_out <= rom_array(5820);
		when "0001011010111101" => data_out <= rom_array(5821);
		when "0001011010111110" => data_out <= rom_array(5822);
		when "0001011010111111" => data_out <= rom_array(5823);
		when "0001011011000000" => data_out <= rom_array(5824);
		when "0001011011000001" => data_out <= rom_array(5825);
		when "0001011011000010" => data_out <= rom_array(5826);
		when "0001011011000011" => data_out <= rom_array(5827);
		when "0001011011000100" => data_out <= rom_array(5828);
		when "0001011011000101" => data_out <= rom_array(5829);
		when "0001011011000110" => data_out <= rom_array(5830);
		when "0001011011000111" => data_out <= rom_array(5831);
		when "0001011011001000" => data_out <= rom_array(5832);
		when "0001011011001001" => data_out <= rom_array(5833);
		when "0001011011001010" => data_out <= rom_array(5834);
		when "0001011011001011" => data_out <= rom_array(5835);
		when "0001011011001100" => data_out <= rom_array(5836);
		when "0001011011001101" => data_out <= rom_array(5837);
		when "0001011011001110" => data_out <= rom_array(5838);
		when "0001011011001111" => data_out <= rom_array(5839);
		when "0001011011010000" => data_out <= rom_array(5840);
		when "0001011011010001" => data_out <= rom_array(5841);
		when "0001011011010010" => data_out <= rom_array(5842);
		when "0001011011010011" => data_out <= rom_array(5843);
		when "0001011011010100" => data_out <= rom_array(5844);
		when "0001011011010101" => data_out <= rom_array(5845);
		when "0001011011010110" => data_out <= rom_array(5846);
		when "0001011011010111" => data_out <= rom_array(5847);
		when "0001011011011000" => data_out <= rom_array(5848);
		when "0001011011011001" => data_out <= rom_array(5849);
		when "0001011011011010" => data_out <= rom_array(5850);
		when "0001011011011011" => data_out <= rom_array(5851);
		when "0001011011011100" => data_out <= rom_array(5852);
		when "0001011011011101" => data_out <= rom_array(5853);
		when "0001011011011110" => data_out <= rom_array(5854);
		when "0001011011011111" => data_out <= rom_array(5855);
		when "0001011011100000" => data_out <= rom_array(5856);
		when "0001011011100001" => data_out <= rom_array(5857);
		when "0001011011100010" => data_out <= rom_array(5858);
		when "0001011011100011" => data_out <= rom_array(5859);
		when "0001011011100100" => data_out <= rom_array(5860);
		when "0001011011100101" => data_out <= rom_array(5861);
		when "0001011011100110" => data_out <= rom_array(5862);
		when "0001011011100111" => data_out <= rom_array(5863);
		when "0001011011101000" => data_out <= rom_array(5864);
		when "0001011011101001" => data_out <= rom_array(5865);
		when "0001011011101010" => data_out <= rom_array(5866);
		when "0001011011101011" => data_out <= rom_array(5867);
		when "0001011011101100" => data_out <= rom_array(5868);
		when "0001011011101101" => data_out <= rom_array(5869);
		when "0001011011101110" => data_out <= rom_array(5870);
		when "0001011011101111" => data_out <= rom_array(5871);
		when "0001011011110000" => data_out <= rom_array(5872);
		when "0001011011110001" => data_out <= rom_array(5873);
		when "0001011011110010" => data_out <= rom_array(5874);
		when "0001011011110011" => data_out <= rom_array(5875);
		when "0001011011110100" => data_out <= rom_array(5876);
		when "0001011011110101" => data_out <= rom_array(5877);
		when "0001011011110110" => data_out <= rom_array(5878);
		when "0001011011110111" => data_out <= rom_array(5879);
		when "0001011011111000" => data_out <= rom_array(5880);
		when "0001011011111001" => data_out <= rom_array(5881);
		when "0001011011111010" => data_out <= rom_array(5882);
		when "0001011011111011" => data_out <= rom_array(5883);
		when "0001011011111100" => data_out <= rom_array(5884);
		when "0001011011111101" => data_out <= rom_array(5885);
		when "0001011011111110" => data_out <= rom_array(5886);
		when "0001011011111111" => data_out <= rom_array(5887);
		when "0001011100000000" => data_out <= rom_array(5888);
		when "0001011100000001" => data_out <= rom_array(5889);
		when "0001011100000010" => data_out <= rom_array(5890);
		when "0001011100000011" => data_out <= rom_array(5891);
		when "0001011100000100" => data_out <= rom_array(5892);
		when "0001011100000101" => data_out <= rom_array(5893);
		when "0001011100000110" => data_out <= rom_array(5894);
		when "0001011100000111" => data_out <= rom_array(5895);
		when "0001011100001000" => data_out <= rom_array(5896);
		when "0001011100001001" => data_out <= rom_array(5897);
		when "0001011100001010" => data_out <= rom_array(5898);
		when "0001011100001011" => data_out <= rom_array(5899);
		when "0001011100001100" => data_out <= rom_array(5900);
		when "0001011100001101" => data_out <= rom_array(5901);
		when "0001011100001110" => data_out <= rom_array(5902);
		when "0001011100001111" => data_out <= rom_array(5903);
		when "0001011100010000" => data_out <= rom_array(5904);
		when "0001011100010001" => data_out <= rom_array(5905);
		when "0001011100010010" => data_out <= rom_array(5906);
		when "0001011100010011" => data_out <= rom_array(5907);
		when "0001011100010100" => data_out <= rom_array(5908);
		when "0001011100010101" => data_out <= rom_array(5909);
		when "0001011100010110" => data_out <= rom_array(5910);
		when "0001011100010111" => data_out <= rom_array(5911);
		when "0001011100011000" => data_out <= rom_array(5912);
		when "0001011100011001" => data_out <= rom_array(5913);
		when "0001011100011010" => data_out <= rom_array(5914);
		when "0001011100011011" => data_out <= rom_array(5915);
		when "0001011100011100" => data_out <= rom_array(5916);
		when "0001011100011101" => data_out <= rom_array(5917);
		when "0001011100011110" => data_out <= rom_array(5918);
		when "0001011100011111" => data_out <= rom_array(5919);
		when "0001011100100000" => data_out <= rom_array(5920);
		when "0001011100100001" => data_out <= rom_array(5921);
		when "0001011100100010" => data_out <= rom_array(5922);
		when "0001011100100011" => data_out <= rom_array(5923);
		when "0001011100100100" => data_out <= rom_array(5924);
		when "0001011100100101" => data_out <= rom_array(5925);
		when "0001011100100110" => data_out <= rom_array(5926);
		when "0001011100100111" => data_out <= rom_array(5927);
		when "0001011100101000" => data_out <= rom_array(5928);
		when "0001011100101001" => data_out <= rom_array(5929);
		when "0001011100101010" => data_out <= rom_array(5930);
		when "0001011100101011" => data_out <= rom_array(5931);
		when "0001011100101100" => data_out <= rom_array(5932);
		when "0001011100101101" => data_out <= rom_array(5933);
		when "0001011100101110" => data_out <= rom_array(5934);
		when "0001011100101111" => data_out <= rom_array(5935);
		when "0001011100110000" => data_out <= rom_array(5936);
		when "0001011100110001" => data_out <= rom_array(5937);
		when "0001011100110010" => data_out <= rom_array(5938);
		when "0001011100110011" => data_out <= rom_array(5939);
		when "0001011100110100" => data_out <= rom_array(5940);
		when "0001011100110101" => data_out <= rom_array(5941);
		when "0001011100110110" => data_out <= rom_array(5942);
		when "0001011100110111" => data_out <= rom_array(5943);
		when "0001011100111000" => data_out <= rom_array(5944);
		when "0001011100111001" => data_out <= rom_array(5945);
		when "0001011100111010" => data_out <= rom_array(5946);
		when "0001011100111011" => data_out <= rom_array(5947);
		when "0001011100111100" => data_out <= rom_array(5948);
		when "0001011100111101" => data_out <= rom_array(5949);
		when "0001011100111110" => data_out <= rom_array(5950);
		when "0001011100111111" => data_out <= rom_array(5951);
		when "0001011101000000" => data_out <= rom_array(5952);
		when "0001011101000001" => data_out <= rom_array(5953);
		when "0001011101000010" => data_out <= rom_array(5954);
		when "0001011101000011" => data_out <= rom_array(5955);
		when "0001011101000100" => data_out <= rom_array(5956);
		when "0001011101000101" => data_out <= rom_array(5957);
		when "0001011101000110" => data_out <= rom_array(5958);
		when "0001011101000111" => data_out <= rom_array(5959);
		when "0001011101001000" => data_out <= rom_array(5960);
		when "0001011101001001" => data_out <= rom_array(5961);
		when "0001011101001010" => data_out <= rom_array(5962);
		when "0001011101001011" => data_out <= rom_array(5963);
		when "0001011101001100" => data_out <= rom_array(5964);
		when "0001011101001101" => data_out <= rom_array(5965);
		when "0001011101001110" => data_out <= rom_array(5966);
		when "0001011101001111" => data_out <= rom_array(5967);
		when "0001011101010000" => data_out <= rom_array(5968);
		when "0001011101010001" => data_out <= rom_array(5969);
		when "0001011101010010" => data_out <= rom_array(5970);
		when "0001011101010011" => data_out <= rom_array(5971);
		when "0001011101010100" => data_out <= rom_array(5972);
		when "0001011101010101" => data_out <= rom_array(5973);
		when "0001011101010110" => data_out <= rom_array(5974);
		when "0001011101010111" => data_out <= rom_array(5975);
		when "0001011101011000" => data_out <= rom_array(5976);
		when "0001011101011001" => data_out <= rom_array(5977);
		when "0001011101011010" => data_out <= rom_array(5978);
		when "0001011101011011" => data_out <= rom_array(5979);
		when "0001011101011100" => data_out <= rom_array(5980);
		when "0001011101011101" => data_out <= rom_array(5981);
		when "0001011101011110" => data_out <= rom_array(5982);
		when "0001011101011111" => data_out <= rom_array(5983);
		when "0001011101100000" => data_out <= rom_array(5984);
		when "0001011101100001" => data_out <= rom_array(5985);
		when "0001011101100010" => data_out <= rom_array(5986);
		when "0001011101100011" => data_out <= rom_array(5987);
		when "0001011101100100" => data_out <= rom_array(5988);
		when "0001011101100101" => data_out <= rom_array(5989);
		when "0001011101100110" => data_out <= rom_array(5990);
		when "0001011101100111" => data_out <= rom_array(5991);
		when "0001011101101000" => data_out <= rom_array(5992);
		when "0001011101101001" => data_out <= rom_array(5993);
		when "0001011101101010" => data_out <= rom_array(5994);
		when "0001011101101011" => data_out <= rom_array(5995);
		when "0001011101101100" => data_out <= rom_array(5996);
		when "0001011101101101" => data_out <= rom_array(5997);
		when "0001011101101110" => data_out <= rom_array(5998);
		when "0001011101101111" => data_out <= rom_array(5999);
		when "0001011101110000" => data_out <= rom_array(6000);
		when "0001011101110001" => data_out <= rom_array(6001);
		when "0001011101110010" => data_out <= rom_array(6002);
		when "0001011101110011" => data_out <= rom_array(6003);
		when "0001011101110100" => data_out <= rom_array(6004);
		when "0001011101110101" => data_out <= rom_array(6005);
		when "0001011101110110" => data_out <= rom_array(6006);
		when "0001011101110111" => data_out <= rom_array(6007);
		when "0001011101111000" => data_out <= rom_array(6008);
		when "0001011101111001" => data_out <= rom_array(6009);
		when "0001011101111010" => data_out <= rom_array(6010);
		when "0001011101111011" => data_out <= rom_array(6011);
		when "0001011101111100" => data_out <= rom_array(6012);
		when "0001011101111101" => data_out <= rom_array(6013);
		when "0001011101111110" => data_out <= rom_array(6014);
		when "0001011101111111" => data_out <= rom_array(6015);
		when "0001011110000000" => data_out <= rom_array(6016);
		when "0001011110000001" => data_out <= rom_array(6017);
		when "0001011110000010" => data_out <= rom_array(6018);
		when "0001011110000011" => data_out <= rom_array(6019);
		when "0001011110000100" => data_out <= rom_array(6020);
		when "0001011110000101" => data_out <= rom_array(6021);
		when "0001011110000110" => data_out <= rom_array(6022);
		when "0001011110000111" => data_out <= rom_array(6023);
		when "0001011110001000" => data_out <= rom_array(6024);
		when "0001011110001001" => data_out <= rom_array(6025);
		when "0001011110001010" => data_out <= rom_array(6026);
		when "0001011110001011" => data_out <= rom_array(6027);
		when "0001011110001100" => data_out <= rom_array(6028);
		when "0001011110001101" => data_out <= rom_array(6029);
		when "0001011110001110" => data_out <= rom_array(6030);
		when "0001011110001111" => data_out <= rom_array(6031);
		when "0001011110010000" => data_out <= rom_array(6032);
		when "0001011110010001" => data_out <= rom_array(6033);
		when "0001011110010010" => data_out <= rom_array(6034);
		when "0001011110010011" => data_out <= rom_array(6035);
		when "0001011110010100" => data_out <= rom_array(6036);
		when "0001011110010101" => data_out <= rom_array(6037);
		when "0001011110010110" => data_out <= rom_array(6038);
		when "0001011110010111" => data_out <= rom_array(6039);
		when "0001011110011000" => data_out <= rom_array(6040);
		when "0001011110011001" => data_out <= rom_array(6041);
		when "0001011110011010" => data_out <= rom_array(6042);
		when "0001011110011011" => data_out <= rom_array(6043);
		when "0001011110011100" => data_out <= rom_array(6044);
		when "0001011110011101" => data_out <= rom_array(6045);
		when "0001011110011110" => data_out <= rom_array(6046);
		when "0001011110011111" => data_out <= rom_array(6047);
		when "0001011110100000" => data_out <= rom_array(6048);
		when "0001011110100001" => data_out <= rom_array(6049);
		when "0001011110100010" => data_out <= rom_array(6050);
		when "0001011110100011" => data_out <= rom_array(6051);
		when "0001011110100100" => data_out <= rom_array(6052);
		when "0001011110100101" => data_out <= rom_array(6053);
		when "0001011110100110" => data_out <= rom_array(6054);
		when "0001011110100111" => data_out <= rom_array(6055);
		when "0001011110101000" => data_out <= rom_array(6056);
		when "0001011110101001" => data_out <= rom_array(6057);
		when "0001011110101010" => data_out <= rom_array(6058);
		when "0001011110101011" => data_out <= rom_array(6059);
		when "0001011110101100" => data_out <= rom_array(6060);
		when "0001011110101101" => data_out <= rom_array(6061);
		when "0001011110101110" => data_out <= rom_array(6062);
		when "0001011110101111" => data_out <= rom_array(6063);
		when "0001011110110000" => data_out <= rom_array(6064);
		when "0001011110110001" => data_out <= rom_array(6065);
		when "0001011110110010" => data_out <= rom_array(6066);
		when "0001011110110011" => data_out <= rom_array(6067);
		when "0001011110110100" => data_out <= rom_array(6068);
		when "0001011110110101" => data_out <= rom_array(6069);
		when "0001011110110110" => data_out <= rom_array(6070);
		when "0001011110110111" => data_out <= rom_array(6071);
		when "0001011110111000" => data_out <= rom_array(6072);
		when "0001011110111001" => data_out <= rom_array(6073);
		when "0001011110111010" => data_out <= rom_array(6074);
		when "0001011110111011" => data_out <= rom_array(6075);
		when "0001011110111100" => data_out <= rom_array(6076);
		when "0001011110111101" => data_out <= rom_array(6077);
		when "0001011110111110" => data_out <= rom_array(6078);
		when "0001011110111111" => data_out <= rom_array(6079);
		when "0001011111000000" => data_out <= rom_array(6080);
		when "0001011111000001" => data_out <= rom_array(6081);
		when "0001011111000010" => data_out <= rom_array(6082);
		when "0001011111000011" => data_out <= rom_array(6083);
		when "0001011111000100" => data_out <= rom_array(6084);
		when "0001011111000101" => data_out <= rom_array(6085);
		when "0001011111000110" => data_out <= rom_array(6086);
		when "0001011111000111" => data_out <= rom_array(6087);
		when "0001011111001000" => data_out <= rom_array(6088);
		when "0001011111001001" => data_out <= rom_array(6089);
		when "0001011111001010" => data_out <= rom_array(6090);
		when "0001011111001011" => data_out <= rom_array(6091);
		when "0001011111001100" => data_out <= rom_array(6092);
		when "0001011111001101" => data_out <= rom_array(6093);
		when "0001011111001110" => data_out <= rom_array(6094);
		when "0001011111001111" => data_out <= rom_array(6095);
		when "0001011111010000" => data_out <= rom_array(6096);
		when "0001011111010001" => data_out <= rom_array(6097);
		when "0001011111010010" => data_out <= rom_array(6098);
		when "0001011111010011" => data_out <= rom_array(6099);
		when "0001011111010100" => data_out <= rom_array(6100);
		when "0001011111010101" => data_out <= rom_array(6101);
		when "0001011111010110" => data_out <= rom_array(6102);
		when "0001011111010111" => data_out <= rom_array(6103);
		when "0001011111011000" => data_out <= rom_array(6104);
		when "0001011111011001" => data_out <= rom_array(6105);
		when "0001011111011010" => data_out <= rom_array(6106);
		when "0001011111011011" => data_out <= rom_array(6107);
		when "0001011111011100" => data_out <= rom_array(6108);
		when "0001011111011101" => data_out <= rom_array(6109);
		when "0001011111011110" => data_out <= rom_array(6110);
		when "0001011111011111" => data_out <= rom_array(6111);
		when "0001011111100000" => data_out <= rom_array(6112);
		when "0001011111100001" => data_out <= rom_array(6113);
		when "0001011111100010" => data_out <= rom_array(6114);
		when "0001011111100011" => data_out <= rom_array(6115);
		when "0001011111100100" => data_out <= rom_array(6116);
		when "0001011111100101" => data_out <= rom_array(6117);
		when "0001011111100110" => data_out <= rom_array(6118);
		when "0001011111100111" => data_out <= rom_array(6119);
		when "0001011111101000" => data_out <= rom_array(6120);
		when "0001011111101001" => data_out <= rom_array(6121);
		when "0001011111101010" => data_out <= rom_array(6122);
		when "0001011111101011" => data_out <= rom_array(6123);
		when "0001011111101100" => data_out <= rom_array(6124);
		when "0001011111101101" => data_out <= rom_array(6125);
		when "0001011111101110" => data_out <= rom_array(6126);
		when "0001011111101111" => data_out <= rom_array(6127);
		when "0001011111110000" => data_out <= rom_array(6128);
		when "0001011111110001" => data_out <= rom_array(6129);
		when "0001011111110010" => data_out <= rom_array(6130);
		when "0001011111110011" => data_out <= rom_array(6131);
		when "0001011111110100" => data_out <= rom_array(6132);
		when "0001011111110101" => data_out <= rom_array(6133);
		when "0001011111110110" => data_out <= rom_array(6134);
		when "0001011111110111" => data_out <= rom_array(6135);
		when "0001011111111000" => data_out <= rom_array(6136);
		when "0001011111111001" => data_out <= rom_array(6137);
		when "0001011111111010" => data_out <= rom_array(6138);
		when "0001011111111011" => data_out <= rom_array(6139);
		when "0001011111111100" => data_out <= rom_array(6140);
		when "0001011111111101" => data_out <= rom_array(6141);
		when "0001011111111110" => data_out <= rom_array(6142);
		when "0001011111111111" => data_out <= rom_array(6143);
		when "0001100000000000" => data_out <= rom_array(6144);
		when "0001100000000001" => data_out <= rom_array(6145);
		when "0001100000000010" => data_out <= rom_array(6146);
		when "0001100000000011" => data_out <= rom_array(6147);
		when "0001100000000100" => data_out <= rom_array(6148);
		when "0001100000000101" => data_out <= rom_array(6149);
		when "0001100000000110" => data_out <= rom_array(6150);
		when "0001100000000111" => data_out <= rom_array(6151);
		when "0001100000001000" => data_out <= rom_array(6152);
		when "0001100000001001" => data_out <= rom_array(6153);
		when "0001100000001010" => data_out <= rom_array(6154);
		when "0001100000001011" => data_out <= rom_array(6155);
		when "0001100000001100" => data_out <= rom_array(6156);
		when "0001100000001101" => data_out <= rom_array(6157);
		when "0001100000001110" => data_out <= rom_array(6158);
		when "0001100000001111" => data_out <= rom_array(6159);
		when "0001100000010000" => data_out <= rom_array(6160);
		when "0001100000010001" => data_out <= rom_array(6161);
		when "0001100000010010" => data_out <= rom_array(6162);
		when "0001100000010011" => data_out <= rom_array(6163);
		when "0001100000010100" => data_out <= rom_array(6164);
		when "0001100000010101" => data_out <= rom_array(6165);
		when "0001100000010110" => data_out <= rom_array(6166);
		when "0001100000010111" => data_out <= rom_array(6167);
		when "0001100000011000" => data_out <= rom_array(6168);
		when "0001100000011001" => data_out <= rom_array(6169);
		when "0001100000011010" => data_out <= rom_array(6170);
		when "0001100000011011" => data_out <= rom_array(6171);
		when "0001100000011100" => data_out <= rom_array(6172);
		when "0001100000011101" => data_out <= rom_array(6173);
		when "0001100000011110" => data_out <= rom_array(6174);
		when "0001100000011111" => data_out <= rom_array(6175);
		when "0001100000100000" => data_out <= rom_array(6176);
		when "0001100000100001" => data_out <= rom_array(6177);
		when "0001100000100010" => data_out <= rom_array(6178);
		when "0001100000100011" => data_out <= rom_array(6179);
		when "0001100000100100" => data_out <= rom_array(6180);
		when "0001100000100101" => data_out <= rom_array(6181);
		when "0001100000100110" => data_out <= rom_array(6182);
		when "0001100000100111" => data_out <= rom_array(6183);
		when "0001100000101000" => data_out <= rom_array(6184);
		when "0001100000101001" => data_out <= rom_array(6185);
		when "0001100000101010" => data_out <= rom_array(6186);
		when "0001100000101011" => data_out <= rom_array(6187);
		when "0001100000101100" => data_out <= rom_array(6188);
		when "0001100000101101" => data_out <= rom_array(6189);
		when "0001100000101110" => data_out <= rom_array(6190);
		when "0001100000101111" => data_out <= rom_array(6191);
		when "0001100000110000" => data_out <= rom_array(6192);
		when "0001100000110001" => data_out <= rom_array(6193);
		when "0001100000110010" => data_out <= rom_array(6194);
		when "0001100000110011" => data_out <= rom_array(6195);
		when "0001100000110100" => data_out <= rom_array(6196);
		when "0001100000110101" => data_out <= rom_array(6197);
		when "0001100000110110" => data_out <= rom_array(6198);
		when "0001100000110111" => data_out <= rom_array(6199);
		when "0001100000111000" => data_out <= rom_array(6200);
		when "0001100000111001" => data_out <= rom_array(6201);
		when "0001100000111010" => data_out <= rom_array(6202);
		when "0001100000111011" => data_out <= rom_array(6203);
		when "0001100000111100" => data_out <= rom_array(6204);
		when "0001100000111101" => data_out <= rom_array(6205);
		when "0001100000111110" => data_out <= rom_array(6206);
		when "0001100000111111" => data_out <= rom_array(6207);
		when "0001100001000000" => data_out <= rom_array(6208);
		when "0001100001000001" => data_out <= rom_array(6209);
		when "0001100001000010" => data_out <= rom_array(6210);
		when "0001100001000011" => data_out <= rom_array(6211);
		when "0001100001000100" => data_out <= rom_array(6212);
		when "0001100001000101" => data_out <= rom_array(6213);
		when "0001100001000110" => data_out <= rom_array(6214);
		when "0001100001000111" => data_out <= rom_array(6215);
		when "0001100001001000" => data_out <= rom_array(6216);
		when "0001100001001001" => data_out <= rom_array(6217);
		when "0001100001001010" => data_out <= rom_array(6218);
		when "0001100001001011" => data_out <= rom_array(6219);
		when "0001100001001100" => data_out <= rom_array(6220);
		when "0001100001001101" => data_out <= rom_array(6221);
		when "0001100001001110" => data_out <= rom_array(6222);
		when "0001100001001111" => data_out <= rom_array(6223);
		when "0001100001010000" => data_out <= rom_array(6224);
		when "0001100001010001" => data_out <= rom_array(6225);
		when "0001100001010010" => data_out <= rom_array(6226);
		when "0001100001010011" => data_out <= rom_array(6227);
		when "0001100001010100" => data_out <= rom_array(6228);
		when "0001100001010101" => data_out <= rom_array(6229);
		when "0001100001010110" => data_out <= rom_array(6230);
		when "0001100001010111" => data_out <= rom_array(6231);
		when "0001100001011000" => data_out <= rom_array(6232);
		when "0001100001011001" => data_out <= rom_array(6233);
		when "0001100001011010" => data_out <= rom_array(6234);
		when "0001100001011011" => data_out <= rom_array(6235);
		when "0001100001011100" => data_out <= rom_array(6236);
		when "0001100001011101" => data_out <= rom_array(6237);
		when "0001100001011110" => data_out <= rom_array(6238);
		when "0001100001011111" => data_out <= rom_array(6239);
		when "0001100001100000" => data_out <= rom_array(6240);
		when "0001100001100001" => data_out <= rom_array(6241);
		when "0001100001100010" => data_out <= rom_array(6242);
		when "0001100001100011" => data_out <= rom_array(6243);
		when "0001100001100100" => data_out <= rom_array(6244);
		when "0001100001100101" => data_out <= rom_array(6245);
		when "0001100001100110" => data_out <= rom_array(6246);
		when "0001100001100111" => data_out <= rom_array(6247);
		when "0001100001101000" => data_out <= rom_array(6248);
		when "0001100001101001" => data_out <= rom_array(6249);
		when "0001100001101010" => data_out <= rom_array(6250);
		when "0001100001101011" => data_out <= rom_array(6251);
		when "0001100001101100" => data_out <= rom_array(6252);
		when "0001100001101101" => data_out <= rom_array(6253);
		when "0001100001101110" => data_out <= rom_array(6254);
		when "0001100001101111" => data_out <= rom_array(6255);
		when "0001100001110000" => data_out <= rom_array(6256);
		when "0001100001110001" => data_out <= rom_array(6257);
		when "0001100001110010" => data_out <= rom_array(6258);
		when "0001100001110011" => data_out <= rom_array(6259);
		when "0001100001110100" => data_out <= rom_array(6260);
		when "0001100001110101" => data_out <= rom_array(6261);
		when "0001100001110110" => data_out <= rom_array(6262);
		when "0001100001110111" => data_out <= rom_array(6263);
		when "0001100001111000" => data_out <= rom_array(6264);
		when "0001100001111001" => data_out <= rom_array(6265);
		when "0001100001111010" => data_out <= rom_array(6266);
		when "0001100001111011" => data_out <= rom_array(6267);
		when "0001100001111100" => data_out <= rom_array(6268);
		when "0001100001111101" => data_out <= rom_array(6269);
		when "0001100001111110" => data_out <= rom_array(6270);
		when "0001100001111111" => data_out <= rom_array(6271);
		when "0001100010000000" => data_out <= rom_array(6272);
		when "0001100010000001" => data_out <= rom_array(6273);
		when "0001100010000010" => data_out <= rom_array(6274);
		when "0001100010000011" => data_out <= rom_array(6275);
		when "0001100010000100" => data_out <= rom_array(6276);
		when "0001100010000101" => data_out <= rom_array(6277);
		when "0001100010000110" => data_out <= rom_array(6278);
		when "0001100010000111" => data_out <= rom_array(6279);
		when "0001100010001000" => data_out <= rom_array(6280);
		when "0001100010001001" => data_out <= rom_array(6281);
		when "0001100010001010" => data_out <= rom_array(6282);
		when "0001100010001011" => data_out <= rom_array(6283);
		when "0001100010001100" => data_out <= rom_array(6284);
		when "0001100010001101" => data_out <= rom_array(6285);
		when "0001100010001110" => data_out <= rom_array(6286);
		when "0001100010001111" => data_out <= rom_array(6287);
		when "0001100010010000" => data_out <= rom_array(6288);
		when "0001100010010001" => data_out <= rom_array(6289);
		when "0001100010010010" => data_out <= rom_array(6290);
		when "0001100010010011" => data_out <= rom_array(6291);
		when "0001100010010100" => data_out <= rom_array(6292);
		when "0001100010010101" => data_out <= rom_array(6293);
		when "0001100010010110" => data_out <= rom_array(6294);
		when "0001100010010111" => data_out <= rom_array(6295);
		when "0001100010011000" => data_out <= rom_array(6296);
		when "0001100010011001" => data_out <= rom_array(6297);
		when "0001100010011010" => data_out <= rom_array(6298);
		when "0001100010011011" => data_out <= rom_array(6299);
		when "0001100010011100" => data_out <= rom_array(6300);
		when "0001100010011101" => data_out <= rom_array(6301);
		when "0001100010011110" => data_out <= rom_array(6302);
		when "0001100010011111" => data_out <= rom_array(6303);
		when "0001100010100000" => data_out <= rom_array(6304);
		when "0001100010100001" => data_out <= rom_array(6305);
		when "0001100010100010" => data_out <= rom_array(6306);
		when "0001100010100011" => data_out <= rom_array(6307);
		when "0001100010100100" => data_out <= rom_array(6308);
		when "0001100010100101" => data_out <= rom_array(6309);
		when "0001100010100110" => data_out <= rom_array(6310);
		when "0001100010100111" => data_out <= rom_array(6311);
		when "0001100010101000" => data_out <= rom_array(6312);
		when "0001100010101001" => data_out <= rom_array(6313);
		when "0001100010101010" => data_out <= rom_array(6314);
		when "0001100010101011" => data_out <= rom_array(6315);
		when "0001100010101100" => data_out <= rom_array(6316);
		when "0001100010101101" => data_out <= rom_array(6317);
		when "0001100010101110" => data_out <= rom_array(6318);
		when "0001100010101111" => data_out <= rom_array(6319);
		when "0001100010110000" => data_out <= rom_array(6320);
		when "0001100010110001" => data_out <= rom_array(6321);
		when "0001100010110010" => data_out <= rom_array(6322);
		when "0001100010110011" => data_out <= rom_array(6323);
		when "0001100010110100" => data_out <= rom_array(6324);
		when "0001100010110101" => data_out <= rom_array(6325);
		when "0001100010110110" => data_out <= rom_array(6326);
		when "0001100010110111" => data_out <= rom_array(6327);
		when "0001100010111000" => data_out <= rom_array(6328);
		when "0001100010111001" => data_out <= rom_array(6329);
		when "0001100010111010" => data_out <= rom_array(6330);
		when "0001100010111011" => data_out <= rom_array(6331);
		when "0001100010111100" => data_out <= rom_array(6332);
		when "0001100010111101" => data_out <= rom_array(6333);
		when "0001100010111110" => data_out <= rom_array(6334);
		when "0001100010111111" => data_out <= rom_array(6335);
		when "0001100011000000" => data_out <= rom_array(6336);
		when "0001100011000001" => data_out <= rom_array(6337);
		when "0001100011000010" => data_out <= rom_array(6338);
		when "0001100011000011" => data_out <= rom_array(6339);
		when "0001100011000100" => data_out <= rom_array(6340);
		when "0001100011000101" => data_out <= rom_array(6341);
		when "0001100011000110" => data_out <= rom_array(6342);
		when "0001100011000111" => data_out <= rom_array(6343);
		when "0001100011001000" => data_out <= rom_array(6344);
		when "0001100011001001" => data_out <= rom_array(6345);
		when "0001100011001010" => data_out <= rom_array(6346);
		when "0001100011001011" => data_out <= rom_array(6347);
		when "0001100011001100" => data_out <= rom_array(6348);
		when "0001100011001101" => data_out <= rom_array(6349);
		when "0001100011001110" => data_out <= rom_array(6350);
		when "0001100011001111" => data_out <= rom_array(6351);
		when "0001100011010000" => data_out <= rom_array(6352);
		when "0001100011010001" => data_out <= rom_array(6353);
		when "0001100011010010" => data_out <= rom_array(6354);
		when "0001100011010011" => data_out <= rom_array(6355);
		when "0001100011010100" => data_out <= rom_array(6356);
		when "0001100011010101" => data_out <= rom_array(6357);
		when "0001100011010110" => data_out <= rom_array(6358);
		when "0001100011010111" => data_out <= rom_array(6359);
		when "0001100011011000" => data_out <= rom_array(6360);
		when "0001100011011001" => data_out <= rom_array(6361);
		when "0001100011011010" => data_out <= rom_array(6362);
		when "0001100011011011" => data_out <= rom_array(6363);
		when "0001100011011100" => data_out <= rom_array(6364);
		when "0001100011011101" => data_out <= rom_array(6365);
		when "0001100011011110" => data_out <= rom_array(6366);
		when "0001100011011111" => data_out <= rom_array(6367);
		when "0001100011100000" => data_out <= rom_array(6368);
		when "0001100011100001" => data_out <= rom_array(6369);
		when "0001100011100010" => data_out <= rom_array(6370);
		when "0001100011100011" => data_out <= rom_array(6371);
		when "0001100011100100" => data_out <= rom_array(6372);
		when "0001100011100101" => data_out <= rom_array(6373);
		when "0001100011100110" => data_out <= rom_array(6374);
		when "0001100011100111" => data_out <= rom_array(6375);
		when "0001100011101000" => data_out <= rom_array(6376);
		when "0001100011101001" => data_out <= rom_array(6377);
		when "0001100011101010" => data_out <= rom_array(6378);
		when "0001100011101011" => data_out <= rom_array(6379);
		when "0001100011101100" => data_out <= rom_array(6380);
		when "0001100011101101" => data_out <= rom_array(6381);
		when "0001100011101110" => data_out <= rom_array(6382);
		when "0001100011101111" => data_out <= rom_array(6383);
		when "0001100011110000" => data_out <= rom_array(6384);
		when "0001100011110001" => data_out <= rom_array(6385);
		when "0001100011110010" => data_out <= rom_array(6386);
		when "0001100011110011" => data_out <= rom_array(6387);
		when "0001100011110100" => data_out <= rom_array(6388);
		when "0001100011110101" => data_out <= rom_array(6389);
		when "0001100011110110" => data_out <= rom_array(6390);
		when "0001100011110111" => data_out <= rom_array(6391);
		when "0001100011111000" => data_out <= rom_array(6392);
		when "0001100011111001" => data_out <= rom_array(6393);
		when "0001100011111010" => data_out <= rom_array(6394);
		when "0001100011111011" => data_out <= rom_array(6395);
		when "0001100011111100" => data_out <= rom_array(6396);
		when "0001100011111101" => data_out <= rom_array(6397);
		when "0001100011111110" => data_out <= rom_array(6398);
		when "0001100011111111" => data_out <= rom_array(6399);
		when "0001100100000000" => data_out <= rom_array(6400);
		when "0001100100000001" => data_out <= rom_array(6401);
		when "0001100100000010" => data_out <= rom_array(6402);
		when "0001100100000011" => data_out <= rom_array(6403);
		when "0001100100000100" => data_out <= rom_array(6404);
		when "0001100100000101" => data_out <= rom_array(6405);
		when "0001100100000110" => data_out <= rom_array(6406);
		when "0001100100000111" => data_out <= rom_array(6407);
		when "0001100100001000" => data_out <= rom_array(6408);
		when "0001100100001001" => data_out <= rom_array(6409);
		when "0001100100001010" => data_out <= rom_array(6410);
		when "0001100100001011" => data_out <= rom_array(6411);
		when "0001100100001100" => data_out <= rom_array(6412);
		when "0001100100001101" => data_out <= rom_array(6413);
		when "0001100100001110" => data_out <= rom_array(6414);
		when "0001100100001111" => data_out <= rom_array(6415);
		when "0001100100010000" => data_out <= rom_array(6416);
		when "0001100100010001" => data_out <= rom_array(6417);
		when "0001100100010010" => data_out <= rom_array(6418);
		when "0001100100010011" => data_out <= rom_array(6419);
		when "0001100100010100" => data_out <= rom_array(6420);
		when "0001100100010101" => data_out <= rom_array(6421);
		when "0001100100010110" => data_out <= rom_array(6422);
		when "0001100100010111" => data_out <= rom_array(6423);
		when "0001100100011000" => data_out <= rom_array(6424);
		when "0001100100011001" => data_out <= rom_array(6425);
		when "0001100100011010" => data_out <= rom_array(6426);
		when "0001100100011011" => data_out <= rom_array(6427);
		when "0001100100011100" => data_out <= rom_array(6428);
		when "0001100100011101" => data_out <= rom_array(6429);
		when "0001100100011110" => data_out <= rom_array(6430);
		when "0001100100011111" => data_out <= rom_array(6431);
		when "0001100100100000" => data_out <= rom_array(6432);
		when "0001100100100001" => data_out <= rom_array(6433);
		when "0001100100100010" => data_out <= rom_array(6434);
		when "0001100100100011" => data_out <= rom_array(6435);
		when "0001100100100100" => data_out <= rom_array(6436);
		when "0001100100100101" => data_out <= rom_array(6437);
		when "0001100100100110" => data_out <= rom_array(6438);
		when "0001100100100111" => data_out <= rom_array(6439);
		when "0001100100101000" => data_out <= rom_array(6440);
		when "0001100100101001" => data_out <= rom_array(6441);
		when "0001100100101010" => data_out <= rom_array(6442);
		when "0001100100101011" => data_out <= rom_array(6443);
		when "0001100100101100" => data_out <= rom_array(6444);
		when "0001100100101101" => data_out <= rom_array(6445);
		when "0001100100101110" => data_out <= rom_array(6446);
		when "0001100100101111" => data_out <= rom_array(6447);
		when "0001100100110000" => data_out <= rom_array(6448);
		when "0001100100110001" => data_out <= rom_array(6449);
		when "0001100100110010" => data_out <= rom_array(6450);
		when "0001100100110011" => data_out <= rom_array(6451);
		when "0001100100110100" => data_out <= rom_array(6452);
		when "0001100100110101" => data_out <= rom_array(6453);
		when "0001100100110110" => data_out <= rom_array(6454);
		when "0001100100110111" => data_out <= rom_array(6455);
		when "0001100100111000" => data_out <= rom_array(6456);
		when "0001100100111001" => data_out <= rom_array(6457);
		when "0001100100111010" => data_out <= rom_array(6458);
		when "0001100100111011" => data_out <= rom_array(6459);
		when "0001100100111100" => data_out <= rom_array(6460);
		when "0001100100111101" => data_out <= rom_array(6461);
		when "0001100100111110" => data_out <= rom_array(6462);
		when "0001100100111111" => data_out <= rom_array(6463);
		when "0001100101000000" => data_out <= rom_array(6464);
		when "0001100101000001" => data_out <= rom_array(6465);
		when "0001100101000010" => data_out <= rom_array(6466);
		when "0001100101000011" => data_out <= rom_array(6467);
		when "0001100101000100" => data_out <= rom_array(6468);
		when "0001100101000101" => data_out <= rom_array(6469);
		when "0001100101000110" => data_out <= rom_array(6470);
		when "0001100101000111" => data_out <= rom_array(6471);
		when "0001100101001000" => data_out <= rom_array(6472);
		when "0001100101001001" => data_out <= rom_array(6473);
		when "0001100101001010" => data_out <= rom_array(6474);
		when "0001100101001011" => data_out <= rom_array(6475);
		when "0001100101001100" => data_out <= rom_array(6476);
		when "0001100101001101" => data_out <= rom_array(6477);
		when "0001100101001110" => data_out <= rom_array(6478);
		when "0001100101001111" => data_out <= rom_array(6479);
		when "0001100101010000" => data_out <= rom_array(6480);
		when "0001100101010001" => data_out <= rom_array(6481);
		when "0001100101010010" => data_out <= rom_array(6482);
		when "0001100101010011" => data_out <= rom_array(6483);
		when "0001100101010100" => data_out <= rom_array(6484);
		when "0001100101010101" => data_out <= rom_array(6485);
		when "0001100101010110" => data_out <= rom_array(6486);
		when "0001100101010111" => data_out <= rom_array(6487);
		when "0001100101011000" => data_out <= rom_array(6488);
		when "0001100101011001" => data_out <= rom_array(6489);
		when "0001100101011010" => data_out <= rom_array(6490);
		when "0001100101011011" => data_out <= rom_array(6491);
		when "0001100101011100" => data_out <= rom_array(6492);
		when "0001100101011101" => data_out <= rom_array(6493);
		when "0001100101011110" => data_out <= rom_array(6494);
		when "0001100101011111" => data_out <= rom_array(6495);
		when "0001100101100000" => data_out <= rom_array(6496);
		when "0001100101100001" => data_out <= rom_array(6497);
		when "0001100101100010" => data_out <= rom_array(6498);
		when "0001100101100011" => data_out <= rom_array(6499);
		when "0001100101100100" => data_out <= rom_array(6500);
		when "0001100101100101" => data_out <= rom_array(6501);
		when "0001100101100110" => data_out <= rom_array(6502);
		when "0001100101100111" => data_out <= rom_array(6503);
		when "0001100101101000" => data_out <= rom_array(6504);
		when "0001100101101001" => data_out <= rom_array(6505);
		when "0001100101101010" => data_out <= rom_array(6506);
		when "0001100101101011" => data_out <= rom_array(6507);
		when "0001100101101100" => data_out <= rom_array(6508);
		when "0001100101101101" => data_out <= rom_array(6509);
		when "0001100101101110" => data_out <= rom_array(6510);
		when "0001100101101111" => data_out <= rom_array(6511);
		when "0001100101110000" => data_out <= rom_array(6512);
		when "0001100101110001" => data_out <= rom_array(6513);
		when "0001100101110010" => data_out <= rom_array(6514);
		when "0001100101110011" => data_out <= rom_array(6515);
		when "0001100101110100" => data_out <= rom_array(6516);
		when "0001100101110101" => data_out <= rom_array(6517);
		when "0001100101110110" => data_out <= rom_array(6518);
		when "0001100101110111" => data_out <= rom_array(6519);
		when "0001100101111000" => data_out <= rom_array(6520);
		when "0001100101111001" => data_out <= rom_array(6521);
		when "0001100101111010" => data_out <= rom_array(6522);
		when "0001100101111011" => data_out <= rom_array(6523);
		when "0001100101111100" => data_out <= rom_array(6524);
		when "0001100101111101" => data_out <= rom_array(6525);
		when "0001100101111110" => data_out <= rom_array(6526);
		when "0001100101111111" => data_out <= rom_array(6527);
		when "0001100110000000" => data_out <= rom_array(6528);
		when "0001100110000001" => data_out <= rom_array(6529);
		when "0001100110000010" => data_out <= rom_array(6530);
		when "0001100110000011" => data_out <= rom_array(6531);
		when "0001100110000100" => data_out <= rom_array(6532);
		when "0001100110000101" => data_out <= rom_array(6533);
		when "0001100110000110" => data_out <= rom_array(6534);
		when "0001100110000111" => data_out <= rom_array(6535);
		when "0001100110001000" => data_out <= rom_array(6536);
		when "0001100110001001" => data_out <= rom_array(6537);
		when "0001100110001010" => data_out <= rom_array(6538);
		when "0001100110001011" => data_out <= rom_array(6539);
		when "0001100110001100" => data_out <= rom_array(6540);
		when "0001100110001101" => data_out <= rom_array(6541);
		when "0001100110001110" => data_out <= rom_array(6542);
		when "0001100110001111" => data_out <= rom_array(6543);
		when "0001100110010000" => data_out <= rom_array(6544);
		when "0001100110010001" => data_out <= rom_array(6545);
		when "0001100110010010" => data_out <= rom_array(6546);
		when "0001100110010011" => data_out <= rom_array(6547);
		when "0001100110010100" => data_out <= rom_array(6548);
		when "0001100110010101" => data_out <= rom_array(6549);
		when "0001100110010110" => data_out <= rom_array(6550);
		when "0001100110010111" => data_out <= rom_array(6551);
		when "0001100110011000" => data_out <= rom_array(6552);
		when "0001100110011001" => data_out <= rom_array(6553);
		when "0001100110011010" => data_out <= rom_array(6554);
		when "0001100110011011" => data_out <= rom_array(6555);
		when "0001100110011100" => data_out <= rom_array(6556);
		when "0001100110011101" => data_out <= rom_array(6557);
		when "0001100110011110" => data_out <= rom_array(6558);
		when "0001100110011111" => data_out <= rom_array(6559);
		when "0001100110100000" => data_out <= rom_array(6560);
		when "0001100110100001" => data_out <= rom_array(6561);
		when "0001100110100010" => data_out <= rom_array(6562);
		when "0001100110100011" => data_out <= rom_array(6563);
		when "0001100110100100" => data_out <= rom_array(6564);
		when "0001100110100101" => data_out <= rom_array(6565);
		when "0001100110100110" => data_out <= rom_array(6566);
		when "0001100110100111" => data_out <= rom_array(6567);
		when "0001100110101000" => data_out <= rom_array(6568);
		when "0001100110101001" => data_out <= rom_array(6569);
		when "0001100110101010" => data_out <= rom_array(6570);
		when "0001100110101011" => data_out <= rom_array(6571);
		when "0001100110101100" => data_out <= rom_array(6572);
		when "0001100110101101" => data_out <= rom_array(6573);
		when "0001100110101110" => data_out <= rom_array(6574);
		when "0001100110101111" => data_out <= rom_array(6575);
		when "0001100110110000" => data_out <= rom_array(6576);
		when "0001100110110001" => data_out <= rom_array(6577);
		when "0001100110110010" => data_out <= rom_array(6578);
		when "0001100110110011" => data_out <= rom_array(6579);
		when "0001100110110100" => data_out <= rom_array(6580);
		when "0001100110110101" => data_out <= rom_array(6581);
		when "0001100110110110" => data_out <= rom_array(6582);
		when "0001100110110111" => data_out <= rom_array(6583);
		when "0001100110111000" => data_out <= rom_array(6584);
		when "0001100110111001" => data_out <= rom_array(6585);
		when "0001100110111010" => data_out <= rom_array(6586);
		when "0001100110111011" => data_out <= rom_array(6587);
		when "0001100110111100" => data_out <= rom_array(6588);
		when "0001100110111101" => data_out <= rom_array(6589);
		when "0001100110111110" => data_out <= rom_array(6590);
		when "0001100110111111" => data_out <= rom_array(6591);
		when "0001100111000000" => data_out <= rom_array(6592);
		when "0001100111000001" => data_out <= rom_array(6593);
		when "0001100111000010" => data_out <= rom_array(6594);
		when "0001100111000011" => data_out <= rom_array(6595);
		when "0001100111000100" => data_out <= rom_array(6596);
		when "0001100111000101" => data_out <= rom_array(6597);
		when "0001100111000110" => data_out <= rom_array(6598);
		when "0001100111000111" => data_out <= rom_array(6599);
		when "0001100111001000" => data_out <= rom_array(6600);
		when "0001100111001001" => data_out <= rom_array(6601);
		when "0001100111001010" => data_out <= rom_array(6602);
		when "0001100111001011" => data_out <= rom_array(6603);
		when "0001100111001100" => data_out <= rom_array(6604);
		when "0001100111001101" => data_out <= rom_array(6605);
		when "0001100111001110" => data_out <= rom_array(6606);
		when "0001100111001111" => data_out <= rom_array(6607);
		when "0001100111010000" => data_out <= rom_array(6608);
		when "0001100111010001" => data_out <= rom_array(6609);
		when "0001100111010010" => data_out <= rom_array(6610);
		when "0001100111010011" => data_out <= rom_array(6611);
		when "0001100111010100" => data_out <= rom_array(6612);
		when "0001100111010101" => data_out <= rom_array(6613);
		when "0001100111010110" => data_out <= rom_array(6614);
		when "0001100111010111" => data_out <= rom_array(6615);
		when "0001100111011000" => data_out <= rom_array(6616);
		when "0001100111011001" => data_out <= rom_array(6617);
		when "0001100111011010" => data_out <= rom_array(6618);
		when "0001100111011011" => data_out <= rom_array(6619);
		when "0001100111011100" => data_out <= rom_array(6620);
		when "0001100111011101" => data_out <= rom_array(6621);
		when "0001100111011110" => data_out <= rom_array(6622);
		when "0001100111011111" => data_out <= rom_array(6623);
		when "0001100111100000" => data_out <= rom_array(6624);
		when "0001100111100001" => data_out <= rom_array(6625);
		when "0001100111100010" => data_out <= rom_array(6626);
		when "0001100111100011" => data_out <= rom_array(6627);
		when "0001100111100100" => data_out <= rom_array(6628);
		when "0001100111100101" => data_out <= rom_array(6629);
		when "0001100111100110" => data_out <= rom_array(6630);
		when "0001100111100111" => data_out <= rom_array(6631);
		when "0001100111101000" => data_out <= rom_array(6632);
		when "0001100111101001" => data_out <= rom_array(6633);
		when "0001100111101010" => data_out <= rom_array(6634);
		when "0001100111101011" => data_out <= rom_array(6635);
		when "0001100111101100" => data_out <= rom_array(6636);
		when "0001100111101101" => data_out <= rom_array(6637);
		when "0001100111101110" => data_out <= rom_array(6638);
		when "0001100111101111" => data_out <= rom_array(6639);
		when "0001100111110000" => data_out <= rom_array(6640);
		when "0001100111110001" => data_out <= rom_array(6641);
		when "0001100111110010" => data_out <= rom_array(6642);
		when "0001100111110011" => data_out <= rom_array(6643);
		when "0001100111110100" => data_out <= rom_array(6644);
		when "0001100111110101" => data_out <= rom_array(6645);
		when "0001100111110110" => data_out <= rom_array(6646);
		when "0001100111110111" => data_out <= rom_array(6647);
		when "0001100111111000" => data_out <= rom_array(6648);
		when "0001100111111001" => data_out <= rom_array(6649);
		when "0001100111111010" => data_out <= rom_array(6650);
		when "0001100111111011" => data_out <= rom_array(6651);
		when "0001100111111100" => data_out <= rom_array(6652);
		when "0001100111111101" => data_out <= rom_array(6653);
		when "0001100111111110" => data_out <= rom_array(6654);
		when "0001100111111111" => data_out <= rom_array(6655);
		when "0001101000000000" => data_out <= rom_array(6656);
		when "0001101000000001" => data_out <= rom_array(6657);
		when "0001101000000010" => data_out <= rom_array(6658);
		when "0001101000000011" => data_out <= rom_array(6659);
		when "0001101000000100" => data_out <= rom_array(6660);
		when "0001101000000101" => data_out <= rom_array(6661);
		when "0001101000000110" => data_out <= rom_array(6662);
		when "0001101000000111" => data_out <= rom_array(6663);
		when "0001101000001000" => data_out <= rom_array(6664);
		when "0001101000001001" => data_out <= rom_array(6665);
		when "0001101000001010" => data_out <= rom_array(6666);
		when "0001101000001011" => data_out <= rom_array(6667);
		when "0001101000001100" => data_out <= rom_array(6668);
		when "0001101000001101" => data_out <= rom_array(6669);
		when "0001101000001110" => data_out <= rom_array(6670);
		when "0001101000001111" => data_out <= rom_array(6671);
		when "0001101000010000" => data_out <= rom_array(6672);
		when "0001101000010001" => data_out <= rom_array(6673);
		when "0001101000010010" => data_out <= rom_array(6674);
		when "0001101000010011" => data_out <= rom_array(6675);
		when "0001101000010100" => data_out <= rom_array(6676);
		when "0001101000010101" => data_out <= rom_array(6677);
		when "0001101000010110" => data_out <= rom_array(6678);
		when "0001101000010111" => data_out <= rom_array(6679);
		when "0001101000011000" => data_out <= rom_array(6680);
		when "0001101000011001" => data_out <= rom_array(6681);
		when "0001101000011010" => data_out <= rom_array(6682);
		when "0001101000011011" => data_out <= rom_array(6683);
		when "0001101000011100" => data_out <= rom_array(6684);
		when "0001101000011101" => data_out <= rom_array(6685);
		when "0001101000011110" => data_out <= rom_array(6686);
		when "0001101000011111" => data_out <= rom_array(6687);
		when "0001101000100000" => data_out <= rom_array(6688);
		when "0001101000100001" => data_out <= rom_array(6689);
		when "0001101000100010" => data_out <= rom_array(6690);
		when "0001101000100011" => data_out <= rom_array(6691);
		when "0001101000100100" => data_out <= rom_array(6692);
		when "0001101000100101" => data_out <= rom_array(6693);
		when "0001101000100110" => data_out <= rom_array(6694);
		when "0001101000100111" => data_out <= rom_array(6695);
		when "0001101000101000" => data_out <= rom_array(6696);
		when "0001101000101001" => data_out <= rom_array(6697);
		when "0001101000101010" => data_out <= rom_array(6698);
		when "0001101000101011" => data_out <= rom_array(6699);
		when "0001101000101100" => data_out <= rom_array(6700);
		when "0001101000101101" => data_out <= rom_array(6701);
		when "0001101000101110" => data_out <= rom_array(6702);
		when "0001101000101111" => data_out <= rom_array(6703);
		when "0001101000110000" => data_out <= rom_array(6704);
		when "0001101000110001" => data_out <= rom_array(6705);
		when "0001101000110010" => data_out <= rom_array(6706);
		when "0001101000110011" => data_out <= rom_array(6707);
		when "0001101000110100" => data_out <= rom_array(6708);
		when "0001101000110101" => data_out <= rom_array(6709);
		when "0001101000110110" => data_out <= rom_array(6710);
		when "0001101000110111" => data_out <= rom_array(6711);
		when "0001101000111000" => data_out <= rom_array(6712);
		when "0001101000111001" => data_out <= rom_array(6713);
		when "0001101000111010" => data_out <= rom_array(6714);
		when "0001101000111011" => data_out <= rom_array(6715);
		when "0001101000111100" => data_out <= rom_array(6716);
		when "0001101000111101" => data_out <= rom_array(6717);
		when "0001101000111110" => data_out <= rom_array(6718);
		when "0001101000111111" => data_out <= rom_array(6719);
		when "0001101001000000" => data_out <= rom_array(6720);
		when "0001101001000001" => data_out <= rom_array(6721);
		when "0001101001000010" => data_out <= rom_array(6722);
		when "0001101001000011" => data_out <= rom_array(6723);
		when "0001101001000100" => data_out <= rom_array(6724);
		when "0001101001000101" => data_out <= rom_array(6725);
		when "0001101001000110" => data_out <= rom_array(6726);
		when "0001101001000111" => data_out <= rom_array(6727);
		when "0001101001001000" => data_out <= rom_array(6728);
		when "0001101001001001" => data_out <= rom_array(6729);
		when "0001101001001010" => data_out <= rom_array(6730);
		when "0001101001001011" => data_out <= rom_array(6731);
		when "0001101001001100" => data_out <= rom_array(6732);
		when "0001101001001101" => data_out <= rom_array(6733);
		when "0001101001001110" => data_out <= rom_array(6734);
		when "0001101001001111" => data_out <= rom_array(6735);
		when "0001101001010000" => data_out <= rom_array(6736);
		when "0001101001010001" => data_out <= rom_array(6737);
		when "0001101001010010" => data_out <= rom_array(6738);
		when "0001101001010011" => data_out <= rom_array(6739);
		when "0001101001010100" => data_out <= rom_array(6740);
		when "0001101001010101" => data_out <= rom_array(6741);
		when "0001101001010110" => data_out <= rom_array(6742);
		when "0001101001010111" => data_out <= rom_array(6743);
		when "0001101001011000" => data_out <= rom_array(6744);
		when "0001101001011001" => data_out <= rom_array(6745);
		when "0001101001011010" => data_out <= rom_array(6746);
		when "0001101001011011" => data_out <= rom_array(6747);
		when "0001101001011100" => data_out <= rom_array(6748);
		when "0001101001011101" => data_out <= rom_array(6749);
		when "0001101001011110" => data_out <= rom_array(6750);
		when "0001101001011111" => data_out <= rom_array(6751);
		when "0001101001100000" => data_out <= rom_array(6752);
		when "0001101001100001" => data_out <= rom_array(6753);
		when "0001101001100010" => data_out <= rom_array(6754);
		when "0001101001100011" => data_out <= rom_array(6755);
		when "0001101001100100" => data_out <= rom_array(6756);
		when "0001101001100101" => data_out <= rom_array(6757);
		when "0001101001100110" => data_out <= rom_array(6758);
		when "0001101001100111" => data_out <= rom_array(6759);
		when "0001101001101000" => data_out <= rom_array(6760);
		when "0001101001101001" => data_out <= rom_array(6761);
		when "0001101001101010" => data_out <= rom_array(6762);
		when "0001101001101011" => data_out <= rom_array(6763);
		when "0001101001101100" => data_out <= rom_array(6764);
		when "0001101001101101" => data_out <= rom_array(6765);
		when "0001101001101110" => data_out <= rom_array(6766);
		when "0001101001101111" => data_out <= rom_array(6767);
		when "0001101001110000" => data_out <= rom_array(6768);
		when "0001101001110001" => data_out <= rom_array(6769);
		when "0001101001110010" => data_out <= rom_array(6770);
		when "0001101001110011" => data_out <= rom_array(6771);
		when "0001101001110100" => data_out <= rom_array(6772);
		when "0001101001110101" => data_out <= rom_array(6773);
		when "0001101001110110" => data_out <= rom_array(6774);
		when "0001101001110111" => data_out <= rom_array(6775);
		when "0001101001111000" => data_out <= rom_array(6776);
		when "0001101001111001" => data_out <= rom_array(6777);
		when "0001101001111010" => data_out <= rom_array(6778);
		when "0001101001111011" => data_out <= rom_array(6779);
		when "0001101001111100" => data_out <= rom_array(6780);
		when "0001101001111101" => data_out <= rom_array(6781);
		when "0001101001111110" => data_out <= rom_array(6782);
		when "0001101001111111" => data_out <= rom_array(6783);
		when "0001101010000000" => data_out <= rom_array(6784);
		when "0001101010000001" => data_out <= rom_array(6785);
		when "0001101010000010" => data_out <= rom_array(6786);
		when "0001101010000011" => data_out <= rom_array(6787);
		when "0001101010000100" => data_out <= rom_array(6788);
		when "0001101010000101" => data_out <= rom_array(6789);
		when "0001101010000110" => data_out <= rom_array(6790);
		when "0001101010000111" => data_out <= rom_array(6791);
		when "0001101010001000" => data_out <= rom_array(6792);
		when "0001101010001001" => data_out <= rom_array(6793);
		when "0001101010001010" => data_out <= rom_array(6794);
		when "0001101010001011" => data_out <= rom_array(6795);
		when "0001101010001100" => data_out <= rom_array(6796);
		when "0001101010001101" => data_out <= rom_array(6797);
		when "0001101010001110" => data_out <= rom_array(6798);
		when "0001101010001111" => data_out <= rom_array(6799);
		when "0001101010010000" => data_out <= rom_array(6800);
		when "0001101010010001" => data_out <= rom_array(6801);
		when "0001101010010010" => data_out <= rom_array(6802);
		when "0001101010010011" => data_out <= rom_array(6803);
		when "0001101010010100" => data_out <= rom_array(6804);
		when "0001101010010101" => data_out <= rom_array(6805);
		when "0001101010010110" => data_out <= rom_array(6806);
		when "0001101010010111" => data_out <= rom_array(6807);
		when "0001101010011000" => data_out <= rom_array(6808);
		when "0001101010011001" => data_out <= rom_array(6809);
		when "0001101010011010" => data_out <= rom_array(6810);
		when "0001101010011011" => data_out <= rom_array(6811);
		when "0001101010011100" => data_out <= rom_array(6812);
		when "0001101010011101" => data_out <= rom_array(6813);
		when "0001101010011110" => data_out <= rom_array(6814);
		when "0001101010011111" => data_out <= rom_array(6815);
		when "0001101010100000" => data_out <= rom_array(6816);
		when "0001101010100001" => data_out <= rom_array(6817);
		when "0001101010100010" => data_out <= rom_array(6818);
		when "0001101010100011" => data_out <= rom_array(6819);
		when "0001101010100100" => data_out <= rom_array(6820);
		when "0001101010100101" => data_out <= rom_array(6821);
		when "0001101010100110" => data_out <= rom_array(6822);
		when "0001101010100111" => data_out <= rom_array(6823);
		when "0001101010101000" => data_out <= rom_array(6824);
		when "0001101010101001" => data_out <= rom_array(6825);
		when "0001101010101010" => data_out <= rom_array(6826);
		when "0001101010101011" => data_out <= rom_array(6827);
		when "0001101010101100" => data_out <= rom_array(6828);
		when "0001101010101101" => data_out <= rom_array(6829);
		when "0001101010101110" => data_out <= rom_array(6830);
		when "0001101010101111" => data_out <= rom_array(6831);
		when "0001101010110000" => data_out <= rom_array(6832);
		when "0001101010110001" => data_out <= rom_array(6833);
		when "0001101010110010" => data_out <= rom_array(6834);
		when "0001101010110011" => data_out <= rom_array(6835);
		when "0001101010110100" => data_out <= rom_array(6836);
		when "0001101010110101" => data_out <= rom_array(6837);
		when "0001101010110110" => data_out <= rom_array(6838);
		when "0001101010110111" => data_out <= rom_array(6839);
		when "0001101010111000" => data_out <= rom_array(6840);
		when "0001101010111001" => data_out <= rom_array(6841);
		when "0001101010111010" => data_out <= rom_array(6842);
		when "0001101010111011" => data_out <= rom_array(6843);
		when "0001101010111100" => data_out <= rom_array(6844);
		when "0001101010111101" => data_out <= rom_array(6845);
		when "0001101010111110" => data_out <= rom_array(6846);
		when "0001101010111111" => data_out <= rom_array(6847);
		when "0001101011000000" => data_out <= rom_array(6848);
		when "0001101011000001" => data_out <= rom_array(6849);
		when "0001101011000010" => data_out <= rom_array(6850);
		when "0001101011000011" => data_out <= rom_array(6851);
		when "0001101011000100" => data_out <= rom_array(6852);
		when "0001101011000101" => data_out <= rom_array(6853);
		when "0001101011000110" => data_out <= rom_array(6854);
		when "0001101011000111" => data_out <= rom_array(6855);
		when "0001101011001000" => data_out <= rom_array(6856);
		when "0001101011001001" => data_out <= rom_array(6857);
		when "0001101011001010" => data_out <= rom_array(6858);
		when "0001101011001011" => data_out <= rom_array(6859);
		when "0001101011001100" => data_out <= rom_array(6860);
		when "0001101011001101" => data_out <= rom_array(6861);
		when "0001101011001110" => data_out <= rom_array(6862);
		when "0001101011001111" => data_out <= rom_array(6863);
		when "0001101011010000" => data_out <= rom_array(6864);
		when "0001101011010001" => data_out <= rom_array(6865);
		when "0001101011010010" => data_out <= rom_array(6866);
		when "0001101011010011" => data_out <= rom_array(6867);
		when "0001101011010100" => data_out <= rom_array(6868);
		when "0001101011010101" => data_out <= rom_array(6869);
		when "0001101011010110" => data_out <= rom_array(6870);
		when "0001101011010111" => data_out <= rom_array(6871);
		when "0001101011011000" => data_out <= rom_array(6872);
		when "0001101011011001" => data_out <= rom_array(6873);
		when "0001101011011010" => data_out <= rom_array(6874);
		when "0001101011011011" => data_out <= rom_array(6875);
		when "0001101011011100" => data_out <= rom_array(6876);
		when "0001101011011101" => data_out <= rom_array(6877);
		when "0001101011011110" => data_out <= rom_array(6878);
		when "0001101011011111" => data_out <= rom_array(6879);
		when "0001101011100000" => data_out <= rom_array(6880);
		when "0001101011100001" => data_out <= rom_array(6881);
		when "0001101011100010" => data_out <= rom_array(6882);
		when "0001101011100011" => data_out <= rom_array(6883);
		when "0001101011100100" => data_out <= rom_array(6884);
		when "0001101011100101" => data_out <= rom_array(6885);
		when "0001101011100110" => data_out <= rom_array(6886);
		when "0001101011100111" => data_out <= rom_array(6887);
		when "0001101011101000" => data_out <= rom_array(6888);
		when "0001101011101001" => data_out <= rom_array(6889);
		when "0001101011101010" => data_out <= rom_array(6890);
		when "0001101011101011" => data_out <= rom_array(6891);
		when "0001101011101100" => data_out <= rom_array(6892);
		when "0001101011101101" => data_out <= rom_array(6893);
		when "0001101011101110" => data_out <= rom_array(6894);
		when "0001101011101111" => data_out <= rom_array(6895);
		when "0001101011110000" => data_out <= rom_array(6896);
		when "0001101011110001" => data_out <= rom_array(6897);
		when "0001101011110010" => data_out <= rom_array(6898);
		when "0001101011110011" => data_out <= rom_array(6899);
		when "0001101011110100" => data_out <= rom_array(6900);
		when "0001101011110101" => data_out <= rom_array(6901);
		when "0001101011110110" => data_out <= rom_array(6902);
		when "0001101011110111" => data_out <= rom_array(6903);
		when "0001101011111000" => data_out <= rom_array(6904);
		when "0001101011111001" => data_out <= rom_array(6905);
		when "0001101011111010" => data_out <= rom_array(6906);
		when "0001101011111011" => data_out <= rom_array(6907);
		when "0001101011111100" => data_out <= rom_array(6908);
		when "0001101011111101" => data_out <= rom_array(6909);
		when "0001101011111110" => data_out <= rom_array(6910);
		when "0001101011111111" => data_out <= rom_array(6911);
		when "0001101100000000" => data_out <= rom_array(6912);
		when "0001101100000001" => data_out <= rom_array(6913);
		when "0001101100000010" => data_out <= rom_array(6914);
		when "0001101100000011" => data_out <= rom_array(6915);
		when "0001101100000100" => data_out <= rom_array(6916);
		when "0001101100000101" => data_out <= rom_array(6917);
		when "0001101100000110" => data_out <= rom_array(6918);
		when "0001101100000111" => data_out <= rom_array(6919);
		when "0001101100001000" => data_out <= rom_array(6920);
		when "0001101100001001" => data_out <= rom_array(6921);
		when "0001101100001010" => data_out <= rom_array(6922);
		when "0001101100001011" => data_out <= rom_array(6923);
		when "0001101100001100" => data_out <= rom_array(6924);
		when "0001101100001101" => data_out <= rom_array(6925);
		when "0001101100001110" => data_out <= rom_array(6926);
		when "0001101100001111" => data_out <= rom_array(6927);
		when "0001101100010000" => data_out <= rom_array(6928);
		when "0001101100010001" => data_out <= rom_array(6929);
		when "0001101100010010" => data_out <= rom_array(6930);
		when "0001101100010011" => data_out <= rom_array(6931);
		when "0001101100010100" => data_out <= rom_array(6932);
		when "0001101100010101" => data_out <= rom_array(6933);
		when "0001101100010110" => data_out <= rom_array(6934);
		when "0001101100010111" => data_out <= rom_array(6935);
		when "0001101100011000" => data_out <= rom_array(6936);
		when "0001101100011001" => data_out <= rom_array(6937);
		when "0001101100011010" => data_out <= rom_array(6938);
		when "0001101100011011" => data_out <= rom_array(6939);
		when "0001101100011100" => data_out <= rom_array(6940);
		when "0001101100011101" => data_out <= rom_array(6941);
		when "0001101100011110" => data_out <= rom_array(6942);
		when "0001101100011111" => data_out <= rom_array(6943);
		when "0001101100100000" => data_out <= rom_array(6944);
		when "0001101100100001" => data_out <= rom_array(6945);
		when "0001101100100010" => data_out <= rom_array(6946);
		when "0001101100100011" => data_out <= rom_array(6947);
		when "0001101100100100" => data_out <= rom_array(6948);
		when "0001101100100101" => data_out <= rom_array(6949);
		when "0001101100100110" => data_out <= rom_array(6950);
		when "0001101100100111" => data_out <= rom_array(6951);
		when "0001101100101000" => data_out <= rom_array(6952);
		when "0001101100101001" => data_out <= rom_array(6953);
		when "0001101100101010" => data_out <= rom_array(6954);
		when "0001101100101011" => data_out <= rom_array(6955);
		when "0001101100101100" => data_out <= rom_array(6956);
		when "0001101100101101" => data_out <= rom_array(6957);
		when "0001101100101110" => data_out <= rom_array(6958);
		when "0001101100101111" => data_out <= rom_array(6959);
		when "0001101100110000" => data_out <= rom_array(6960);
		when "0001101100110001" => data_out <= rom_array(6961);
		when "0001101100110010" => data_out <= rom_array(6962);
		when "0001101100110011" => data_out <= rom_array(6963);
		when "0001101100110100" => data_out <= rom_array(6964);
		when "0001101100110101" => data_out <= rom_array(6965);
		when "0001101100110110" => data_out <= rom_array(6966);
		when "0001101100110111" => data_out <= rom_array(6967);
		when "0001101100111000" => data_out <= rom_array(6968);
		when "0001101100111001" => data_out <= rom_array(6969);
		when "0001101100111010" => data_out <= rom_array(6970);
		when "0001101100111011" => data_out <= rom_array(6971);
		when "0001101100111100" => data_out <= rom_array(6972);
		when "0001101100111101" => data_out <= rom_array(6973);
		when "0001101100111110" => data_out <= rom_array(6974);
		when "0001101100111111" => data_out <= rom_array(6975);
		when "0001101101000000" => data_out <= rom_array(6976);
		when "0001101101000001" => data_out <= rom_array(6977);
		when "0001101101000010" => data_out <= rom_array(6978);
		when "0001101101000011" => data_out <= rom_array(6979);
		when "0001101101000100" => data_out <= rom_array(6980);
		when "0001101101000101" => data_out <= rom_array(6981);
		when "0001101101000110" => data_out <= rom_array(6982);
		when "0001101101000111" => data_out <= rom_array(6983);
		when "0001101101001000" => data_out <= rom_array(6984);
		when "0001101101001001" => data_out <= rom_array(6985);
		when "0001101101001010" => data_out <= rom_array(6986);
		when "0001101101001011" => data_out <= rom_array(6987);
		when "0001101101001100" => data_out <= rom_array(6988);
		when "0001101101001101" => data_out <= rom_array(6989);
		when "0001101101001110" => data_out <= rom_array(6990);
		when "0001101101001111" => data_out <= rom_array(6991);
		when "0001101101010000" => data_out <= rom_array(6992);
		when "0001101101010001" => data_out <= rom_array(6993);
		when "0001101101010010" => data_out <= rom_array(6994);
		when "0001101101010011" => data_out <= rom_array(6995);
		when "0001101101010100" => data_out <= rom_array(6996);
		when "0001101101010101" => data_out <= rom_array(6997);
		when "0001101101010110" => data_out <= rom_array(6998);
		when "0001101101010111" => data_out <= rom_array(6999);
		when "0001101101011000" => data_out <= rom_array(7000);
		when "0001101101011001" => data_out <= rom_array(7001);
		when "0001101101011010" => data_out <= rom_array(7002);
		when "0001101101011011" => data_out <= rom_array(7003);
		when "0001101101011100" => data_out <= rom_array(7004);
		when "0001101101011101" => data_out <= rom_array(7005);
		when "0001101101011110" => data_out <= rom_array(7006);
		when "0001101101011111" => data_out <= rom_array(7007);
		when "0001101101100000" => data_out <= rom_array(7008);
		when "0001101101100001" => data_out <= rom_array(7009);
		when "0001101101100010" => data_out <= rom_array(7010);
		when "0001101101100011" => data_out <= rom_array(7011);
		when "0001101101100100" => data_out <= rom_array(7012);
		when "0001101101100101" => data_out <= rom_array(7013);
		when "0001101101100110" => data_out <= rom_array(7014);
		when "0001101101100111" => data_out <= rom_array(7015);
		when "0001101101101000" => data_out <= rom_array(7016);
		when "0001101101101001" => data_out <= rom_array(7017);
		when "0001101101101010" => data_out <= rom_array(7018);
		when "0001101101101011" => data_out <= rom_array(7019);
		when "0001101101101100" => data_out <= rom_array(7020);
		when "0001101101101101" => data_out <= rom_array(7021);
		when "0001101101101110" => data_out <= rom_array(7022);
		when "0001101101101111" => data_out <= rom_array(7023);
		when "0001101101110000" => data_out <= rom_array(7024);
		when "0001101101110001" => data_out <= rom_array(7025);
		when "0001101101110010" => data_out <= rom_array(7026);
		when "0001101101110011" => data_out <= rom_array(7027);
		when "0001101101110100" => data_out <= rom_array(7028);
		when "0001101101110101" => data_out <= rom_array(7029);
		when "0001101101110110" => data_out <= rom_array(7030);
		when "0001101101110111" => data_out <= rom_array(7031);
		when "0001101101111000" => data_out <= rom_array(7032);
		when "0001101101111001" => data_out <= rom_array(7033);
		when "0001101101111010" => data_out <= rom_array(7034);
		when "0001101101111011" => data_out <= rom_array(7035);
		when "0001101101111100" => data_out <= rom_array(7036);
		when "0001101101111101" => data_out <= rom_array(7037);
		when "0001101101111110" => data_out <= rom_array(7038);
		when "0001101101111111" => data_out <= rom_array(7039);
		when "0001101110000000" => data_out <= rom_array(7040);
		when "0001101110000001" => data_out <= rom_array(7041);
		when "0001101110000010" => data_out <= rom_array(7042);
		when "0001101110000011" => data_out <= rom_array(7043);
		when "0001101110000100" => data_out <= rom_array(7044);
		when "0001101110000101" => data_out <= rom_array(7045);
		when "0001101110000110" => data_out <= rom_array(7046);
		when "0001101110000111" => data_out <= rom_array(7047);
		when "0001101110001000" => data_out <= rom_array(7048);
		when "0001101110001001" => data_out <= rom_array(7049);
		when "0001101110001010" => data_out <= rom_array(7050);
		when "0001101110001011" => data_out <= rom_array(7051);
		when "0001101110001100" => data_out <= rom_array(7052);
		when "0001101110001101" => data_out <= rom_array(7053);
		when "0001101110001110" => data_out <= rom_array(7054);
		when "0001101110001111" => data_out <= rom_array(7055);
		when "0001101110010000" => data_out <= rom_array(7056);
		when "0001101110010001" => data_out <= rom_array(7057);
		when "0001101110010010" => data_out <= rom_array(7058);
		when "0001101110010011" => data_out <= rom_array(7059);
		when "0001101110010100" => data_out <= rom_array(7060);
		when "0001101110010101" => data_out <= rom_array(7061);
		when "0001101110010110" => data_out <= rom_array(7062);
		when "0001101110010111" => data_out <= rom_array(7063);
		when "0001101110011000" => data_out <= rom_array(7064);
		when "0001101110011001" => data_out <= rom_array(7065);
		when "0001101110011010" => data_out <= rom_array(7066);
		when "0001101110011011" => data_out <= rom_array(7067);
		when "0001101110011100" => data_out <= rom_array(7068);
		when "0001101110011101" => data_out <= rom_array(7069);
		when "0001101110011110" => data_out <= rom_array(7070);
		when "0001101110011111" => data_out <= rom_array(7071);
		when "0001101110100000" => data_out <= rom_array(7072);
		when "0001101110100001" => data_out <= rom_array(7073);
		when "0001101110100010" => data_out <= rom_array(7074);
		when "0001101110100011" => data_out <= rom_array(7075);
		when "0001101110100100" => data_out <= rom_array(7076);
		when "0001101110100101" => data_out <= rom_array(7077);
		when "0001101110100110" => data_out <= rom_array(7078);
		when "0001101110100111" => data_out <= rom_array(7079);
		when "0001101110101000" => data_out <= rom_array(7080);
		when "0001101110101001" => data_out <= rom_array(7081);
		when "0001101110101010" => data_out <= rom_array(7082);
		when "0001101110101011" => data_out <= rom_array(7083);
		when "0001101110101100" => data_out <= rom_array(7084);
		when "0001101110101101" => data_out <= rom_array(7085);
		when "0001101110101110" => data_out <= rom_array(7086);
		when "0001101110101111" => data_out <= rom_array(7087);
		when "0001101110110000" => data_out <= rom_array(7088);
		when "0001101110110001" => data_out <= rom_array(7089);
		when "0001101110110010" => data_out <= rom_array(7090);
		when "0001101110110011" => data_out <= rom_array(7091);
		when "0001101110110100" => data_out <= rom_array(7092);
		when "0001101110110101" => data_out <= rom_array(7093);
		when "0001101110110110" => data_out <= rom_array(7094);
		when "0001101110110111" => data_out <= rom_array(7095);
		when "0001101110111000" => data_out <= rom_array(7096);
		when "0001101110111001" => data_out <= rom_array(7097);
		when "0001101110111010" => data_out <= rom_array(7098);
		when "0001101110111011" => data_out <= rom_array(7099);
		when "0001101110111100" => data_out <= rom_array(7100);
		when "0001101110111101" => data_out <= rom_array(7101);
		when "0001101110111110" => data_out <= rom_array(7102);
		when "0001101110111111" => data_out <= rom_array(7103);
		when "0001101111000000" => data_out <= rom_array(7104);
		when "0001101111000001" => data_out <= rom_array(7105);
		when "0001101111000010" => data_out <= rom_array(7106);
		when "0001101111000011" => data_out <= rom_array(7107);
		when "0001101111000100" => data_out <= rom_array(7108);
		when "0001101111000101" => data_out <= rom_array(7109);
		when "0001101111000110" => data_out <= rom_array(7110);
		when "0001101111000111" => data_out <= rom_array(7111);
		when "0001101111001000" => data_out <= rom_array(7112);
		when "0001101111001001" => data_out <= rom_array(7113);
		when "0001101111001010" => data_out <= rom_array(7114);
		when "0001101111001011" => data_out <= rom_array(7115);
		when "0001101111001100" => data_out <= rom_array(7116);
		when "0001101111001101" => data_out <= rom_array(7117);
		when "0001101111001110" => data_out <= rom_array(7118);
		when "0001101111001111" => data_out <= rom_array(7119);
		when "0001101111010000" => data_out <= rom_array(7120);
		when "0001101111010001" => data_out <= rom_array(7121);
		when "0001101111010010" => data_out <= rom_array(7122);
		when "0001101111010011" => data_out <= rom_array(7123);
		when "0001101111010100" => data_out <= rom_array(7124);
		when "0001101111010101" => data_out <= rom_array(7125);
		when "0001101111010110" => data_out <= rom_array(7126);
		when "0001101111010111" => data_out <= rom_array(7127);
		when "0001101111011000" => data_out <= rom_array(7128);
		when "0001101111011001" => data_out <= rom_array(7129);
		when "0001101111011010" => data_out <= rom_array(7130);
		when "0001101111011011" => data_out <= rom_array(7131);
		when "0001101111011100" => data_out <= rom_array(7132);
		when "0001101111011101" => data_out <= rom_array(7133);
		when "0001101111011110" => data_out <= rom_array(7134);
		when "0001101111011111" => data_out <= rom_array(7135);
		when "0001101111100000" => data_out <= rom_array(7136);
		when "0001101111100001" => data_out <= rom_array(7137);
		when "0001101111100010" => data_out <= rom_array(7138);
		when "0001101111100011" => data_out <= rom_array(7139);
		when "0001101111100100" => data_out <= rom_array(7140);
		when "0001101111100101" => data_out <= rom_array(7141);
		when "0001101111100110" => data_out <= rom_array(7142);
		when "0001101111100111" => data_out <= rom_array(7143);
		when "0001101111101000" => data_out <= rom_array(7144);
		when "0001101111101001" => data_out <= rom_array(7145);
		when "0001101111101010" => data_out <= rom_array(7146);
		when "0001101111101011" => data_out <= rom_array(7147);
		when "0001101111101100" => data_out <= rom_array(7148);
		when "0001101111101101" => data_out <= rom_array(7149);
		when "0001101111101110" => data_out <= rom_array(7150);
		when "0001101111101111" => data_out <= rom_array(7151);
		when "0001101111110000" => data_out <= rom_array(7152);
		when "0001101111110001" => data_out <= rom_array(7153);
		when "0001101111110010" => data_out <= rom_array(7154);
		when "0001101111110011" => data_out <= rom_array(7155);
		when "0001101111110100" => data_out <= rom_array(7156);
		when "0001101111110101" => data_out <= rom_array(7157);
		when "0001101111110110" => data_out <= rom_array(7158);
		when "0001101111110111" => data_out <= rom_array(7159);
		when "0001101111111000" => data_out <= rom_array(7160);
		when "0001101111111001" => data_out <= rom_array(7161);
		when "0001101111111010" => data_out <= rom_array(7162);
		when "0001101111111011" => data_out <= rom_array(7163);
		when "0001101111111100" => data_out <= rom_array(7164);
		when "0001101111111101" => data_out <= rom_array(7165);
		when "0001101111111110" => data_out <= rom_array(7166);
		when "0001101111111111" => data_out <= rom_array(7167);
		when "0001110000000000" => data_out <= rom_array(7168);
		when "0001110000000001" => data_out <= rom_array(7169);
		when "0001110000000010" => data_out <= rom_array(7170);
		when "0001110000000011" => data_out <= rom_array(7171);
		when "0001110000000100" => data_out <= rom_array(7172);
		when "0001110000000101" => data_out <= rom_array(7173);
		when "0001110000000110" => data_out <= rom_array(7174);
		when "0001110000000111" => data_out <= rom_array(7175);
		when "0001110000001000" => data_out <= rom_array(7176);
		when "0001110000001001" => data_out <= rom_array(7177);
		when "0001110000001010" => data_out <= rom_array(7178);
		when "0001110000001011" => data_out <= rom_array(7179);
		when "0001110000001100" => data_out <= rom_array(7180);
		when "0001110000001101" => data_out <= rom_array(7181);
		when "0001110000001110" => data_out <= rom_array(7182);
		when "0001110000001111" => data_out <= rom_array(7183);
		when "0001110000010000" => data_out <= rom_array(7184);
		when "0001110000010001" => data_out <= rom_array(7185);
		when "0001110000010010" => data_out <= rom_array(7186);
		when "0001110000010011" => data_out <= rom_array(7187);
		when "0001110000010100" => data_out <= rom_array(7188);
		when "0001110000010101" => data_out <= rom_array(7189);
		when "0001110000010110" => data_out <= rom_array(7190);
		when "0001110000010111" => data_out <= rom_array(7191);
		when "0001110000011000" => data_out <= rom_array(7192);
		when "0001110000011001" => data_out <= rom_array(7193);
		when "0001110000011010" => data_out <= rom_array(7194);
		when "0001110000011011" => data_out <= rom_array(7195);
		when "0001110000011100" => data_out <= rom_array(7196);
		when "0001110000011101" => data_out <= rom_array(7197);
		when "0001110000011110" => data_out <= rom_array(7198);
		when "0001110000011111" => data_out <= rom_array(7199);
		when "0001110000100000" => data_out <= rom_array(7200);
		when "0001110000100001" => data_out <= rom_array(7201);
		when "0001110000100010" => data_out <= rom_array(7202);
		when "0001110000100011" => data_out <= rom_array(7203);
		when "0001110000100100" => data_out <= rom_array(7204);
		when "0001110000100101" => data_out <= rom_array(7205);
		when "0001110000100110" => data_out <= rom_array(7206);
		when "0001110000100111" => data_out <= rom_array(7207);
		when "0001110000101000" => data_out <= rom_array(7208);
		when "0001110000101001" => data_out <= rom_array(7209);
		when "0001110000101010" => data_out <= rom_array(7210);
		when "0001110000101011" => data_out <= rom_array(7211);
		when "0001110000101100" => data_out <= rom_array(7212);
		when "0001110000101101" => data_out <= rom_array(7213);
		when "0001110000101110" => data_out <= rom_array(7214);
		when "0001110000101111" => data_out <= rom_array(7215);
		when "0001110000110000" => data_out <= rom_array(7216);
		when "0001110000110001" => data_out <= rom_array(7217);
		when "0001110000110010" => data_out <= rom_array(7218);
		when "0001110000110011" => data_out <= rom_array(7219);
		when "0001110000110100" => data_out <= rom_array(7220);
		when "0001110000110101" => data_out <= rom_array(7221);
		when "0001110000110110" => data_out <= rom_array(7222);
		when "0001110000110111" => data_out <= rom_array(7223);
		when "0001110000111000" => data_out <= rom_array(7224);
		when "0001110000111001" => data_out <= rom_array(7225);
		when "0001110000111010" => data_out <= rom_array(7226);
		when "0001110000111011" => data_out <= rom_array(7227);
		when "0001110000111100" => data_out <= rom_array(7228);
		when "0001110000111101" => data_out <= rom_array(7229);
		when "0001110000111110" => data_out <= rom_array(7230);
		when "0001110000111111" => data_out <= rom_array(7231);
		when "0001110001000000" => data_out <= rom_array(7232);
		when "0001110001000001" => data_out <= rom_array(7233);
		when "0001110001000010" => data_out <= rom_array(7234);
		when "0001110001000011" => data_out <= rom_array(7235);
		when "0001110001000100" => data_out <= rom_array(7236);
		when "0001110001000101" => data_out <= rom_array(7237);
		when "0001110001000110" => data_out <= rom_array(7238);
		when "0001110001000111" => data_out <= rom_array(7239);
		when "0001110001001000" => data_out <= rom_array(7240);
		when "0001110001001001" => data_out <= rom_array(7241);
		when "0001110001001010" => data_out <= rom_array(7242);
		when "0001110001001011" => data_out <= rom_array(7243);
		when "0001110001001100" => data_out <= rom_array(7244);
		when "0001110001001101" => data_out <= rom_array(7245);
		when "0001110001001110" => data_out <= rom_array(7246);
		when "0001110001001111" => data_out <= rom_array(7247);
		when "0001110001010000" => data_out <= rom_array(7248);
		when "0001110001010001" => data_out <= rom_array(7249);
		when "0001110001010010" => data_out <= rom_array(7250);
		when "0001110001010011" => data_out <= rom_array(7251);
		when "0001110001010100" => data_out <= rom_array(7252);
		when "0001110001010101" => data_out <= rom_array(7253);
		when "0001110001010110" => data_out <= rom_array(7254);
		when "0001110001010111" => data_out <= rom_array(7255);
		when "0001110001011000" => data_out <= rom_array(7256);
		when "0001110001011001" => data_out <= rom_array(7257);
		when "0001110001011010" => data_out <= rom_array(7258);
		when "0001110001011011" => data_out <= rom_array(7259);
		when "0001110001011100" => data_out <= rom_array(7260);
		when "0001110001011101" => data_out <= rom_array(7261);
		when "0001110001011110" => data_out <= rom_array(7262);
		when "0001110001011111" => data_out <= rom_array(7263);
		when "0001110001100000" => data_out <= rom_array(7264);
		when "0001110001100001" => data_out <= rom_array(7265);
		when "0001110001100010" => data_out <= rom_array(7266);
		when "0001110001100011" => data_out <= rom_array(7267);
		when "0001110001100100" => data_out <= rom_array(7268);
		when "0001110001100101" => data_out <= rom_array(7269);
		when "0001110001100110" => data_out <= rom_array(7270);
		when "0001110001100111" => data_out <= rom_array(7271);
		when "0001110001101000" => data_out <= rom_array(7272);
		when "0001110001101001" => data_out <= rom_array(7273);
		when "0001110001101010" => data_out <= rom_array(7274);
		when "0001110001101011" => data_out <= rom_array(7275);
		when "0001110001101100" => data_out <= rom_array(7276);
		when "0001110001101101" => data_out <= rom_array(7277);
		when "0001110001101110" => data_out <= rom_array(7278);
		when "0001110001101111" => data_out <= rom_array(7279);
		when "0001110001110000" => data_out <= rom_array(7280);
		when "0001110001110001" => data_out <= rom_array(7281);
		when "0001110001110010" => data_out <= rom_array(7282);
		when "0001110001110011" => data_out <= rom_array(7283);
		when "0001110001110100" => data_out <= rom_array(7284);
		when "0001110001110101" => data_out <= rom_array(7285);
		when "0001110001110110" => data_out <= rom_array(7286);
		when "0001110001110111" => data_out <= rom_array(7287);
		when "0001110001111000" => data_out <= rom_array(7288);
		when "0001110001111001" => data_out <= rom_array(7289);
		when "0001110001111010" => data_out <= rom_array(7290);
		when "0001110001111011" => data_out <= rom_array(7291);
		when "0001110001111100" => data_out <= rom_array(7292);
		when "0001110001111101" => data_out <= rom_array(7293);
		when "0001110001111110" => data_out <= rom_array(7294);
		when "0001110001111111" => data_out <= rom_array(7295);
		when "0001110010000000" => data_out <= rom_array(7296);
		when "0001110010000001" => data_out <= rom_array(7297);
		when "0001110010000010" => data_out <= rom_array(7298);
		when "0001110010000011" => data_out <= rom_array(7299);
		when "0001110010000100" => data_out <= rom_array(7300);
		when "0001110010000101" => data_out <= rom_array(7301);
		when "0001110010000110" => data_out <= rom_array(7302);
		when "0001110010000111" => data_out <= rom_array(7303);
		when "0001110010001000" => data_out <= rom_array(7304);
		when "0001110010001001" => data_out <= rom_array(7305);
		when "0001110010001010" => data_out <= rom_array(7306);
		when "0001110010001011" => data_out <= rom_array(7307);
		when "0001110010001100" => data_out <= rom_array(7308);
		when "0001110010001101" => data_out <= rom_array(7309);
		when "0001110010001110" => data_out <= rom_array(7310);
		when "0001110010001111" => data_out <= rom_array(7311);
		when "0001110010010000" => data_out <= rom_array(7312);
		when "0001110010010001" => data_out <= rom_array(7313);
		when "0001110010010010" => data_out <= rom_array(7314);
		when "0001110010010011" => data_out <= rom_array(7315);
		when "0001110010010100" => data_out <= rom_array(7316);
		when "0001110010010101" => data_out <= rom_array(7317);
		when "0001110010010110" => data_out <= rom_array(7318);
		when "0001110010010111" => data_out <= rom_array(7319);
		when "0001110010011000" => data_out <= rom_array(7320);
		when "0001110010011001" => data_out <= rom_array(7321);
		when "0001110010011010" => data_out <= rom_array(7322);
		when "0001110010011011" => data_out <= rom_array(7323);
		when "0001110010011100" => data_out <= rom_array(7324);
		when "0001110010011101" => data_out <= rom_array(7325);
		when "0001110010011110" => data_out <= rom_array(7326);
		when "0001110010011111" => data_out <= rom_array(7327);
		when "0001110010100000" => data_out <= rom_array(7328);
		when "0001110010100001" => data_out <= rom_array(7329);
		when "0001110010100010" => data_out <= rom_array(7330);
		when "0001110010100011" => data_out <= rom_array(7331);
		when "0001110010100100" => data_out <= rom_array(7332);
		when "0001110010100101" => data_out <= rom_array(7333);
		when "0001110010100110" => data_out <= rom_array(7334);
		when "0001110010100111" => data_out <= rom_array(7335);
		when "0001110010101000" => data_out <= rom_array(7336);
		when "0001110010101001" => data_out <= rom_array(7337);
		when "0001110010101010" => data_out <= rom_array(7338);
		when "0001110010101011" => data_out <= rom_array(7339);
		when "0001110010101100" => data_out <= rom_array(7340);
		when "0001110010101101" => data_out <= rom_array(7341);
		when "0001110010101110" => data_out <= rom_array(7342);
		when "0001110010101111" => data_out <= rom_array(7343);
		when "0001110010110000" => data_out <= rom_array(7344);
		when "0001110010110001" => data_out <= rom_array(7345);
		when "0001110010110010" => data_out <= rom_array(7346);
		when "0001110010110011" => data_out <= rom_array(7347);
		when "0001110010110100" => data_out <= rom_array(7348);
		when "0001110010110101" => data_out <= rom_array(7349);
		when "0001110010110110" => data_out <= rom_array(7350);
		when "0001110010110111" => data_out <= rom_array(7351);
		when "0001110010111000" => data_out <= rom_array(7352);
		when "0001110010111001" => data_out <= rom_array(7353);
		when "0001110010111010" => data_out <= rom_array(7354);
		when "0001110010111011" => data_out <= rom_array(7355);
		when "0001110010111100" => data_out <= rom_array(7356);
		when "0001110010111101" => data_out <= rom_array(7357);
		when "0001110010111110" => data_out <= rom_array(7358);
		when "0001110010111111" => data_out <= rom_array(7359);
		when "0001110011000000" => data_out <= rom_array(7360);
		when "0001110011000001" => data_out <= rom_array(7361);
		when "0001110011000010" => data_out <= rom_array(7362);
		when "0001110011000011" => data_out <= rom_array(7363);
		when "0001110011000100" => data_out <= rom_array(7364);
		when "0001110011000101" => data_out <= rom_array(7365);
		when "0001110011000110" => data_out <= rom_array(7366);
		when "0001110011000111" => data_out <= rom_array(7367);
		when "0001110011001000" => data_out <= rom_array(7368);
		when "0001110011001001" => data_out <= rom_array(7369);
		when "0001110011001010" => data_out <= rom_array(7370);
		when "0001110011001011" => data_out <= rom_array(7371);
		when "0001110011001100" => data_out <= rom_array(7372);
		when "0001110011001101" => data_out <= rom_array(7373);
		when "0001110011001110" => data_out <= rom_array(7374);
		when "0001110011001111" => data_out <= rom_array(7375);
		when "0001110011010000" => data_out <= rom_array(7376);
		when "0001110011010001" => data_out <= rom_array(7377);
		when "0001110011010010" => data_out <= rom_array(7378);
		when "0001110011010011" => data_out <= rom_array(7379);
		when "0001110011010100" => data_out <= rom_array(7380);
		when "0001110011010101" => data_out <= rom_array(7381);
		when "0001110011010110" => data_out <= rom_array(7382);
		when "0001110011010111" => data_out <= rom_array(7383);
		when "0001110011011000" => data_out <= rom_array(7384);
		when "0001110011011001" => data_out <= rom_array(7385);
		when "0001110011011010" => data_out <= rom_array(7386);
		when "0001110011011011" => data_out <= rom_array(7387);
		when "0001110011011100" => data_out <= rom_array(7388);
		when "0001110011011101" => data_out <= rom_array(7389);
		when "0001110011011110" => data_out <= rom_array(7390);
		when "0001110011011111" => data_out <= rom_array(7391);
		when "0001110011100000" => data_out <= rom_array(7392);
		when "0001110011100001" => data_out <= rom_array(7393);
		when "0001110011100010" => data_out <= rom_array(7394);
		when "0001110011100011" => data_out <= rom_array(7395);
		when "0001110011100100" => data_out <= rom_array(7396);
		when "0001110011100101" => data_out <= rom_array(7397);
		when "0001110011100110" => data_out <= rom_array(7398);
		when "0001110011100111" => data_out <= rom_array(7399);
		when "0001110011101000" => data_out <= rom_array(7400);
		when "0001110011101001" => data_out <= rom_array(7401);
		when "0001110011101010" => data_out <= rom_array(7402);
		when "0001110011101011" => data_out <= rom_array(7403);
		when "0001110011101100" => data_out <= rom_array(7404);
		when "0001110011101101" => data_out <= rom_array(7405);
		when "0001110011101110" => data_out <= rom_array(7406);
		when "0001110011101111" => data_out <= rom_array(7407);
		when "0001110011110000" => data_out <= rom_array(7408);
		when "0001110011110001" => data_out <= rom_array(7409);
		when "0001110011110010" => data_out <= rom_array(7410);
		when "0001110011110011" => data_out <= rom_array(7411);
		when "0001110011110100" => data_out <= rom_array(7412);
		when "0001110011110101" => data_out <= rom_array(7413);
		when "0001110011110110" => data_out <= rom_array(7414);
		when "0001110011110111" => data_out <= rom_array(7415);
		when "0001110011111000" => data_out <= rom_array(7416);
		when "0001110011111001" => data_out <= rom_array(7417);
		when "0001110011111010" => data_out <= rom_array(7418);
		when "0001110011111011" => data_out <= rom_array(7419);
		when "0001110011111100" => data_out <= rom_array(7420);
		when "0001110011111101" => data_out <= rom_array(7421);
		when "0001110011111110" => data_out <= rom_array(7422);
		when "0001110011111111" => data_out <= rom_array(7423);
		when "0001110100000000" => data_out <= rom_array(7424);
		when "0001110100000001" => data_out <= rom_array(7425);
		when "0001110100000010" => data_out <= rom_array(7426);
		when "0001110100000011" => data_out <= rom_array(7427);
		when "0001110100000100" => data_out <= rom_array(7428);
		when "0001110100000101" => data_out <= rom_array(7429);
		when "0001110100000110" => data_out <= rom_array(7430);
		when "0001110100000111" => data_out <= rom_array(7431);
		when "0001110100001000" => data_out <= rom_array(7432);
		when "0001110100001001" => data_out <= rom_array(7433);
		when "0001110100001010" => data_out <= rom_array(7434);
		when "0001110100001011" => data_out <= rom_array(7435);
		when "0001110100001100" => data_out <= rom_array(7436);
		when "0001110100001101" => data_out <= rom_array(7437);
		when "0001110100001110" => data_out <= rom_array(7438);
		when "0001110100001111" => data_out <= rom_array(7439);
		when "0001110100010000" => data_out <= rom_array(7440);
		when "0001110100010001" => data_out <= rom_array(7441);
		when "0001110100010010" => data_out <= rom_array(7442);
		when "0001110100010011" => data_out <= rom_array(7443);
		when "0001110100010100" => data_out <= rom_array(7444);
		when "0001110100010101" => data_out <= rom_array(7445);
		when "0001110100010110" => data_out <= rom_array(7446);
		when "0001110100010111" => data_out <= rom_array(7447);
		when "0001110100011000" => data_out <= rom_array(7448);
		when "0001110100011001" => data_out <= rom_array(7449);
		when "0001110100011010" => data_out <= rom_array(7450);
		when "0001110100011011" => data_out <= rom_array(7451);
		when "0001110100011100" => data_out <= rom_array(7452);
		when "0001110100011101" => data_out <= rom_array(7453);
		when "0001110100011110" => data_out <= rom_array(7454);
		when "0001110100011111" => data_out <= rom_array(7455);
		when "0001110100100000" => data_out <= rom_array(7456);
		when "0001110100100001" => data_out <= rom_array(7457);
		when "0001110100100010" => data_out <= rom_array(7458);
		when "0001110100100011" => data_out <= rom_array(7459);
		when "0001110100100100" => data_out <= rom_array(7460);
		when "0001110100100101" => data_out <= rom_array(7461);
		when "0001110100100110" => data_out <= rom_array(7462);
		when "0001110100100111" => data_out <= rom_array(7463);
		when "0001110100101000" => data_out <= rom_array(7464);
		when "0001110100101001" => data_out <= rom_array(7465);
		when "0001110100101010" => data_out <= rom_array(7466);
		when "0001110100101011" => data_out <= rom_array(7467);
		when "0001110100101100" => data_out <= rom_array(7468);
		when "0001110100101101" => data_out <= rom_array(7469);
		when "0001110100101110" => data_out <= rom_array(7470);
		when "0001110100101111" => data_out <= rom_array(7471);
		when "0001110100110000" => data_out <= rom_array(7472);
		when "0001110100110001" => data_out <= rom_array(7473);
		when "0001110100110010" => data_out <= rom_array(7474);
		when "0001110100110011" => data_out <= rom_array(7475);
		when "0001110100110100" => data_out <= rom_array(7476);
		when "0001110100110101" => data_out <= rom_array(7477);
		when "0001110100110110" => data_out <= rom_array(7478);
		when "0001110100110111" => data_out <= rom_array(7479);
		when "0001110100111000" => data_out <= rom_array(7480);
		when "0001110100111001" => data_out <= rom_array(7481);
		when "0001110100111010" => data_out <= rom_array(7482);
		when "0001110100111011" => data_out <= rom_array(7483);
		when "0001110100111100" => data_out <= rom_array(7484);
		when "0001110100111101" => data_out <= rom_array(7485);
		when "0001110100111110" => data_out <= rom_array(7486);
		when "0001110100111111" => data_out <= rom_array(7487);
		when "0001110101000000" => data_out <= rom_array(7488);
		when "0001110101000001" => data_out <= rom_array(7489);
		when "0001110101000010" => data_out <= rom_array(7490);
		when "0001110101000011" => data_out <= rom_array(7491);
		when "0001110101000100" => data_out <= rom_array(7492);
		when "0001110101000101" => data_out <= rom_array(7493);
		when "0001110101000110" => data_out <= rom_array(7494);
		when "0001110101000111" => data_out <= rom_array(7495);
		when "0001110101001000" => data_out <= rom_array(7496);
		when "0001110101001001" => data_out <= rom_array(7497);
		when "0001110101001010" => data_out <= rom_array(7498);
		when "0001110101001011" => data_out <= rom_array(7499);
		when "0001110101001100" => data_out <= rom_array(7500);
		when "0001110101001101" => data_out <= rom_array(7501);
		when "0001110101001110" => data_out <= rom_array(7502);
		when "0001110101001111" => data_out <= rom_array(7503);
		when "0001110101010000" => data_out <= rom_array(7504);
		when "0001110101010001" => data_out <= rom_array(7505);
		when "0001110101010010" => data_out <= rom_array(7506);
		when "0001110101010011" => data_out <= rom_array(7507);
		when "0001110101010100" => data_out <= rom_array(7508);
		when "0001110101010101" => data_out <= rom_array(7509);
		when "0001110101010110" => data_out <= rom_array(7510);
		when "0001110101010111" => data_out <= rom_array(7511);
		when "0001110101011000" => data_out <= rom_array(7512);
		when "0001110101011001" => data_out <= rom_array(7513);
		when "0001110101011010" => data_out <= rom_array(7514);
		when "0001110101011011" => data_out <= rom_array(7515);
		when "0001110101011100" => data_out <= rom_array(7516);
		when "0001110101011101" => data_out <= rom_array(7517);
		when "0001110101011110" => data_out <= rom_array(7518);
		when "0001110101011111" => data_out <= rom_array(7519);
		when "0001110101100000" => data_out <= rom_array(7520);
		when "0001110101100001" => data_out <= rom_array(7521);
		when "0001110101100010" => data_out <= rom_array(7522);
		when "0001110101100011" => data_out <= rom_array(7523);
		when "0001110101100100" => data_out <= rom_array(7524);
		when "0001110101100101" => data_out <= rom_array(7525);
		when "0001110101100110" => data_out <= rom_array(7526);
		when "0001110101100111" => data_out <= rom_array(7527);
		when "0001110101101000" => data_out <= rom_array(7528);
		when "0001110101101001" => data_out <= rom_array(7529);
		when "0001110101101010" => data_out <= rom_array(7530);
		when "0001110101101011" => data_out <= rom_array(7531);
		when "0001110101101100" => data_out <= rom_array(7532);
		when "0001110101101101" => data_out <= rom_array(7533);
		when "0001110101101110" => data_out <= rom_array(7534);
		when "0001110101101111" => data_out <= rom_array(7535);
		when "0001110101110000" => data_out <= rom_array(7536);
		when "0001110101110001" => data_out <= rom_array(7537);
		when "0001110101110010" => data_out <= rom_array(7538);
		when "0001110101110011" => data_out <= rom_array(7539);
		when "0001110101110100" => data_out <= rom_array(7540);
		when "0001110101110101" => data_out <= rom_array(7541);
		when "0001110101110110" => data_out <= rom_array(7542);
		when "0001110101110111" => data_out <= rom_array(7543);
		when "0001110101111000" => data_out <= rom_array(7544);
		when "0001110101111001" => data_out <= rom_array(7545);
		when "0001110101111010" => data_out <= rom_array(7546);
		when "0001110101111011" => data_out <= rom_array(7547);
		when "0001110101111100" => data_out <= rom_array(7548);
		when "0001110101111101" => data_out <= rom_array(7549);
		when "0001110101111110" => data_out <= rom_array(7550);
		when "0001110101111111" => data_out <= rom_array(7551);
		when "0001110110000000" => data_out <= rom_array(7552);
		when "0001110110000001" => data_out <= rom_array(7553);
		when "0001110110000010" => data_out <= rom_array(7554);
		when "0001110110000011" => data_out <= rom_array(7555);
		when "0001110110000100" => data_out <= rom_array(7556);
		when "0001110110000101" => data_out <= rom_array(7557);
		when "0001110110000110" => data_out <= rom_array(7558);
		when "0001110110000111" => data_out <= rom_array(7559);
		when "0001110110001000" => data_out <= rom_array(7560);
		when "0001110110001001" => data_out <= rom_array(7561);
		when "0001110110001010" => data_out <= rom_array(7562);
		when "0001110110001011" => data_out <= rom_array(7563);
		when "0001110110001100" => data_out <= rom_array(7564);
		when "0001110110001101" => data_out <= rom_array(7565);
		when "0001110110001110" => data_out <= rom_array(7566);
		when "0001110110001111" => data_out <= rom_array(7567);
		when "0001110110010000" => data_out <= rom_array(7568);
		when "0001110110010001" => data_out <= rom_array(7569);
		when "0001110110010010" => data_out <= rom_array(7570);
		when "0001110110010011" => data_out <= rom_array(7571);
		when "0001110110010100" => data_out <= rom_array(7572);
		when "0001110110010101" => data_out <= rom_array(7573);
		when "0001110110010110" => data_out <= rom_array(7574);
		when "0001110110010111" => data_out <= rom_array(7575);
		when "0001110110011000" => data_out <= rom_array(7576);
		when "0001110110011001" => data_out <= rom_array(7577);
		when "0001110110011010" => data_out <= rom_array(7578);
		when "0001110110011011" => data_out <= rom_array(7579);
		when "0001110110011100" => data_out <= rom_array(7580);
		when "0001110110011101" => data_out <= rom_array(7581);
		when "0001110110011110" => data_out <= rom_array(7582);
		when "0001110110011111" => data_out <= rom_array(7583);
		when "0001110110100000" => data_out <= rom_array(7584);
		when "0001110110100001" => data_out <= rom_array(7585);
		when "0001110110100010" => data_out <= rom_array(7586);
		when "0001110110100011" => data_out <= rom_array(7587);
		when "0001110110100100" => data_out <= rom_array(7588);
		when "0001110110100101" => data_out <= rom_array(7589);
		when "0001110110100110" => data_out <= rom_array(7590);
		when "0001110110100111" => data_out <= rom_array(7591);
		when "0001110110101000" => data_out <= rom_array(7592);
		when "0001110110101001" => data_out <= rom_array(7593);
		when "0001110110101010" => data_out <= rom_array(7594);
		when "0001110110101011" => data_out <= rom_array(7595);
		when "0001110110101100" => data_out <= rom_array(7596);
		when "0001110110101101" => data_out <= rom_array(7597);
		when "0001110110101110" => data_out <= rom_array(7598);
		when "0001110110101111" => data_out <= rom_array(7599);
		when "0001110110110000" => data_out <= rom_array(7600);
		when "0001110110110001" => data_out <= rom_array(7601);
		when "0001110110110010" => data_out <= rom_array(7602);
		when "0001110110110011" => data_out <= rom_array(7603);
		when "0001110110110100" => data_out <= rom_array(7604);
		when "0001110110110101" => data_out <= rom_array(7605);
		when "0001110110110110" => data_out <= rom_array(7606);
		when "0001110110110111" => data_out <= rom_array(7607);
		when "0001110110111000" => data_out <= rom_array(7608);
		when "0001110110111001" => data_out <= rom_array(7609);
		when "0001110110111010" => data_out <= rom_array(7610);
		when "0001110110111011" => data_out <= rom_array(7611);
		when "0001110110111100" => data_out <= rom_array(7612);
		when "0001110110111101" => data_out <= rom_array(7613);
		when "0001110110111110" => data_out <= rom_array(7614);
		when "0001110110111111" => data_out <= rom_array(7615);
		when "0001110111000000" => data_out <= rom_array(7616);
		when "0001110111000001" => data_out <= rom_array(7617);
		when "0001110111000010" => data_out <= rom_array(7618);
		when "0001110111000011" => data_out <= rom_array(7619);
		when "0001110111000100" => data_out <= rom_array(7620);
		when "0001110111000101" => data_out <= rom_array(7621);
		when "0001110111000110" => data_out <= rom_array(7622);
		when "0001110111000111" => data_out <= rom_array(7623);
		when "0001110111001000" => data_out <= rom_array(7624);
		when "0001110111001001" => data_out <= rom_array(7625);
		when "0001110111001010" => data_out <= rom_array(7626);
		when "0001110111001011" => data_out <= rom_array(7627);
		when "0001110111001100" => data_out <= rom_array(7628);
		when "0001110111001101" => data_out <= rom_array(7629);
		when "0001110111001110" => data_out <= rom_array(7630);
		when "0001110111001111" => data_out <= rom_array(7631);
		when "0001110111010000" => data_out <= rom_array(7632);
		when "0001110111010001" => data_out <= rom_array(7633);
		when "0001110111010010" => data_out <= rom_array(7634);
		when "0001110111010011" => data_out <= rom_array(7635);
		when "0001110111010100" => data_out <= rom_array(7636);
		when "0001110111010101" => data_out <= rom_array(7637);
		when "0001110111010110" => data_out <= rom_array(7638);
		when "0001110111010111" => data_out <= rom_array(7639);
		when "0001110111011000" => data_out <= rom_array(7640);
		when "0001110111011001" => data_out <= rom_array(7641);
		when "0001110111011010" => data_out <= rom_array(7642);
		when "0001110111011011" => data_out <= rom_array(7643);
		when "0001110111011100" => data_out <= rom_array(7644);
		when "0001110111011101" => data_out <= rom_array(7645);
		when "0001110111011110" => data_out <= rom_array(7646);
		when "0001110111011111" => data_out <= rom_array(7647);
		when "0001110111100000" => data_out <= rom_array(7648);
		when "0001110111100001" => data_out <= rom_array(7649);
		when "0001110111100010" => data_out <= rom_array(7650);
		when "0001110111100011" => data_out <= rom_array(7651);
		when "0001110111100100" => data_out <= rom_array(7652);
		when "0001110111100101" => data_out <= rom_array(7653);
		when "0001110111100110" => data_out <= rom_array(7654);
		when "0001110111100111" => data_out <= rom_array(7655);
		when "0001110111101000" => data_out <= rom_array(7656);
		when "0001110111101001" => data_out <= rom_array(7657);
		when "0001110111101010" => data_out <= rom_array(7658);
		when "0001110111101011" => data_out <= rom_array(7659);
		when "0001110111101100" => data_out <= rom_array(7660);
		when "0001110111101101" => data_out <= rom_array(7661);
		when "0001110111101110" => data_out <= rom_array(7662);
		when "0001110111101111" => data_out <= rom_array(7663);
		when "0001110111110000" => data_out <= rom_array(7664);
		when "0001110111110001" => data_out <= rom_array(7665);
		when "0001110111110010" => data_out <= rom_array(7666);
		when "0001110111110011" => data_out <= rom_array(7667);
		when "0001110111110100" => data_out <= rom_array(7668);
		when "0001110111110101" => data_out <= rom_array(7669);
		when "0001110111110110" => data_out <= rom_array(7670);
		when "0001110111110111" => data_out <= rom_array(7671);
		when "0001110111111000" => data_out <= rom_array(7672);
		when "0001110111111001" => data_out <= rom_array(7673);
		when "0001110111111010" => data_out <= rom_array(7674);
		when "0001110111111011" => data_out <= rom_array(7675);
		when "0001110111111100" => data_out <= rom_array(7676);
		when "0001110111111101" => data_out <= rom_array(7677);
		when "0001110111111110" => data_out <= rom_array(7678);
		when "0001110111111111" => data_out <= rom_array(7679);
		when "0001111000000000" => data_out <= rom_array(7680);
		when "0001111000000001" => data_out <= rom_array(7681);
		when "0001111000000010" => data_out <= rom_array(7682);
		when "0001111000000011" => data_out <= rom_array(7683);
		when "0001111000000100" => data_out <= rom_array(7684);
		when "0001111000000101" => data_out <= rom_array(7685);
		when "0001111000000110" => data_out <= rom_array(7686);
		when "0001111000000111" => data_out <= rom_array(7687);
		when "0001111000001000" => data_out <= rom_array(7688);
		when "0001111000001001" => data_out <= rom_array(7689);
		when "0001111000001010" => data_out <= rom_array(7690);
		when "0001111000001011" => data_out <= rom_array(7691);
		when "0001111000001100" => data_out <= rom_array(7692);
		when "0001111000001101" => data_out <= rom_array(7693);
		when "0001111000001110" => data_out <= rom_array(7694);
		when "0001111000001111" => data_out <= rom_array(7695);
		when "0001111000010000" => data_out <= rom_array(7696);
		when "0001111000010001" => data_out <= rom_array(7697);
		when "0001111000010010" => data_out <= rom_array(7698);
		when "0001111000010011" => data_out <= rom_array(7699);
		when "0001111000010100" => data_out <= rom_array(7700);
		when "0001111000010101" => data_out <= rom_array(7701);
		when "0001111000010110" => data_out <= rom_array(7702);
		when "0001111000010111" => data_out <= rom_array(7703);
		when "0001111000011000" => data_out <= rom_array(7704);
		when "0001111000011001" => data_out <= rom_array(7705);
		when "0001111000011010" => data_out <= rom_array(7706);
		when "0001111000011011" => data_out <= rom_array(7707);
		when "0001111000011100" => data_out <= rom_array(7708);
		when "0001111000011101" => data_out <= rom_array(7709);
		when "0001111000011110" => data_out <= rom_array(7710);
		when "0001111000011111" => data_out <= rom_array(7711);
		when "0001111000100000" => data_out <= rom_array(7712);
		when "0001111000100001" => data_out <= rom_array(7713);
		when "0001111000100010" => data_out <= rom_array(7714);
		when "0001111000100011" => data_out <= rom_array(7715);
		when "0001111000100100" => data_out <= rom_array(7716);
		when "0001111000100101" => data_out <= rom_array(7717);
		when "0001111000100110" => data_out <= rom_array(7718);
		when "0001111000100111" => data_out <= rom_array(7719);
		when "0001111000101000" => data_out <= rom_array(7720);
		when "0001111000101001" => data_out <= rom_array(7721);
		when "0001111000101010" => data_out <= rom_array(7722);
		when "0001111000101011" => data_out <= rom_array(7723);
		when "0001111000101100" => data_out <= rom_array(7724);
		when "0001111000101101" => data_out <= rom_array(7725);
		when "0001111000101110" => data_out <= rom_array(7726);
		when "0001111000101111" => data_out <= rom_array(7727);
		when "0001111000110000" => data_out <= rom_array(7728);
		when "0001111000110001" => data_out <= rom_array(7729);
		when "0001111000110010" => data_out <= rom_array(7730);
		when "0001111000110011" => data_out <= rom_array(7731);
		when "0001111000110100" => data_out <= rom_array(7732);
		when "0001111000110101" => data_out <= rom_array(7733);
		when "0001111000110110" => data_out <= rom_array(7734);
		when "0001111000110111" => data_out <= rom_array(7735);
		when "0001111000111000" => data_out <= rom_array(7736);
		when "0001111000111001" => data_out <= rom_array(7737);
		when "0001111000111010" => data_out <= rom_array(7738);
		when "0001111000111011" => data_out <= rom_array(7739);
		when "0001111000111100" => data_out <= rom_array(7740);
		when "0001111000111101" => data_out <= rom_array(7741);
		when "0001111000111110" => data_out <= rom_array(7742);
		when "0001111000111111" => data_out <= rom_array(7743);
		when "0001111001000000" => data_out <= rom_array(7744);
		when "0001111001000001" => data_out <= rom_array(7745);
		when "0001111001000010" => data_out <= rom_array(7746);
		when "0001111001000011" => data_out <= rom_array(7747);
		when "0001111001000100" => data_out <= rom_array(7748);
		when "0001111001000101" => data_out <= rom_array(7749);
		when "0001111001000110" => data_out <= rom_array(7750);
		when "0001111001000111" => data_out <= rom_array(7751);
		when "0001111001001000" => data_out <= rom_array(7752);
		when "0001111001001001" => data_out <= rom_array(7753);
		when "0001111001001010" => data_out <= rom_array(7754);
		when "0001111001001011" => data_out <= rom_array(7755);
		when "0001111001001100" => data_out <= rom_array(7756);
		when "0001111001001101" => data_out <= rom_array(7757);
		when "0001111001001110" => data_out <= rom_array(7758);
		when "0001111001001111" => data_out <= rom_array(7759);
		when "0001111001010000" => data_out <= rom_array(7760);
		when "0001111001010001" => data_out <= rom_array(7761);
		when "0001111001010010" => data_out <= rom_array(7762);
		when "0001111001010011" => data_out <= rom_array(7763);
		when "0001111001010100" => data_out <= rom_array(7764);
		when "0001111001010101" => data_out <= rom_array(7765);
		when "0001111001010110" => data_out <= rom_array(7766);
		when "0001111001010111" => data_out <= rom_array(7767);
		when "0001111001011000" => data_out <= rom_array(7768);
		when "0001111001011001" => data_out <= rom_array(7769);
		when "0001111001011010" => data_out <= rom_array(7770);
		when "0001111001011011" => data_out <= rom_array(7771);
		when "0001111001011100" => data_out <= rom_array(7772);
		when "0001111001011101" => data_out <= rom_array(7773);
		when "0001111001011110" => data_out <= rom_array(7774);
		when "0001111001011111" => data_out <= rom_array(7775);
		when "0001111001100000" => data_out <= rom_array(7776);
		when "0001111001100001" => data_out <= rom_array(7777);
		when "0001111001100010" => data_out <= rom_array(7778);
		when "0001111001100011" => data_out <= rom_array(7779);
		when "0001111001100100" => data_out <= rom_array(7780);
		when "0001111001100101" => data_out <= rom_array(7781);
		when "0001111001100110" => data_out <= rom_array(7782);
		when "0001111001100111" => data_out <= rom_array(7783);
		when "0001111001101000" => data_out <= rom_array(7784);
		when "0001111001101001" => data_out <= rom_array(7785);
		when "0001111001101010" => data_out <= rom_array(7786);
		when "0001111001101011" => data_out <= rom_array(7787);
		when "0001111001101100" => data_out <= rom_array(7788);
		when "0001111001101101" => data_out <= rom_array(7789);
		when "0001111001101110" => data_out <= rom_array(7790);
		when "0001111001101111" => data_out <= rom_array(7791);
		when "0001111001110000" => data_out <= rom_array(7792);
		when "0001111001110001" => data_out <= rom_array(7793);
		when "0001111001110010" => data_out <= rom_array(7794);
		when "0001111001110011" => data_out <= rom_array(7795);
		when "0001111001110100" => data_out <= rom_array(7796);
		when "0001111001110101" => data_out <= rom_array(7797);
		when "0001111001110110" => data_out <= rom_array(7798);
		when "0001111001110111" => data_out <= rom_array(7799);
		when "0001111001111000" => data_out <= rom_array(7800);
		when "0001111001111001" => data_out <= rom_array(7801);
		when "0001111001111010" => data_out <= rom_array(7802);
		when "0001111001111011" => data_out <= rom_array(7803);
		when "0001111001111100" => data_out <= rom_array(7804);
		when "0001111001111101" => data_out <= rom_array(7805);
		when "0001111001111110" => data_out <= rom_array(7806);
		when "0001111001111111" => data_out <= rom_array(7807);
		when "0001111010000000" => data_out <= rom_array(7808);
		when "0001111010000001" => data_out <= rom_array(7809);
		when "0001111010000010" => data_out <= rom_array(7810);
		when "0001111010000011" => data_out <= rom_array(7811);
		when "0001111010000100" => data_out <= rom_array(7812);
		when "0001111010000101" => data_out <= rom_array(7813);
		when "0001111010000110" => data_out <= rom_array(7814);
		when "0001111010000111" => data_out <= rom_array(7815);
		when "0001111010001000" => data_out <= rom_array(7816);
		when "0001111010001001" => data_out <= rom_array(7817);
		when "0001111010001010" => data_out <= rom_array(7818);
		when "0001111010001011" => data_out <= rom_array(7819);
		when "0001111010001100" => data_out <= rom_array(7820);
		when "0001111010001101" => data_out <= rom_array(7821);
		when "0001111010001110" => data_out <= rom_array(7822);
		when "0001111010001111" => data_out <= rom_array(7823);
		when "0001111010010000" => data_out <= rom_array(7824);
		when "0001111010010001" => data_out <= rom_array(7825);
		when "0001111010010010" => data_out <= rom_array(7826);
		when "0001111010010011" => data_out <= rom_array(7827);
		when "0001111010010100" => data_out <= rom_array(7828);
		when "0001111010010101" => data_out <= rom_array(7829);
		when "0001111010010110" => data_out <= rom_array(7830);
		when "0001111010010111" => data_out <= rom_array(7831);
		when "0001111010011000" => data_out <= rom_array(7832);
		when "0001111010011001" => data_out <= rom_array(7833);
		when "0001111010011010" => data_out <= rom_array(7834);
		when "0001111010011011" => data_out <= rom_array(7835);
		when "0001111010011100" => data_out <= rom_array(7836);
		when "0001111010011101" => data_out <= rom_array(7837);
		when "0001111010011110" => data_out <= rom_array(7838);
		when "0001111010011111" => data_out <= rom_array(7839);
		when "0001111010100000" => data_out <= rom_array(7840);
		when "0001111010100001" => data_out <= rom_array(7841);
		when "0001111010100010" => data_out <= rom_array(7842);
		when "0001111010100011" => data_out <= rom_array(7843);
		when "0001111010100100" => data_out <= rom_array(7844);
		when "0001111010100101" => data_out <= rom_array(7845);
		when "0001111010100110" => data_out <= rom_array(7846);
		when "0001111010100111" => data_out <= rom_array(7847);
		when "0001111010101000" => data_out <= rom_array(7848);
		when "0001111010101001" => data_out <= rom_array(7849);
		when "0001111010101010" => data_out <= rom_array(7850);
		when "0001111010101011" => data_out <= rom_array(7851);
		when "0001111010101100" => data_out <= rom_array(7852);
		when "0001111010101101" => data_out <= rom_array(7853);
		when "0001111010101110" => data_out <= rom_array(7854);
		when "0001111010101111" => data_out <= rom_array(7855);
		when "0001111010110000" => data_out <= rom_array(7856);
		when "0001111010110001" => data_out <= rom_array(7857);
		when "0001111010110010" => data_out <= rom_array(7858);
		when "0001111010110011" => data_out <= rom_array(7859);
		when "0001111010110100" => data_out <= rom_array(7860);
		when "0001111010110101" => data_out <= rom_array(7861);
		when "0001111010110110" => data_out <= rom_array(7862);
		when "0001111010110111" => data_out <= rom_array(7863);
		when "0001111010111000" => data_out <= rom_array(7864);
		when "0001111010111001" => data_out <= rom_array(7865);
		when "0001111010111010" => data_out <= rom_array(7866);
		when "0001111010111011" => data_out <= rom_array(7867);
		when "0001111010111100" => data_out <= rom_array(7868);
		when "0001111010111101" => data_out <= rom_array(7869);
		when "0001111010111110" => data_out <= rom_array(7870);
		when "0001111010111111" => data_out <= rom_array(7871);
		when "0001111011000000" => data_out <= rom_array(7872);
		when "0001111011000001" => data_out <= rom_array(7873);
		when "0001111011000010" => data_out <= rom_array(7874);
		when "0001111011000011" => data_out <= rom_array(7875);
		when "0001111011000100" => data_out <= rom_array(7876);
		when "0001111011000101" => data_out <= rom_array(7877);
		when "0001111011000110" => data_out <= rom_array(7878);
		when "0001111011000111" => data_out <= rom_array(7879);
		when "0001111011001000" => data_out <= rom_array(7880);
		when "0001111011001001" => data_out <= rom_array(7881);
		when "0001111011001010" => data_out <= rom_array(7882);
		when "0001111011001011" => data_out <= rom_array(7883);
		when "0001111011001100" => data_out <= rom_array(7884);
		when "0001111011001101" => data_out <= rom_array(7885);
		when "0001111011001110" => data_out <= rom_array(7886);
		when "0001111011001111" => data_out <= rom_array(7887);
		when "0001111011010000" => data_out <= rom_array(7888);
		when "0001111011010001" => data_out <= rom_array(7889);
		when "0001111011010010" => data_out <= rom_array(7890);
		when "0001111011010011" => data_out <= rom_array(7891);
		when "0001111011010100" => data_out <= rom_array(7892);
		when "0001111011010101" => data_out <= rom_array(7893);
		when "0001111011010110" => data_out <= rom_array(7894);
		when "0001111011010111" => data_out <= rom_array(7895);
		when "0001111011011000" => data_out <= rom_array(7896);
		when "0001111011011001" => data_out <= rom_array(7897);
		when "0001111011011010" => data_out <= rom_array(7898);
		when "0001111011011011" => data_out <= rom_array(7899);
		when "0001111011011100" => data_out <= rom_array(7900);
		when "0001111011011101" => data_out <= rom_array(7901);
		when "0001111011011110" => data_out <= rom_array(7902);
		when "0001111011011111" => data_out <= rom_array(7903);
		when "0001111011100000" => data_out <= rom_array(7904);
		when "0001111011100001" => data_out <= rom_array(7905);
		when "0001111011100010" => data_out <= rom_array(7906);
		when "0001111011100011" => data_out <= rom_array(7907);
		when "0001111011100100" => data_out <= rom_array(7908);
		when "0001111011100101" => data_out <= rom_array(7909);
		when "0001111011100110" => data_out <= rom_array(7910);
		when "0001111011100111" => data_out <= rom_array(7911);
		when "0001111011101000" => data_out <= rom_array(7912);
		when "0001111011101001" => data_out <= rom_array(7913);
		when "0001111011101010" => data_out <= rom_array(7914);
		when "0001111011101011" => data_out <= rom_array(7915);
		when "0001111011101100" => data_out <= rom_array(7916);
		when "0001111011101101" => data_out <= rom_array(7917);
		when "0001111011101110" => data_out <= rom_array(7918);
		when "0001111011101111" => data_out <= rom_array(7919);
		when "0001111011110000" => data_out <= rom_array(7920);
		when "0001111011110001" => data_out <= rom_array(7921);
		when "0001111011110010" => data_out <= rom_array(7922);
		when "0001111011110011" => data_out <= rom_array(7923);
		when "0001111011110100" => data_out <= rom_array(7924);
		when "0001111011110101" => data_out <= rom_array(7925);
		when "0001111011110110" => data_out <= rom_array(7926);
		when "0001111011110111" => data_out <= rom_array(7927);
		when "0001111011111000" => data_out <= rom_array(7928);
		when "0001111011111001" => data_out <= rom_array(7929);
		when "0001111011111010" => data_out <= rom_array(7930);
		when "0001111011111011" => data_out <= rom_array(7931);
		when "0001111011111100" => data_out <= rom_array(7932);
		when "0001111011111101" => data_out <= rom_array(7933);
		when "0001111011111110" => data_out <= rom_array(7934);
		when "0001111011111111" => data_out <= rom_array(7935);
		when "0001111100000000" => data_out <= rom_array(7936);
		when "0001111100000001" => data_out <= rom_array(7937);
		when "0001111100000010" => data_out <= rom_array(7938);
		when "0001111100000011" => data_out <= rom_array(7939);
		when "0001111100000100" => data_out <= rom_array(7940);
		when "0001111100000101" => data_out <= rom_array(7941);
		when "0001111100000110" => data_out <= rom_array(7942);
		when "0001111100000111" => data_out <= rom_array(7943);
		when "0001111100001000" => data_out <= rom_array(7944);
		when "0001111100001001" => data_out <= rom_array(7945);
		when "0001111100001010" => data_out <= rom_array(7946);
		when "0001111100001011" => data_out <= rom_array(7947);
		when "0001111100001100" => data_out <= rom_array(7948);
		when "0001111100001101" => data_out <= rom_array(7949);
		when "0001111100001110" => data_out <= rom_array(7950);
		when "0001111100001111" => data_out <= rom_array(7951);
		when "0001111100010000" => data_out <= rom_array(7952);
		when "0001111100010001" => data_out <= rom_array(7953);
		when "0001111100010010" => data_out <= rom_array(7954);
		when "0001111100010011" => data_out <= rom_array(7955);
		when "0001111100010100" => data_out <= rom_array(7956);
		when "0001111100010101" => data_out <= rom_array(7957);
		when "0001111100010110" => data_out <= rom_array(7958);
		when "0001111100010111" => data_out <= rom_array(7959);
		when "0001111100011000" => data_out <= rom_array(7960);
		when "0001111100011001" => data_out <= rom_array(7961);
		when "0001111100011010" => data_out <= rom_array(7962);
		when "0001111100011011" => data_out <= rom_array(7963);
		when "0001111100011100" => data_out <= rom_array(7964);
		when "0001111100011101" => data_out <= rom_array(7965);
		when "0001111100011110" => data_out <= rom_array(7966);
		when "0001111100011111" => data_out <= rom_array(7967);
		when "0001111100100000" => data_out <= rom_array(7968);
		when "0001111100100001" => data_out <= rom_array(7969);
		when "0001111100100010" => data_out <= rom_array(7970);
		when "0001111100100011" => data_out <= rom_array(7971);
		when "0001111100100100" => data_out <= rom_array(7972);
		when "0001111100100101" => data_out <= rom_array(7973);
		when "0001111100100110" => data_out <= rom_array(7974);
		when "0001111100100111" => data_out <= rom_array(7975);
		when "0001111100101000" => data_out <= rom_array(7976);
		when "0001111100101001" => data_out <= rom_array(7977);
		when "0001111100101010" => data_out <= rom_array(7978);
		when "0001111100101011" => data_out <= rom_array(7979);
		when "0001111100101100" => data_out <= rom_array(7980);
		when "0001111100101101" => data_out <= rom_array(7981);
		when "0001111100101110" => data_out <= rom_array(7982);
		when "0001111100101111" => data_out <= rom_array(7983);
		when "0001111100110000" => data_out <= rom_array(7984);
		when "0001111100110001" => data_out <= rom_array(7985);
		when "0001111100110010" => data_out <= rom_array(7986);
		when "0001111100110011" => data_out <= rom_array(7987);
		when "0001111100110100" => data_out <= rom_array(7988);
		when "0001111100110101" => data_out <= rom_array(7989);
		when "0001111100110110" => data_out <= rom_array(7990);
		when "0001111100110111" => data_out <= rom_array(7991);
		when "0001111100111000" => data_out <= rom_array(7992);
		when "0001111100111001" => data_out <= rom_array(7993);
		when "0001111100111010" => data_out <= rom_array(7994);
		when "0001111100111011" => data_out <= rom_array(7995);
		when "0001111100111100" => data_out <= rom_array(7996);
		when "0001111100111101" => data_out <= rom_array(7997);
		when "0001111100111110" => data_out <= rom_array(7998);
		when "0001111100111111" => data_out <= rom_array(7999);
		when "0001111101000000" => data_out <= rom_array(8000);
		when "0001111101000001" => data_out <= rom_array(8001);
		when "0001111101000010" => data_out <= rom_array(8002);
		when "0001111101000011" => data_out <= rom_array(8003);
		when "0001111101000100" => data_out <= rom_array(8004);
		when "0001111101000101" => data_out <= rom_array(8005);
		when "0001111101000110" => data_out <= rom_array(8006);
		when "0001111101000111" => data_out <= rom_array(8007);
		when "0001111101001000" => data_out <= rom_array(8008);
		when "0001111101001001" => data_out <= rom_array(8009);
		when "0001111101001010" => data_out <= rom_array(8010);
		when "0001111101001011" => data_out <= rom_array(8011);
		when "0001111101001100" => data_out <= rom_array(8012);
		when "0001111101001101" => data_out <= rom_array(8013);
		when "0001111101001110" => data_out <= rom_array(8014);
		when "0001111101001111" => data_out <= rom_array(8015);
		when "0001111101010000" => data_out <= rom_array(8016);
		when "0001111101010001" => data_out <= rom_array(8017);
		when "0001111101010010" => data_out <= rom_array(8018);
		when "0001111101010011" => data_out <= rom_array(8019);
		when "0001111101010100" => data_out <= rom_array(8020);
		when "0001111101010101" => data_out <= rom_array(8021);
		when "0001111101010110" => data_out <= rom_array(8022);
		when "0001111101010111" => data_out <= rom_array(8023);
		when "0001111101011000" => data_out <= rom_array(8024);
		when "0001111101011001" => data_out <= rom_array(8025);
		when "0001111101011010" => data_out <= rom_array(8026);
		when "0001111101011011" => data_out <= rom_array(8027);
		when "0001111101011100" => data_out <= rom_array(8028);
		when "0001111101011101" => data_out <= rom_array(8029);
		when "0001111101011110" => data_out <= rom_array(8030);
		when "0001111101011111" => data_out <= rom_array(8031);
		when "0001111101100000" => data_out <= rom_array(8032);
		when "0001111101100001" => data_out <= rom_array(8033);
		when "0001111101100010" => data_out <= rom_array(8034);
		when "0001111101100011" => data_out <= rom_array(8035);
		when "0001111101100100" => data_out <= rom_array(8036);
		when "0001111101100101" => data_out <= rom_array(8037);
		when "0001111101100110" => data_out <= rom_array(8038);
		when "0001111101100111" => data_out <= rom_array(8039);
		when "0001111101101000" => data_out <= rom_array(8040);
		when "0001111101101001" => data_out <= rom_array(8041);
		when "0001111101101010" => data_out <= rom_array(8042);
		when "0001111101101011" => data_out <= rom_array(8043);
		when "0001111101101100" => data_out <= rom_array(8044);
		when "0001111101101101" => data_out <= rom_array(8045);
		when "0001111101101110" => data_out <= rom_array(8046);
		when "0001111101101111" => data_out <= rom_array(8047);
		when "0001111101110000" => data_out <= rom_array(8048);
		when "0001111101110001" => data_out <= rom_array(8049);
		when "0001111101110010" => data_out <= rom_array(8050);
		when "0001111101110011" => data_out <= rom_array(8051);
		when "0001111101110100" => data_out <= rom_array(8052);
		when "0001111101110101" => data_out <= rom_array(8053);
		when "0001111101110110" => data_out <= rom_array(8054);
		when "0001111101110111" => data_out <= rom_array(8055);
		when "0001111101111000" => data_out <= rom_array(8056);
		when "0001111101111001" => data_out <= rom_array(8057);
		when "0001111101111010" => data_out <= rom_array(8058);
		when "0001111101111011" => data_out <= rom_array(8059);
		when "0001111101111100" => data_out <= rom_array(8060);
		when "0001111101111101" => data_out <= rom_array(8061);
		when "0001111101111110" => data_out <= rom_array(8062);
		when "0001111101111111" => data_out <= rom_array(8063);
		when "0001111110000000" => data_out <= rom_array(8064);
		when "0001111110000001" => data_out <= rom_array(8065);
		when "0001111110000010" => data_out <= rom_array(8066);
		when "0001111110000011" => data_out <= rom_array(8067);
		when "0001111110000100" => data_out <= rom_array(8068);
		when "0001111110000101" => data_out <= rom_array(8069);
		when "0001111110000110" => data_out <= rom_array(8070);
		when "0001111110000111" => data_out <= rom_array(8071);
		when "0001111110001000" => data_out <= rom_array(8072);
		when "0001111110001001" => data_out <= rom_array(8073);
		when "0001111110001010" => data_out <= rom_array(8074);
		when "0001111110001011" => data_out <= rom_array(8075);
		when "0001111110001100" => data_out <= rom_array(8076);
		when "0001111110001101" => data_out <= rom_array(8077);
		when "0001111110001110" => data_out <= rom_array(8078);
		when "0001111110001111" => data_out <= rom_array(8079);
		when "0001111110010000" => data_out <= rom_array(8080);
		when "0001111110010001" => data_out <= rom_array(8081);
		when "0001111110010010" => data_out <= rom_array(8082);
		when "0001111110010011" => data_out <= rom_array(8083);
		when "0001111110010100" => data_out <= rom_array(8084);
		when "0001111110010101" => data_out <= rom_array(8085);
		when "0001111110010110" => data_out <= rom_array(8086);
		when "0001111110010111" => data_out <= rom_array(8087);
		when "0001111110011000" => data_out <= rom_array(8088);
		when "0001111110011001" => data_out <= rom_array(8089);
		when "0001111110011010" => data_out <= rom_array(8090);
		when "0001111110011011" => data_out <= rom_array(8091);
		when "0001111110011100" => data_out <= rom_array(8092);
		when "0001111110011101" => data_out <= rom_array(8093);
		when "0001111110011110" => data_out <= rom_array(8094);
		when "0001111110011111" => data_out <= rom_array(8095);
		when "0001111110100000" => data_out <= rom_array(8096);
		when "0001111110100001" => data_out <= rom_array(8097);
		when "0001111110100010" => data_out <= rom_array(8098);
		when "0001111110100011" => data_out <= rom_array(8099);
		when "0001111110100100" => data_out <= rom_array(8100);
		when "0001111110100101" => data_out <= rom_array(8101);
		when "0001111110100110" => data_out <= rom_array(8102);
		when "0001111110100111" => data_out <= rom_array(8103);
		when "0001111110101000" => data_out <= rom_array(8104);
		when "0001111110101001" => data_out <= rom_array(8105);
		when "0001111110101010" => data_out <= rom_array(8106);
		when "0001111110101011" => data_out <= rom_array(8107);
		when "0001111110101100" => data_out <= rom_array(8108);
		when "0001111110101101" => data_out <= rom_array(8109);
		when "0001111110101110" => data_out <= rom_array(8110);
		when "0001111110101111" => data_out <= rom_array(8111);
		when "0001111110110000" => data_out <= rom_array(8112);
		when "0001111110110001" => data_out <= rom_array(8113);
		when "0001111110110010" => data_out <= rom_array(8114);
		when "0001111110110011" => data_out <= rom_array(8115);
		when "0001111110110100" => data_out <= rom_array(8116);
		when "0001111110110101" => data_out <= rom_array(8117);
		when "0001111110110110" => data_out <= rom_array(8118);
		when "0001111110110111" => data_out <= rom_array(8119);
		when "0001111110111000" => data_out <= rom_array(8120);
		when "0001111110111001" => data_out <= rom_array(8121);
		when "0001111110111010" => data_out <= rom_array(8122);
		when "0001111110111011" => data_out <= rom_array(8123);
		when "0001111110111100" => data_out <= rom_array(8124);
		when "0001111110111101" => data_out <= rom_array(8125);
		when "0001111110111110" => data_out <= rom_array(8126);
		when "0001111110111111" => data_out <= rom_array(8127);
		when "0001111111000000" => data_out <= rom_array(8128);
		when "0001111111000001" => data_out <= rom_array(8129);
		when "0001111111000010" => data_out <= rom_array(8130);
		when "0001111111000011" => data_out <= rom_array(8131);
		when "0001111111000100" => data_out <= rom_array(8132);
		when "0001111111000101" => data_out <= rom_array(8133);
		when "0001111111000110" => data_out <= rom_array(8134);
		when "0001111111000111" => data_out <= rom_array(8135);
		when "0001111111001000" => data_out <= rom_array(8136);
		when "0001111111001001" => data_out <= rom_array(8137);
		when "0001111111001010" => data_out <= rom_array(8138);
		when "0001111111001011" => data_out <= rom_array(8139);
		when "0001111111001100" => data_out <= rom_array(8140);
		when "0001111111001101" => data_out <= rom_array(8141);
		when "0001111111001110" => data_out <= rom_array(8142);
		when "0001111111001111" => data_out <= rom_array(8143);
		when "0001111111010000" => data_out <= rom_array(8144);
		when "0001111111010001" => data_out <= rom_array(8145);
		when "0001111111010010" => data_out <= rom_array(8146);
		when "0001111111010011" => data_out <= rom_array(8147);
		when "0001111111010100" => data_out <= rom_array(8148);
		when "0001111111010101" => data_out <= rom_array(8149);
		when "0001111111010110" => data_out <= rom_array(8150);
		when "0001111111010111" => data_out <= rom_array(8151);
		when "0001111111011000" => data_out <= rom_array(8152);
		when "0001111111011001" => data_out <= rom_array(8153);
		when "0001111111011010" => data_out <= rom_array(8154);
		when "0001111111011011" => data_out <= rom_array(8155);
		when "0001111111011100" => data_out <= rom_array(8156);
		when "0001111111011101" => data_out <= rom_array(8157);
		when "0001111111011110" => data_out <= rom_array(8158);
		when "0001111111011111" => data_out <= rom_array(8159);
		when "0001111111100000" => data_out <= rom_array(8160);
		when "0001111111100001" => data_out <= rom_array(8161);
		when "0001111111100010" => data_out <= rom_array(8162);
		when "0001111111100011" => data_out <= rom_array(8163);
		when "0001111111100100" => data_out <= rom_array(8164);
		when "0001111111100101" => data_out <= rom_array(8165);
		when "0001111111100110" => data_out <= rom_array(8166);
		when "0001111111100111" => data_out <= rom_array(8167);
		when "0001111111101000" => data_out <= rom_array(8168);
		when "0001111111101001" => data_out <= rom_array(8169);
		when "0001111111101010" => data_out <= rom_array(8170);
		when "0001111111101011" => data_out <= rom_array(8171);
		when "0001111111101100" => data_out <= rom_array(8172);
		when "0001111111101101" => data_out <= rom_array(8173);
		when "0001111111101110" => data_out <= rom_array(8174);
		when "0001111111101111" => data_out <= rom_array(8175);
		when "0001111111110000" => data_out <= rom_array(8176);
		when "0001111111110001" => data_out <= rom_array(8177);
		when "0001111111110010" => data_out <= rom_array(8178);
		when "0001111111110011" => data_out <= rom_array(8179);
		when "0001111111110100" => data_out <= rom_array(8180);
		when "0001111111110101" => data_out <= rom_array(8181);
		when "0001111111110110" => data_out <= rom_array(8182);
		when "0001111111110111" => data_out <= rom_array(8183);
		when "0001111111111000" => data_out <= rom_array(8184);
		when "0001111111111001" => data_out <= rom_array(8185);
		when "0001111111111010" => data_out <= rom_array(8186);
		when "0001111111111011" => data_out <= rom_array(8187);
		when "0001111111111100" => data_out <= rom_array(8188);
		when "0001111111111101" => data_out <= rom_array(8189);
		when "0001111111111110" => data_out <= rom_array(8190);
		when "0001111111111111" => data_out <= rom_array(8191);
		when "0010000000000000" => data_out <= rom_array(8192);
		when "0010000000000001" => data_out <= rom_array(8193);
		when "0010000000000010" => data_out <= rom_array(8194);
		when "0010000000000011" => data_out <= rom_array(8195);
		when "0010000000000100" => data_out <= rom_array(8196);
		when "0010000000000101" => data_out <= rom_array(8197);
		when "0010000000000110" => data_out <= rom_array(8198);
		when "0010000000000111" => data_out <= rom_array(8199);
		when "0010000000001000" => data_out <= rom_array(8200);
		when "0010000000001001" => data_out <= rom_array(8201);
		when "0010000000001010" => data_out <= rom_array(8202);
		when "0010000000001011" => data_out <= rom_array(8203);
		when "0010000000001100" => data_out <= rom_array(8204);
		when "0010000000001101" => data_out <= rom_array(8205);
		when "0010000000001110" => data_out <= rom_array(8206);
		when "0010000000001111" => data_out <= rom_array(8207);
		when "0010000000010000" => data_out <= rom_array(8208);
		when "0010000000010001" => data_out <= rom_array(8209);
		when "0010000000010010" => data_out <= rom_array(8210);
		when "0010000000010011" => data_out <= rom_array(8211);
		when "0010000000010100" => data_out <= rom_array(8212);
		when "0010000000010101" => data_out <= rom_array(8213);
		when "0010000000010110" => data_out <= rom_array(8214);
		when "0010000000010111" => data_out <= rom_array(8215);
		when "0010000000011000" => data_out <= rom_array(8216);
		when "0010000000011001" => data_out <= rom_array(8217);
		when "0010000000011010" => data_out <= rom_array(8218);
		when "0010000000011011" => data_out <= rom_array(8219);
		when "0010000000011100" => data_out <= rom_array(8220);
		when "0010000000011101" => data_out <= rom_array(8221);
		when "0010000000011110" => data_out <= rom_array(8222);
		when "0010000000011111" => data_out <= rom_array(8223);
		when "0010000000100000" => data_out <= rom_array(8224);
		when "0010000000100001" => data_out <= rom_array(8225);
		when "0010000000100010" => data_out <= rom_array(8226);
		when "0010000000100011" => data_out <= rom_array(8227);
		when "0010000000100100" => data_out <= rom_array(8228);
		when "0010000000100101" => data_out <= rom_array(8229);
		when "0010000000100110" => data_out <= rom_array(8230);
		when "0010000000100111" => data_out <= rom_array(8231);
		when "0010000000101000" => data_out <= rom_array(8232);
		when "0010000000101001" => data_out <= rom_array(8233);
		when "0010000000101010" => data_out <= rom_array(8234);
		when "0010000000101011" => data_out <= rom_array(8235);
		when "0010000000101100" => data_out <= rom_array(8236);
		when "0010000000101101" => data_out <= rom_array(8237);
		when "0010000000101110" => data_out <= rom_array(8238);
		when "0010000000101111" => data_out <= rom_array(8239);
		when "0010000000110000" => data_out <= rom_array(8240);
		when "0010000000110001" => data_out <= rom_array(8241);
		when "0010000000110010" => data_out <= rom_array(8242);
		when "0010000000110011" => data_out <= rom_array(8243);
		when "0010000000110100" => data_out <= rom_array(8244);
		when "0010000000110101" => data_out <= rom_array(8245);
		when "0010000000110110" => data_out <= rom_array(8246);
		when "0010000000110111" => data_out <= rom_array(8247);
		when "0010000000111000" => data_out <= rom_array(8248);
		when "0010000000111001" => data_out <= rom_array(8249);
		when "0010000000111010" => data_out <= rom_array(8250);
		when "0010000000111011" => data_out <= rom_array(8251);
		when "0010000000111100" => data_out <= rom_array(8252);
		when "0010000000111101" => data_out <= rom_array(8253);
		when "0010000000111110" => data_out <= rom_array(8254);
		when "0010000000111111" => data_out <= rom_array(8255);
		when "0010000001000000" => data_out <= rom_array(8256);
		when "0010000001000001" => data_out <= rom_array(8257);
		when "0010000001000010" => data_out <= rom_array(8258);
		when "0010000001000011" => data_out <= rom_array(8259);
		when "0010000001000100" => data_out <= rom_array(8260);
		when "0010000001000101" => data_out <= rom_array(8261);
		when "0010000001000110" => data_out <= rom_array(8262);
		when "0010000001000111" => data_out <= rom_array(8263);
		when "0010000001001000" => data_out <= rom_array(8264);
		when "0010000001001001" => data_out <= rom_array(8265);
		when "0010000001001010" => data_out <= rom_array(8266);
		when "0010000001001011" => data_out <= rom_array(8267);
		when "0010000001001100" => data_out <= rom_array(8268);
		when "0010000001001101" => data_out <= rom_array(8269);
		when "0010000001001110" => data_out <= rom_array(8270);
		when "0010000001001111" => data_out <= rom_array(8271);
		when "0010000001010000" => data_out <= rom_array(8272);
		when "0010000001010001" => data_out <= rom_array(8273);
		when "0010000001010010" => data_out <= rom_array(8274);
		when "0010000001010011" => data_out <= rom_array(8275);
		when "0010000001010100" => data_out <= rom_array(8276);
		when "0010000001010101" => data_out <= rom_array(8277);
		when "0010000001010110" => data_out <= rom_array(8278);
		when "0010000001010111" => data_out <= rom_array(8279);
		when "0010000001011000" => data_out <= rom_array(8280);
		when "0010000001011001" => data_out <= rom_array(8281);
		when "0010000001011010" => data_out <= rom_array(8282);
		when "0010000001011011" => data_out <= rom_array(8283);
		when "0010000001011100" => data_out <= rom_array(8284);
		when "0010000001011101" => data_out <= rom_array(8285);
		when "0010000001011110" => data_out <= rom_array(8286);
		when "0010000001011111" => data_out <= rom_array(8287);
		when "0010000001100000" => data_out <= rom_array(8288);
		when "0010000001100001" => data_out <= rom_array(8289);
		when "0010000001100010" => data_out <= rom_array(8290);
		when "0010000001100011" => data_out <= rom_array(8291);
		when "0010000001100100" => data_out <= rom_array(8292);
		when "0010000001100101" => data_out <= rom_array(8293);
		when "0010000001100110" => data_out <= rom_array(8294);
		when "0010000001100111" => data_out <= rom_array(8295);
		when "0010000001101000" => data_out <= rom_array(8296);
		when "0010000001101001" => data_out <= rom_array(8297);
		when "0010000001101010" => data_out <= rom_array(8298);
		when "0010000001101011" => data_out <= rom_array(8299);
		when "0010000001101100" => data_out <= rom_array(8300);
		when "0010000001101101" => data_out <= rom_array(8301);
		when "0010000001101110" => data_out <= rom_array(8302);
		when "0010000001101111" => data_out <= rom_array(8303);
		when "0010000001110000" => data_out <= rom_array(8304);
		when "0010000001110001" => data_out <= rom_array(8305);
		when "0010000001110010" => data_out <= rom_array(8306);
		when "0010000001110011" => data_out <= rom_array(8307);
		when "0010000001110100" => data_out <= rom_array(8308);
		when "0010000001110101" => data_out <= rom_array(8309);
		when "0010000001110110" => data_out <= rom_array(8310);
		when "0010000001110111" => data_out <= rom_array(8311);
		when "0010000001111000" => data_out <= rom_array(8312);
		when "0010000001111001" => data_out <= rom_array(8313);
		when "0010000001111010" => data_out <= rom_array(8314);
		when "0010000001111011" => data_out <= rom_array(8315);
		when "0010000001111100" => data_out <= rom_array(8316);
		when "0010000001111101" => data_out <= rom_array(8317);
		when "0010000001111110" => data_out <= rom_array(8318);
		when "0010000001111111" => data_out <= rom_array(8319);
		when "0010000010000000" => data_out <= rom_array(8320);
		when "0010000010000001" => data_out <= rom_array(8321);
		when "0010000010000010" => data_out <= rom_array(8322);
		when "0010000010000011" => data_out <= rom_array(8323);
		when "0010000010000100" => data_out <= rom_array(8324);
		when "0010000010000101" => data_out <= rom_array(8325);
		when "0010000010000110" => data_out <= rom_array(8326);
		when "0010000010000111" => data_out <= rom_array(8327);
		when "0010000010001000" => data_out <= rom_array(8328);
		when "0010000010001001" => data_out <= rom_array(8329);
		when "0010000010001010" => data_out <= rom_array(8330);
		when "0010000010001011" => data_out <= rom_array(8331);
		when "0010000010001100" => data_out <= rom_array(8332);
		when "0010000010001101" => data_out <= rom_array(8333);
		when "0010000010001110" => data_out <= rom_array(8334);
		when "0010000010001111" => data_out <= rom_array(8335);
		when "0010000010010000" => data_out <= rom_array(8336);
		when "0010000010010001" => data_out <= rom_array(8337);
		when "0010000010010010" => data_out <= rom_array(8338);
		when "0010000010010011" => data_out <= rom_array(8339);
		when "0010000010010100" => data_out <= rom_array(8340);
		when "0010000010010101" => data_out <= rom_array(8341);
		when "0010000010010110" => data_out <= rom_array(8342);
		when "0010000010010111" => data_out <= rom_array(8343);
		when "0010000010011000" => data_out <= rom_array(8344);
		when "0010000010011001" => data_out <= rom_array(8345);
		when "0010000010011010" => data_out <= rom_array(8346);
		when "0010000010011011" => data_out <= rom_array(8347);
		when "0010000010011100" => data_out <= rom_array(8348);
		when "0010000010011101" => data_out <= rom_array(8349);
		when "0010000010011110" => data_out <= rom_array(8350);
		when "0010000010011111" => data_out <= rom_array(8351);
		when "0010000010100000" => data_out <= rom_array(8352);
		when "0010000010100001" => data_out <= rom_array(8353);
		when "0010000010100010" => data_out <= rom_array(8354);
		when "0010000010100011" => data_out <= rom_array(8355);
		when "0010000010100100" => data_out <= rom_array(8356);
		when "0010000010100101" => data_out <= rom_array(8357);
		when "0010000010100110" => data_out <= rom_array(8358);
		when "0010000010100111" => data_out <= rom_array(8359);
		when "0010000010101000" => data_out <= rom_array(8360);
		when "0010000010101001" => data_out <= rom_array(8361);
		when "0010000010101010" => data_out <= rom_array(8362);
		when "0010000010101011" => data_out <= rom_array(8363);
		when "0010000010101100" => data_out <= rom_array(8364);
		when "0010000010101101" => data_out <= rom_array(8365);
		when "0010000010101110" => data_out <= rom_array(8366);
		when "0010000010101111" => data_out <= rom_array(8367);
		when "0010000010110000" => data_out <= rom_array(8368);
		when "0010000010110001" => data_out <= rom_array(8369);
		when "0010000010110010" => data_out <= rom_array(8370);
		when "0010000010110011" => data_out <= rom_array(8371);
		when "0010000010110100" => data_out <= rom_array(8372);
		when "0010000010110101" => data_out <= rom_array(8373);
		when "0010000010110110" => data_out <= rom_array(8374);
		when "0010000010110111" => data_out <= rom_array(8375);
		when "0010000010111000" => data_out <= rom_array(8376);
		when "0010000010111001" => data_out <= rom_array(8377);
		when "0010000010111010" => data_out <= rom_array(8378);
		when "0010000010111011" => data_out <= rom_array(8379);
		when "0010000010111100" => data_out <= rom_array(8380);
		when "0010000010111101" => data_out <= rom_array(8381);
		when "0010000010111110" => data_out <= rom_array(8382);
		when "0010000010111111" => data_out <= rom_array(8383);
		when "0010000011000000" => data_out <= rom_array(8384);
		when "0010000011000001" => data_out <= rom_array(8385);
		when "0010000011000010" => data_out <= rom_array(8386);
		when "0010000011000011" => data_out <= rom_array(8387);
		when "0010000011000100" => data_out <= rom_array(8388);
		when "0010000011000101" => data_out <= rom_array(8389);
		when "0010000011000110" => data_out <= rom_array(8390);
		when "0010000011000111" => data_out <= rom_array(8391);
		when "0010000011001000" => data_out <= rom_array(8392);
		when "0010000011001001" => data_out <= rom_array(8393);
		when "0010000011001010" => data_out <= rom_array(8394);
		when "0010000011001011" => data_out <= rom_array(8395);
		when "0010000011001100" => data_out <= rom_array(8396);
		when "0010000011001101" => data_out <= rom_array(8397);
		when "0010000011001110" => data_out <= rom_array(8398);
		when "0010000011001111" => data_out <= rom_array(8399);
		when "0010000011010000" => data_out <= rom_array(8400);
		when "0010000011010001" => data_out <= rom_array(8401);
		when "0010000011010010" => data_out <= rom_array(8402);
		when "0010000011010011" => data_out <= rom_array(8403);
		when "0010000011010100" => data_out <= rom_array(8404);
		when "0010000011010101" => data_out <= rom_array(8405);
		when "0010000011010110" => data_out <= rom_array(8406);
		when "0010000011010111" => data_out <= rom_array(8407);
		when "0010000011011000" => data_out <= rom_array(8408);
		when "0010000011011001" => data_out <= rom_array(8409);
		when "0010000011011010" => data_out <= rom_array(8410);
		when "0010000011011011" => data_out <= rom_array(8411);
		when "0010000011011100" => data_out <= rom_array(8412);
		when "0010000011011101" => data_out <= rom_array(8413);
		when "0010000011011110" => data_out <= rom_array(8414);
		when "0010000011011111" => data_out <= rom_array(8415);
		when "0010000011100000" => data_out <= rom_array(8416);
		when "0010000011100001" => data_out <= rom_array(8417);
		when "0010000011100010" => data_out <= rom_array(8418);
		when "0010000011100011" => data_out <= rom_array(8419);
		when "0010000011100100" => data_out <= rom_array(8420);
		when "0010000011100101" => data_out <= rom_array(8421);
		when "0010000011100110" => data_out <= rom_array(8422);
		when "0010000011100111" => data_out <= rom_array(8423);
		when "0010000011101000" => data_out <= rom_array(8424);
		when "0010000011101001" => data_out <= rom_array(8425);
		when "0010000011101010" => data_out <= rom_array(8426);
		when "0010000011101011" => data_out <= rom_array(8427);
		when "0010000011101100" => data_out <= rom_array(8428);
		when "0010000011101101" => data_out <= rom_array(8429);
		when "0010000011101110" => data_out <= rom_array(8430);
		when "0010000011101111" => data_out <= rom_array(8431);
		when "0010000011110000" => data_out <= rom_array(8432);
		when "0010000011110001" => data_out <= rom_array(8433);
		when "0010000011110010" => data_out <= rom_array(8434);
		when "0010000011110011" => data_out <= rom_array(8435);
		when "0010000011110100" => data_out <= rom_array(8436);
		when "0010000011110101" => data_out <= rom_array(8437);
		when "0010000011110110" => data_out <= rom_array(8438);
		when "0010000011110111" => data_out <= rom_array(8439);
		when "0010000011111000" => data_out <= rom_array(8440);
		when "0010000011111001" => data_out <= rom_array(8441);
		when "0010000011111010" => data_out <= rom_array(8442);
		when "0010000011111011" => data_out <= rom_array(8443);
		when "0010000011111100" => data_out <= rom_array(8444);
		when "0010000011111101" => data_out <= rom_array(8445);
		when "0010000011111110" => data_out <= rom_array(8446);
		when "0010000011111111" => data_out <= rom_array(8447);
		when "0010000100000000" => data_out <= rom_array(8448);
		when "0010000100000001" => data_out <= rom_array(8449);
		when "0010000100000010" => data_out <= rom_array(8450);
		when "0010000100000011" => data_out <= rom_array(8451);
		when "0010000100000100" => data_out <= rom_array(8452);
		when "0010000100000101" => data_out <= rom_array(8453);
		when "0010000100000110" => data_out <= rom_array(8454);
		when "0010000100000111" => data_out <= rom_array(8455);
		when "0010000100001000" => data_out <= rom_array(8456);
		when "0010000100001001" => data_out <= rom_array(8457);
		when "0010000100001010" => data_out <= rom_array(8458);
		when "0010000100001011" => data_out <= rom_array(8459);
		when "0010000100001100" => data_out <= rom_array(8460);
		when "0010000100001101" => data_out <= rom_array(8461);
		when "0010000100001110" => data_out <= rom_array(8462);
		when "0010000100001111" => data_out <= rom_array(8463);
		when "0010000100010000" => data_out <= rom_array(8464);
		when "0010000100010001" => data_out <= rom_array(8465);
		when "0010000100010010" => data_out <= rom_array(8466);
		when "0010000100010011" => data_out <= rom_array(8467);
		when "0010000100010100" => data_out <= rom_array(8468);
		when "0010000100010101" => data_out <= rom_array(8469);
		when "0010000100010110" => data_out <= rom_array(8470);
		when "0010000100010111" => data_out <= rom_array(8471);
		when "0010000100011000" => data_out <= rom_array(8472);
		when "0010000100011001" => data_out <= rom_array(8473);
		when "0010000100011010" => data_out <= rom_array(8474);
		when "0010000100011011" => data_out <= rom_array(8475);
		when "0010000100011100" => data_out <= rom_array(8476);
		when "0010000100011101" => data_out <= rom_array(8477);
		when "0010000100011110" => data_out <= rom_array(8478);
		when "0010000100011111" => data_out <= rom_array(8479);
		when "0010000100100000" => data_out <= rom_array(8480);
		when "0010000100100001" => data_out <= rom_array(8481);
		when "0010000100100010" => data_out <= rom_array(8482);
		when "0010000100100011" => data_out <= rom_array(8483);
		when "0010000100100100" => data_out <= rom_array(8484);
		when "0010000100100101" => data_out <= rom_array(8485);
		when "0010000100100110" => data_out <= rom_array(8486);
		when "0010000100100111" => data_out <= rom_array(8487);
		when "0010000100101000" => data_out <= rom_array(8488);
		when "0010000100101001" => data_out <= rom_array(8489);
		when "0010000100101010" => data_out <= rom_array(8490);
		when "0010000100101011" => data_out <= rom_array(8491);
		when "0010000100101100" => data_out <= rom_array(8492);
		when "0010000100101101" => data_out <= rom_array(8493);
		when "0010000100101110" => data_out <= rom_array(8494);
		when "0010000100101111" => data_out <= rom_array(8495);
		when "0010000100110000" => data_out <= rom_array(8496);
		when "0010000100110001" => data_out <= rom_array(8497);
		when "0010000100110010" => data_out <= rom_array(8498);
		when "0010000100110011" => data_out <= rom_array(8499);
		when "0010000100110100" => data_out <= rom_array(8500);
		when "0010000100110101" => data_out <= rom_array(8501);
		when "0010000100110110" => data_out <= rom_array(8502);
		when "0010000100110111" => data_out <= rom_array(8503);
		when "0010000100111000" => data_out <= rom_array(8504);
		when "0010000100111001" => data_out <= rom_array(8505);
		when "0010000100111010" => data_out <= rom_array(8506);
		when "0010000100111011" => data_out <= rom_array(8507);
		when "0010000100111100" => data_out <= rom_array(8508);
		when "0010000100111101" => data_out <= rom_array(8509);
		when "0010000100111110" => data_out <= rom_array(8510);
		when "0010000100111111" => data_out <= rom_array(8511);
		when "0010000101000000" => data_out <= rom_array(8512);
		when "0010000101000001" => data_out <= rom_array(8513);
		when "0010000101000010" => data_out <= rom_array(8514);
		when "0010000101000011" => data_out <= rom_array(8515);
		when "0010000101000100" => data_out <= rom_array(8516);
		when "0010000101000101" => data_out <= rom_array(8517);
		when "0010000101000110" => data_out <= rom_array(8518);
		when "0010000101000111" => data_out <= rom_array(8519);
		when "0010000101001000" => data_out <= rom_array(8520);
		when "0010000101001001" => data_out <= rom_array(8521);
		when "0010000101001010" => data_out <= rom_array(8522);
		when "0010000101001011" => data_out <= rom_array(8523);
		when "0010000101001100" => data_out <= rom_array(8524);
		when "0010000101001101" => data_out <= rom_array(8525);
		when "0010000101001110" => data_out <= rom_array(8526);
		when "0010000101001111" => data_out <= rom_array(8527);
		when "0010000101010000" => data_out <= rom_array(8528);
		when "0010000101010001" => data_out <= rom_array(8529);
		when "0010000101010010" => data_out <= rom_array(8530);
		when "0010000101010011" => data_out <= rom_array(8531);
		when "0010000101010100" => data_out <= rom_array(8532);
		when "0010000101010101" => data_out <= rom_array(8533);
		when "0010000101010110" => data_out <= rom_array(8534);
		when "0010000101010111" => data_out <= rom_array(8535);
		when "0010000101011000" => data_out <= rom_array(8536);
		when "0010000101011001" => data_out <= rom_array(8537);
		when "0010000101011010" => data_out <= rom_array(8538);
		when "0010000101011011" => data_out <= rom_array(8539);
		when "0010000101011100" => data_out <= rom_array(8540);
		when "0010000101011101" => data_out <= rom_array(8541);
		when "0010000101011110" => data_out <= rom_array(8542);
		when "0010000101011111" => data_out <= rom_array(8543);
		when "0010000101100000" => data_out <= rom_array(8544);
		when "0010000101100001" => data_out <= rom_array(8545);
		when "0010000101100010" => data_out <= rom_array(8546);
		when "0010000101100011" => data_out <= rom_array(8547);
		when "0010000101100100" => data_out <= rom_array(8548);
		when "0010000101100101" => data_out <= rom_array(8549);
		when "0010000101100110" => data_out <= rom_array(8550);
		when "0010000101100111" => data_out <= rom_array(8551);
		when "0010000101101000" => data_out <= rom_array(8552);
		when "0010000101101001" => data_out <= rom_array(8553);
		when "0010000101101010" => data_out <= rom_array(8554);
		when "0010000101101011" => data_out <= rom_array(8555);
		when "0010000101101100" => data_out <= rom_array(8556);
		when "0010000101101101" => data_out <= rom_array(8557);
		when "0010000101101110" => data_out <= rom_array(8558);
		when "0010000101101111" => data_out <= rom_array(8559);
		when "0010000101110000" => data_out <= rom_array(8560);
		when "0010000101110001" => data_out <= rom_array(8561);
		when "0010000101110010" => data_out <= rom_array(8562);
		when "0010000101110011" => data_out <= rom_array(8563);
		when "0010000101110100" => data_out <= rom_array(8564);
		when "0010000101110101" => data_out <= rom_array(8565);
		when "0010000101110110" => data_out <= rom_array(8566);
		when "0010000101110111" => data_out <= rom_array(8567);
		when "0010000101111000" => data_out <= rom_array(8568);
		when "0010000101111001" => data_out <= rom_array(8569);
		when "0010000101111010" => data_out <= rom_array(8570);
		when "0010000101111011" => data_out <= rom_array(8571);
		when "0010000101111100" => data_out <= rom_array(8572);
		when "0010000101111101" => data_out <= rom_array(8573);
		when "0010000101111110" => data_out <= rom_array(8574);
		when "0010000101111111" => data_out <= rom_array(8575);
		when "0010000110000000" => data_out <= rom_array(8576);
		when "0010000110000001" => data_out <= rom_array(8577);
		when "0010000110000010" => data_out <= rom_array(8578);
		when "0010000110000011" => data_out <= rom_array(8579);
		when "0010000110000100" => data_out <= rom_array(8580);
		when "0010000110000101" => data_out <= rom_array(8581);
		when "0010000110000110" => data_out <= rom_array(8582);
		when "0010000110000111" => data_out <= rom_array(8583);
		when "0010000110001000" => data_out <= rom_array(8584);
		when "0010000110001001" => data_out <= rom_array(8585);
		when "0010000110001010" => data_out <= rom_array(8586);
		when "0010000110001011" => data_out <= rom_array(8587);
		when "0010000110001100" => data_out <= rom_array(8588);
		when "0010000110001101" => data_out <= rom_array(8589);
		when "0010000110001110" => data_out <= rom_array(8590);
		when "0010000110001111" => data_out <= rom_array(8591);
		when "0010000110010000" => data_out <= rom_array(8592);
		when "0010000110010001" => data_out <= rom_array(8593);
		when "0010000110010010" => data_out <= rom_array(8594);
		when "0010000110010011" => data_out <= rom_array(8595);
		when "0010000110010100" => data_out <= rom_array(8596);
		when "0010000110010101" => data_out <= rom_array(8597);
		when "0010000110010110" => data_out <= rom_array(8598);
		when "0010000110010111" => data_out <= rom_array(8599);
		when "0010000110011000" => data_out <= rom_array(8600);
		when "0010000110011001" => data_out <= rom_array(8601);
		when "0010000110011010" => data_out <= rom_array(8602);
		when "0010000110011011" => data_out <= rom_array(8603);
		when "0010000110011100" => data_out <= rom_array(8604);
		when "0010000110011101" => data_out <= rom_array(8605);
		when "0010000110011110" => data_out <= rom_array(8606);
		when "0010000110011111" => data_out <= rom_array(8607);
		when "0010000110100000" => data_out <= rom_array(8608);
		when "0010000110100001" => data_out <= rom_array(8609);
		when "0010000110100010" => data_out <= rom_array(8610);
		when "0010000110100011" => data_out <= rom_array(8611);
		when "0010000110100100" => data_out <= rom_array(8612);
		when "0010000110100101" => data_out <= rom_array(8613);
		when "0010000110100110" => data_out <= rom_array(8614);
		when "0010000110100111" => data_out <= rom_array(8615);
		when "0010000110101000" => data_out <= rom_array(8616);
		when "0010000110101001" => data_out <= rom_array(8617);
		when "0010000110101010" => data_out <= rom_array(8618);
		when "0010000110101011" => data_out <= rom_array(8619);
		when "0010000110101100" => data_out <= rom_array(8620);
		when "0010000110101101" => data_out <= rom_array(8621);
		when "0010000110101110" => data_out <= rom_array(8622);
		when "0010000110101111" => data_out <= rom_array(8623);
		when "0010000110110000" => data_out <= rom_array(8624);
		when "0010000110110001" => data_out <= rom_array(8625);
		when "0010000110110010" => data_out <= rom_array(8626);
		when "0010000110110011" => data_out <= rom_array(8627);
		when "0010000110110100" => data_out <= rom_array(8628);
		when "0010000110110101" => data_out <= rom_array(8629);
		when "0010000110110110" => data_out <= rom_array(8630);
		when "0010000110110111" => data_out <= rom_array(8631);
		when "0010000110111000" => data_out <= rom_array(8632);
		when "0010000110111001" => data_out <= rom_array(8633);
		when "0010000110111010" => data_out <= rom_array(8634);
		when "0010000110111011" => data_out <= rom_array(8635);
		when "0010000110111100" => data_out <= rom_array(8636);
		when "0010000110111101" => data_out <= rom_array(8637);
		when "0010000110111110" => data_out <= rom_array(8638);
		when "0010000110111111" => data_out <= rom_array(8639);
		when "0010000111000000" => data_out <= rom_array(8640);
		when "0010000111000001" => data_out <= rom_array(8641);
		when "0010000111000010" => data_out <= rom_array(8642);
		when "0010000111000011" => data_out <= rom_array(8643);
		when "0010000111000100" => data_out <= rom_array(8644);
		when "0010000111000101" => data_out <= rom_array(8645);
		when "0010000111000110" => data_out <= rom_array(8646);
		when "0010000111000111" => data_out <= rom_array(8647);
		when "0010000111001000" => data_out <= rom_array(8648);
		when "0010000111001001" => data_out <= rom_array(8649);
		when "0010000111001010" => data_out <= rom_array(8650);
		when "0010000111001011" => data_out <= rom_array(8651);
		when "0010000111001100" => data_out <= rom_array(8652);
		when "0010000111001101" => data_out <= rom_array(8653);
		when "0010000111001110" => data_out <= rom_array(8654);
		when "0010000111001111" => data_out <= rom_array(8655);
		when "0010000111010000" => data_out <= rom_array(8656);
		when "0010000111010001" => data_out <= rom_array(8657);
		when "0010000111010010" => data_out <= rom_array(8658);
		when "0010000111010011" => data_out <= rom_array(8659);
		when "0010000111010100" => data_out <= rom_array(8660);
		when "0010000111010101" => data_out <= rom_array(8661);
		when "0010000111010110" => data_out <= rom_array(8662);
		when "0010000111010111" => data_out <= rom_array(8663);
		when "0010000111011000" => data_out <= rom_array(8664);
		when "0010000111011001" => data_out <= rom_array(8665);
		when "0010000111011010" => data_out <= rom_array(8666);
		when "0010000111011011" => data_out <= rom_array(8667);
		when "0010000111011100" => data_out <= rom_array(8668);
		when "0010000111011101" => data_out <= rom_array(8669);
		when "0010000111011110" => data_out <= rom_array(8670);
		when "0010000111011111" => data_out <= rom_array(8671);
		when "0010000111100000" => data_out <= rom_array(8672);
		when "0010000111100001" => data_out <= rom_array(8673);
		when "0010000111100010" => data_out <= rom_array(8674);
		when "0010000111100011" => data_out <= rom_array(8675);
		when "0010000111100100" => data_out <= rom_array(8676);
		when "0010000111100101" => data_out <= rom_array(8677);
		when "0010000111100110" => data_out <= rom_array(8678);
		when "0010000111100111" => data_out <= rom_array(8679);
		when "0010000111101000" => data_out <= rom_array(8680);
		when "0010000111101001" => data_out <= rom_array(8681);
		when "0010000111101010" => data_out <= rom_array(8682);
		when "0010000111101011" => data_out <= rom_array(8683);
		when "0010000111101100" => data_out <= rom_array(8684);
		when "0010000111101101" => data_out <= rom_array(8685);
		when "0010000111101110" => data_out <= rom_array(8686);
		when "0010000111101111" => data_out <= rom_array(8687);
		when "0010000111110000" => data_out <= rom_array(8688);
		when "0010000111110001" => data_out <= rom_array(8689);
		when "0010000111110010" => data_out <= rom_array(8690);
		when "0010000111110011" => data_out <= rom_array(8691);
		when "0010000111110100" => data_out <= rom_array(8692);
		when "0010000111110101" => data_out <= rom_array(8693);
		when "0010000111110110" => data_out <= rom_array(8694);
		when "0010000111110111" => data_out <= rom_array(8695);
		when "0010000111111000" => data_out <= rom_array(8696);
		when "0010000111111001" => data_out <= rom_array(8697);
		when "0010000111111010" => data_out <= rom_array(8698);
		when "0010000111111011" => data_out <= rom_array(8699);
		when "0010000111111100" => data_out <= rom_array(8700);
		when "0010000111111101" => data_out <= rom_array(8701);
		when "0010000111111110" => data_out <= rom_array(8702);
		when "0010000111111111" => data_out <= rom_array(8703);
		when "0010001000000000" => data_out <= rom_array(8704);
		when "0010001000000001" => data_out <= rom_array(8705);
		when "0010001000000010" => data_out <= rom_array(8706);
		when "0010001000000011" => data_out <= rom_array(8707);
		when "0010001000000100" => data_out <= rom_array(8708);
		when "0010001000000101" => data_out <= rom_array(8709);
		when "0010001000000110" => data_out <= rom_array(8710);
		when "0010001000000111" => data_out <= rom_array(8711);
		when "0010001000001000" => data_out <= rom_array(8712);
		when "0010001000001001" => data_out <= rom_array(8713);
		when "0010001000001010" => data_out <= rom_array(8714);
		when "0010001000001011" => data_out <= rom_array(8715);
		when "0010001000001100" => data_out <= rom_array(8716);
		when "0010001000001101" => data_out <= rom_array(8717);
		when "0010001000001110" => data_out <= rom_array(8718);
		when "0010001000001111" => data_out <= rom_array(8719);
		when "0010001000010000" => data_out <= rom_array(8720);
		when "0010001000010001" => data_out <= rom_array(8721);
		when "0010001000010010" => data_out <= rom_array(8722);
		when "0010001000010011" => data_out <= rom_array(8723);
		when "0010001000010100" => data_out <= rom_array(8724);
		when "0010001000010101" => data_out <= rom_array(8725);
		when "0010001000010110" => data_out <= rom_array(8726);
		when "0010001000010111" => data_out <= rom_array(8727);
		when "0010001000011000" => data_out <= rom_array(8728);
		when "0010001000011001" => data_out <= rom_array(8729);
		when "0010001000011010" => data_out <= rom_array(8730);
		when "0010001000011011" => data_out <= rom_array(8731);
		when "0010001000011100" => data_out <= rom_array(8732);
		when "0010001000011101" => data_out <= rom_array(8733);
		when "0010001000011110" => data_out <= rom_array(8734);
		when "0010001000011111" => data_out <= rom_array(8735);
		when "0010001000100000" => data_out <= rom_array(8736);
		when "0010001000100001" => data_out <= rom_array(8737);
		when "0010001000100010" => data_out <= rom_array(8738);
		when "0010001000100011" => data_out <= rom_array(8739);
		when "0010001000100100" => data_out <= rom_array(8740);
		when "0010001000100101" => data_out <= rom_array(8741);
		when "0010001000100110" => data_out <= rom_array(8742);
		when "0010001000100111" => data_out <= rom_array(8743);
		when "0010001000101000" => data_out <= rom_array(8744);
		when "0010001000101001" => data_out <= rom_array(8745);
		when "0010001000101010" => data_out <= rom_array(8746);
		when "0010001000101011" => data_out <= rom_array(8747);
		when "0010001000101100" => data_out <= rom_array(8748);
		when "0010001000101101" => data_out <= rom_array(8749);
		when "0010001000101110" => data_out <= rom_array(8750);
		when "0010001000101111" => data_out <= rom_array(8751);
		when "0010001000110000" => data_out <= rom_array(8752);
		when "0010001000110001" => data_out <= rom_array(8753);
		when "0010001000110010" => data_out <= rom_array(8754);
		when "0010001000110011" => data_out <= rom_array(8755);
		when "0010001000110100" => data_out <= rom_array(8756);
		when "0010001000110101" => data_out <= rom_array(8757);
		when "0010001000110110" => data_out <= rom_array(8758);
		when "0010001000110111" => data_out <= rom_array(8759);
		when "0010001000111000" => data_out <= rom_array(8760);
		when "0010001000111001" => data_out <= rom_array(8761);
		when "0010001000111010" => data_out <= rom_array(8762);
		when "0010001000111011" => data_out <= rom_array(8763);
		when "0010001000111100" => data_out <= rom_array(8764);
		when "0010001000111101" => data_out <= rom_array(8765);
		when "0010001000111110" => data_out <= rom_array(8766);
		when "0010001000111111" => data_out <= rom_array(8767);
		when "0010001001000000" => data_out <= rom_array(8768);
		when "0010001001000001" => data_out <= rom_array(8769);
		when "0010001001000010" => data_out <= rom_array(8770);
		when "0010001001000011" => data_out <= rom_array(8771);
		when "0010001001000100" => data_out <= rom_array(8772);
		when "0010001001000101" => data_out <= rom_array(8773);
		when "0010001001000110" => data_out <= rom_array(8774);
		when "0010001001000111" => data_out <= rom_array(8775);
		when "0010001001001000" => data_out <= rom_array(8776);
		when "0010001001001001" => data_out <= rom_array(8777);
		when "0010001001001010" => data_out <= rom_array(8778);
		when "0010001001001011" => data_out <= rom_array(8779);
		when "0010001001001100" => data_out <= rom_array(8780);
		when "0010001001001101" => data_out <= rom_array(8781);
		when "0010001001001110" => data_out <= rom_array(8782);
		when "0010001001001111" => data_out <= rom_array(8783);
		when "0010001001010000" => data_out <= rom_array(8784);
		when "0010001001010001" => data_out <= rom_array(8785);
		when "0010001001010010" => data_out <= rom_array(8786);
		when "0010001001010011" => data_out <= rom_array(8787);
		when "0010001001010100" => data_out <= rom_array(8788);
		when "0010001001010101" => data_out <= rom_array(8789);
		when "0010001001010110" => data_out <= rom_array(8790);
		when "0010001001010111" => data_out <= rom_array(8791);
		when "0010001001011000" => data_out <= rom_array(8792);
		when "0010001001011001" => data_out <= rom_array(8793);
		when "0010001001011010" => data_out <= rom_array(8794);
		when "0010001001011011" => data_out <= rom_array(8795);
		when "0010001001011100" => data_out <= rom_array(8796);
		when "0010001001011101" => data_out <= rom_array(8797);
		when "0010001001011110" => data_out <= rom_array(8798);
		when "0010001001011111" => data_out <= rom_array(8799);
		when "0010001001100000" => data_out <= rom_array(8800);
		when "0010001001100001" => data_out <= rom_array(8801);
		when "0010001001100010" => data_out <= rom_array(8802);
		when "0010001001100011" => data_out <= rom_array(8803);
		when "0010001001100100" => data_out <= rom_array(8804);
		when "0010001001100101" => data_out <= rom_array(8805);
		when "0010001001100110" => data_out <= rom_array(8806);
		when "0010001001100111" => data_out <= rom_array(8807);
		when "0010001001101000" => data_out <= rom_array(8808);
		when "0010001001101001" => data_out <= rom_array(8809);
		when "0010001001101010" => data_out <= rom_array(8810);
		when "0010001001101011" => data_out <= rom_array(8811);
		when "0010001001101100" => data_out <= rom_array(8812);
		when "0010001001101101" => data_out <= rom_array(8813);
		when "0010001001101110" => data_out <= rom_array(8814);
		when "0010001001101111" => data_out <= rom_array(8815);
		when "0010001001110000" => data_out <= rom_array(8816);
		when "0010001001110001" => data_out <= rom_array(8817);
		when "0010001001110010" => data_out <= rom_array(8818);
		when "0010001001110011" => data_out <= rom_array(8819);
		when "0010001001110100" => data_out <= rom_array(8820);
		when "0010001001110101" => data_out <= rom_array(8821);
		when "0010001001110110" => data_out <= rom_array(8822);
		when "0010001001110111" => data_out <= rom_array(8823);
		when "0010001001111000" => data_out <= rom_array(8824);
		when "0010001001111001" => data_out <= rom_array(8825);
		when "0010001001111010" => data_out <= rom_array(8826);
		when "0010001001111011" => data_out <= rom_array(8827);
		when "0010001001111100" => data_out <= rom_array(8828);
		when "0010001001111101" => data_out <= rom_array(8829);
		when "0010001001111110" => data_out <= rom_array(8830);
		when "0010001001111111" => data_out <= rom_array(8831);
		when "0010001010000000" => data_out <= rom_array(8832);
		when "0010001010000001" => data_out <= rom_array(8833);
		when "0010001010000010" => data_out <= rom_array(8834);
		when "0010001010000011" => data_out <= rom_array(8835);
		when "0010001010000100" => data_out <= rom_array(8836);
		when "0010001010000101" => data_out <= rom_array(8837);
		when "0010001010000110" => data_out <= rom_array(8838);
		when "0010001010000111" => data_out <= rom_array(8839);
		when "0010001010001000" => data_out <= rom_array(8840);
		when "0010001010001001" => data_out <= rom_array(8841);
		when "0010001010001010" => data_out <= rom_array(8842);
		when "0010001010001011" => data_out <= rom_array(8843);
		when "0010001010001100" => data_out <= rom_array(8844);
		when "0010001010001101" => data_out <= rom_array(8845);
		when "0010001010001110" => data_out <= rom_array(8846);
		when "0010001010001111" => data_out <= rom_array(8847);
		when "0010001010010000" => data_out <= rom_array(8848);
		when "0010001010010001" => data_out <= rom_array(8849);
		when "0010001010010010" => data_out <= rom_array(8850);
		when "0010001010010011" => data_out <= rom_array(8851);
		when "0010001010010100" => data_out <= rom_array(8852);
		when "0010001010010101" => data_out <= rom_array(8853);
		when "0010001010010110" => data_out <= rom_array(8854);
		when "0010001010010111" => data_out <= rom_array(8855);
		when "0010001010011000" => data_out <= rom_array(8856);
		when "0010001010011001" => data_out <= rom_array(8857);
		when "0010001010011010" => data_out <= rom_array(8858);
		when "0010001010011011" => data_out <= rom_array(8859);
		when "0010001010011100" => data_out <= rom_array(8860);
		when "0010001010011101" => data_out <= rom_array(8861);
		when "0010001010011110" => data_out <= rom_array(8862);
		when "0010001010011111" => data_out <= rom_array(8863);
		when "0010001010100000" => data_out <= rom_array(8864);
		when "0010001010100001" => data_out <= rom_array(8865);
		when "0010001010100010" => data_out <= rom_array(8866);
		when "0010001010100011" => data_out <= rom_array(8867);
		when "0010001010100100" => data_out <= rom_array(8868);
		when "0010001010100101" => data_out <= rom_array(8869);
		when "0010001010100110" => data_out <= rom_array(8870);
		when "0010001010100111" => data_out <= rom_array(8871);
		when "0010001010101000" => data_out <= rom_array(8872);
		when "0010001010101001" => data_out <= rom_array(8873);
		when "0010001010101010" => data_out <= rom_array(8874);
		when "0010001010101011" => data_out <= rom_array(8875);
		when "0010001010101100" => data_out <= rom_array(8876);
		when "0010001010101101" => data_out <= rom_array(8877);
		when "0010001010101110" => data_out <= rom_array(8878);
		when "0010001010101111" => data_out <= rom_array(8879);
		when "0010001010110000" => data_out <= rom_array(8880);
		when "0010001010110001" => data_out <= rom_array(8881);
		when "0010001010110010" => data_out <= rom_array(8882);
		when "0010001010110011" => data_out <= rom_array(8883);
		when "0010001010110100" => data_out <= rom_array(8884);
		when "0010001010110101" => data_out <= rom_array(8885);
		when "0010001010110110" => data_out <= rom_array(8886);
		when "0010001010110111" => data_out <= rom_array(8887);
		when "0010001010111000" => data_out <= rom_array(8888);
		when "0010001010111001" => data_out <= rom_array(8889);
		when "0010001010111010" => data_out <= rom_array(8890);
		when "0010001010111011" => data_out <= rom_array(8891);
		when "0010001010111100" => data_out <= rom_array(8892);
		when "0010001010111101" => data_out <= rom_array(8893);
		when "0010001010111110" => data_out <= rom_array(8894);
		when "0010001010111111" => data_out <= rom_array(8895);
		when "0010001011000000" => data_out <= rom_array(8896);
		when "0010001011000001" => data_out <= rom_array(8897);
		when "0010001011000010" => data_out <= rom_array(8898);
		when "0010001011000011" => data_out <= rom_array(8899);
		when "0010001011000100" => data_out <= rom_array(8900);
		when "0010001011000101" => data_out <= rom_array(8901);
		when "0010001011000110" => data_out <= rom_array(8902);
		when "0010001011000111" => data_out <= rom_array(8903);
		when "0010001011001000" => data_out <= rom_array(8904);
		when "0010001011001001" => data_out <= rom_array(8905);
		when "0010001011001010" => data_out <= rom_array(8906);
		when "0010001011001011" => data_out <= rom_array(8907);
		when "0010001011001100" => data_out <= rom_array(8908);
		when "0010001011001101" => data_out <= rom_array(8909);
		when "0010001011001110" => data_out <= rom_array(8910);
		when "0010001011001111" => data_out <= rom_array(8911);
		when "0010001011010000" => data_out <= rom_array(8912);
		when "0010001011010001" => data_out <= rom_array(8913);
		when "0010001011010010" => data_out <= rom_array(8914);
		when "0010001011010011" => data_out <= rom_array(8915);
		when "0010001011010100" => data_out <= rom_array(8916);
		when "0010001011010101" => data_out <= rom_array(8917);
		when "0010001011010110" => data_out <= rom_array(8918);
		when "0010001011010111" => data_out <= rom_array(8919);
		when "0010001011011000" => data_out <= rom_array(8920);
		when "0010001011011001" => data_out <= rom_array(8921);
		when "0010001011011010" => data_out <= rom_array(8922);
		when "0010001011011011" => data_out <= rom_array(8923);
		when "0010001011011100" => data_out <= rom_array(8924);
		when "0010001011011101" => data_out <= rom_array(8925);
		when "0010001011011110" => data_out <= rom_array(8926);
		when "0010001011011111" => data_out <= rom_array(8927);
		when "0010001011100000" => data_out <= rom_array(8928);
		when "0010001011100001" => data_out <= rom_array(8929);
		when "0010001011100010" => data_out <= rom_array(8930);
		when "0010001011100011" => data_out <= rom_array(8931);
		when "0010001011100100" => data_out <= rom_array(8932);
		when "0010001011100101" => data_out <= rom_array(8933);
		when "0010001011100110" => data_out <= rom_array(8934);
		when "0010001011100111" => data_out <= rom_array(8935);
		when "0010001011101000" => data_out <= rom_array(8936);
		when "0010001011101001" => data_out <= rom_array(8937);
		when "0010001011101010" => data_out <= rom_array(8938);
		when "0010001011101011" => data_out <= rom_array(8939);
		when "0010001011101100" => data_out <= rom_array(8940);
		when "0010001011101101" => data_out <= rom_array(8941);
		when "0010001011101110" => data_out <= rom_array(8942);
		when "0010001011101111" => data_out <= rom_array(8943);
		when "0010001011110000" => data_out <= rom_array(8944);
		when "0010001011110001" => data_out <= rom_array(8945);
		when "0010001011110010" => data_out <= rom_array(8946);
		when "0010001011110011" => data_out <= rom_array(8947);
		when "0010001011110100" => data_out <= rom_array(8948);
		when "0010001011110101" => data_out <= rom_array(8949);
		when "0010001011110110" => data_out <= rom_array(8950);
		when "0010001011110111" => data_out <= rom_array(8951);
		when "0010001011111000" => data_out <= rom_array(8952);
		when "0010001011111001" => data_out <= rom_array(8953);
		when "0010001011111010" => data_out <= rom_array(8954);
		when "0010001011111011" => data_out <= rom_array(8955);
		when "0010001011111100" => data_out <= rom_array(8956);
		when "0010001011111101" => data_out <= rom_array(8957);
		when "0010001011111110" => data_out <= rom_array(8958);
		when "0010001011111111" => data_out <= rom_array(8959);
		when "0010001100000000" => data_out <= rom_array(8960);
		when "0010001100000001" => data_out <= rom_array(8961);
		when "0010001100000010" => data_out <= rom_array(8962);
		when "0010001100000011" => data_out <= rom_array(8963);
		when "0010001100000100" => data_out <= rom_array(8964);
		when "0010001100000101" => data_out <= rom_array(8965);
		when "0010001100000110" => data_out <= rom_array(8966);
		when "0010001100000111" => data_out <= rom_array(8967);
		when "0010001100001000" => data_out <= rom_array(8968);
		when "0010001100001001" => data_out <= rom_array(8969);
		when "0010001100001010" => data_out <= rom_array(8970);
		when "0010001100001011" => data_out <= rom_array(8971);
		when "0010001100001100" => data_out <= rom_array(8972);
		when "0010001100001101" => data_out <= rom_array(8973);
		when "0010001100001110" => data_out <= rom_array(8974);
		when "0010001100001111" => data_out <= rom_array(8975);
		when "0010001100010000" => data_out <= rom_array(8976);
		when "0010001100010001" => data_out <= rom_array(8977);
		when "0010001100010010" => data_out <= rom_array(8978);
		when "0010001100010011" => data_out <= rom_array(8979);
		when "0010001100010100" => data_out <= rom_array(8980);
		when "0010001100010101" => data_out <= rom_array(8981);
		when "0010001100010110" => data_out <= rom_array(8982);
		when "0010001100010111" => data_out <= rom_array(8983);
		when "0010001100011000" => data_out <= rom_array(8984);
		when "0010001100011001" => data_out <= rom_array(8985);
		when "0010001100011010" => data_out <= rom_array(8986);
		when "0010001100011011" => data_out <= rom_array(8987);
		when "0010001100011100" => data_out <= rom_array(8988);
		when "0010001100011101" => data_out <= rom_array(8989);
		when "0010001100011110" => data_out <= rom_array(8990);
		when "0010001100011111" => data_out <= rom_array(8991);
		when "0010001100100000" => data_out <= rom_array(8992);
		when "0010001100100001" => data_out <= rom_array(8993);
		when "0010001100100010" => data_out <= rom_array(8994);
		when "0010001100100011" => data_out <= rom_array(8995);
		when "0010001100100100" => data_out <= rom_array(8996);
		when "0010001100100101" => data_out <= rom_array(8997);
		when "0010001100100110" => data_out <= rom_array(8998);
		when "0010001100100111" => data_out <= rom_array(8999);
		when "0010001100101000" => data_out <= rom_array(9000);
		when "0010001100101001" => data_out <= rom_array(9001);
		when "0010001100101010" => data_out <= rom_array(9002);
		when "0010001100101011" => data_out <= rom_array(9003);
		when "0010001100101100" => data_out <= rom_array(9004);
		when "0010001100101101" => data_out <= rom_array(9005);
		when "0010001100101110" => data_out <= rom_array(9006);
		when "0010001100101111" => data_out <= rom_array(9007);
		when "0010001100110000" => data_out <= rom_array(9008);
		when "0010001100110001" => data_out <= rom_array(9009);
		when "0010001100110010" => data_out <= rom_array(9010);
		when "0010001100110011" => data_out <= rom_array(9011);
		when "0010001100110100" => data_out <= rom_array(9012);
		when "0010001100110101" => data_out <= rom_array(9013);
		when "0010001100110110" => data_out <= rom_array(9014);
		when "0010001100110111" => data_out <= rom_array(9015);
		when "0010001100111000" => data_out <= rom_array(9016);
		when "0010001100111001" => data_out <= rom_array(9017);
		when "0010001100111010" => data_out <= rom_array(9018);
		when "0010001100111011" => data_out <= rom_array(9019);
		when "0010001100111100" => data_out <= rom_array(9020);
		when "0010001100111101" => data_out <= rom_array(9021);
		when "0010001100111110" => data_out <= rom_array(9022);
		when "0010001100111111" => data_out <= rom_array(9023);
		when "0010001101000000" => data_out <= rom_array(9024);
		when "0010001101000001" => data_out <= rom_array(9025);
		when "0010001101000010" => data_out <= rom_array(9026);
		when "0010001101000011" => data_out <= rom_array(9027);
		when "0010001101000100" => data_out <= rom_array(9028);
		when "0010001101000101" => data_out <= rom_array(9029);
		when "0010001101000110" => data_out <= rom_array(9030);
		when "0010001101000111" => data_out <= rom_array(9031);
		when "0010001101001000" => data_out <= rom_array(9032);
		when "0010001101001001" => data_out <= rom_array(9033);
		when "0010001101001010" => data_out <= rom_array(9034);
		when "0010001101001011" => data_out <= rom_array(9035);
		when "0010001101001100" => data_out <= rom_array(9036);
		when "0010001101001101" => data_out <= rom_array(9037);
		when "0010001101001110" => data_out <= rom_array(9038);
		when "0010001101001111" => data_out <= rom_array(9039);
		when "0010001101010000" => data_out <= rom_array(9040);
		when "0010001101010001" => data_out <= rom_array(9041);
		when "0010001101010010" => data_out <= rom_array(9042);
		when "0010001101010011" => data_out <= rom_array(9043);
		when "0010001101010100" => data_out <= rom_array(9044);
		when "0010001101010101" => data_out <= rom_array(9045);
		when "0010001101010110" => data_out <= rom_array(9046);
		when "0010001101010111" => data_out <= rom_array(9047);
		when "0010001101011000" => data_out <= rom_array(9048);
		when "0010001101011001" => data_out <= rom_array(9049);
		when "0010001101011010" => data_out <= rom_array(9050);
		when "0010001101011011" => data_out <= rom_array(9051);
		when "0010001101011100" => data_out <= rom_array(9052);
		when "0010001101011101" => data_out <= rom_array(9053);
		when "0010001101011110" => data_out <= rom_array(9054);
		when "0010001101011111" => data_out <= rom_array(9055);
		when "0010001101100000" => data_out <= rom_array(9056);
		when "0010001101100001" => data_out <= rom_array(9057);
		when "0010001101100010" => data_out <= rom_array(9058);
		when "0010001101100011" => data_out <= rom_array(9059);
		when "0010001101100100" => data_out <= rom_array(9060);
		when "0010001101100101" => data_out <= rom_array(9061);
		when "0010001101100110" => data_out <= rom_array(9062);
		when "0010001101100111" => data_out <= rom_array(9063);
		when "0010001101101000" => data_out <= rom_array(9064);
		when "0010001101101001" => data_out <= rom_array(9065);
		when "0010001101101010" => data_out <= rom_array(9066);
		when "0010001101101011" => data_out <= rom_array(9067);
		when "0010001101101100" => data_out <= rom_array(9068);
		when "0010001101101101" => data_out <= rom_array(9069);
		when "0010001101101110" => data_out <= rom_array(9070);
		when "0010001101101111" => data_out <= rom_array(9071);
		when "0010001101110000" => data_out <= rom_array(9072);
		when "0010001101110001" => data_out <= rom_array(9073);
		when "0010001101110010" => data_out <= rom_array(9074);
		when "0010001101110011" => data_out <= rom_array(9075);
		when "0010001101110100" => data_out <= rom_array(9076);
		when "0010001101110101" => data_out <= rom_array(9077);
		when "0010001101110110" => data_out <= rom_array(9078);
		when "0010001101110111" => data_out <= rom_array(9079);
		when "0010001101111000" => data_out <= rom_array(9080);
		when "0010001101111001" => data_out <= rom_array(9081);
		when "0010001101111010" => data_out <= rom_array(9082);
		when "0010001101111011" => data_out <= rom_array(9083);
		when "0010001101111100" => data_out <= rom_array(9084);
		when "0010001101111101" => data_out <= rom_array(9085);
		when "0010001101111110" => data_out <= rom_array(9086);
		when "0010001101111111" => data_out <= rom_array(9087);
		when "0010001110000000" => data_out <= rom_array(9088);
		when "0010001110000001" => data_out <= rom_array(9089);
		when "0010001110000010" => data_out <= rom_array(9090);
		when "0010001110000011" => data_out <= rom_array(9091);
		when "0010001110000100" => data_out <= rom_array(9092);
		when "0010001110000101" => data_out <= rom_array(9093);
		when "0010001110000110" => data_out <= rom_array(9094);
		when "0010001110000111" => data_out <= rom_array(9095);
		when "0010001110001000" => data_out <= rom_array(9096);
		when "0010001110001001" => data_out <= rom_array(9097);
		when "0010001110001010" => data_out <= rom_array(9098);
		when "0010001110001011" => data_out <= rom_array(9099);
		when "0010001110001100" => data_out <= rom_array(9100);
		when "0010001110001101" => data_out <= rom_array(9101);
		when "0010001110001110" => data_out <= rom_array(9102);
		when "0010001110001111" => data_out <= rom_array(9103);
		when "0010001110010000" => data_out <= rom_array(9104);
		when "0010001110010001" => data_out <= rom_array(9105);
		when "0010001110010010" => data_out <= rom_array(9106);
		when "0010001110010011" => data_out <= rom_array(9107);
		when "0010001110010100" => data_out <= rom_array(9108);
		when "0010001110010101" => data_out <= rom_array(9109);
		when "0010001110010110" => data_out <= rom_array(9110);
		when "0010001110010111" => data_out <= rom_array(9111);
		when "0010001110011000" => data_out <= rom_array(9112);
		when "0010001110011001" => data_out <= rom_array(9113);
		when "0010001110011010" => data_out <= rom_array(9114);
		when "0010001110011011" => data_out <= rom_array(9115);
		when "0010001110011100" => data_out <= rom_array(9116);
		when "0010001110011101" => data_out <= rom_array(9117);
		when "0010001110011110" => data_out <= rom_array(9118);
		when "0010001110011111" => data_out <= rom_array(9119);
		when "0010001110100000" => data_out <= rom_array(9120);
		when "0010001110100001" => data_out <= rom_array(9121);
		when "0010001110100010" => data_out <= rom_array(9122);
		when "0010001110100011" => data_out <= rom_array(9123);
		when "0010001110100100" => data_out <= rom_array(9124);
		when "0010001110100101" => data_out <= rom_array(9125);
		when "0010001110100110" => data_out <= rom_array(9126);
		when "0010001110100111" => data_out <= rom_array(9127);
		when "0010001110101000" => data_out <= rom_array(9128);
		when "0010001110101001" => data_out <= rom_array(9129);
		when "0010001110101010" => data_out <= rom_array(9130);
		when "0010001110101011" => data_out <= rom_array(9131);
		when "0010001110101100" => data_out <= rom_array(9132);
		when "0010001110101101" => data_out <= rom_array(9133);
		when "0010001110101110" => data_out <= rom_array(9134);
		when "0010001110101111" => data_out <= rom_array(9135);
		when "0010001110110000" => data_out <= rom_array(9136);
		when "0010001110110001" => data_out <= rom_array(9137);
		when "0010001110110010" => data_out <= rom_array(9138);
		when "0010001110110011" => data_out <= rom_array(9139);
		when "0010001110110100" => data_out <= rom_array(9140);
		when "0010001110110101" => data_out <= rom_array(9141);
		when "0010001110110110" => data_out <= rom_array(9142);
		when "0010001110110111" => data_out <= rom_array(9143);
		when "0010001110111000" => data_out <= rom_array(9144);
		when "0010001110111001" => data_out <= rom_array(9145);
		when "0010001110111010" => data_out <= rom_array(9146);
		when "0010001110111011" => data_out <= rom_array(9147);
		when "0010001110111100" => data_out <= rom_array(9148);
		when "0010001110111101" => data_out <= rom_array(9149);
		when "0010001110111110" => data_out <= rom_array(9150);
		when "0010001110111111" => data_out <= rom_array(9151);
		when "0010001111000000" => data_out <= rom_array(9152);
		when "0010001111000001" => data_out <= rom_array(9153);
		when "0010001111000010" => data_out <= rom_array(9154);
		when "0010001111000011" => data_out <= rom_array(9155);
		when "0010001111000100" => data_out <= rom_array(9156);
		when "0010001111000101" => data_out <= rom_array(9157);
		when "0010001111000110" => data_out <= rom_array(9158);
		when "0010001111000111" => data_out <= rom_array(9159);
		when "0010001111001000" => data_out <= rom_array(9160);
		when "0010001111001001" => data_out <= rom_array(9161);
		when "0010001111001010" => data_out <= rom_array(9162);
		when "0010001111001011" => data_out <= rom_array(9163);
		when "0010001111001100" => data_out <= rom_array(9164);
		when "0010001111001101" => data_out <= rom_array(9165);
		when "0010001111001110" => data_out <= rom_array(9166);
		when "0010001111001111" => data_out <= rom_array(9167);
		when "0010001111010000" => data_out <= rom_array(9168);
		when "0010001111010001" => data_out <= rom_array(9169);
		when "0010001111010010" => data_out <= rom_array(9170);
		when "0010001111010011" => data_out <= rom_array(9171);
		when "0010001111010100" => data_out <= rom_array(9172);
		when "0010001111010101" => data_out <= rom_array(9173);
		when "0010001111010110" => data_out <= rom_array(9174);
		when "0010001111010111" => data_out <= rom_array(9175);
		when "0010001111011000" => data_out <= rom_array(9176);
		when "0010001111011001" => data_out <= rom_array(9177);
		when "0010001111011010" => data_out <= rom_array(9178);
		when "0010001111011011" => data_out <= rom_array(9179);
		when "0010001111011100" => data_out <= rom_array(9180);
		when "0010001111011101" => data_out <= rom_array(9181);
		when "0010001111011110" => data_out <= rom_array(9182);
		when "0010001111011111" => data_out <= rom_array(9183);
		when "0010001111100000" => data_out <= rom_array(9184);
		when "0010001111100001" => data_out <= rom_array(9185);
		when "0010001111100010" => data_out <= rom_array(9186);
		when "0010001111100011" => data_out <= rom_array(9187);
		when "0010001111100100" => data_out <= rom_array(9188);
		when "0010001111100101" => data_out <= rom_array(9189);
		when "0010001111100110" => data_out <= rom_array(9190);
		when "0010001111100111" => data_out <= rom_array(9191);
		when "0010001111101000" => data_out <= rom_array(9192);
		when "0010001111101001" => data_out <= rom_array(9193);
		when "0010001111101010" => data_out <= rom_array(9194);
		when "0010001111101011" => data_out <= rom_array(9195);
		when "0010001111101100" => data_out <= rom_array(9196);
		when "0010001111101101" => data_out <= rom_array(9197);
		when "0010001111101110" => data_out <= rom_array(9198);
		when "0010001111101111" => data_out <= rom_array(9199);
		when "0010001111110000" => data_out <= rom_array(9200);
		when "0010001111110001" => data_out <= rom_array(9201);
		when "0010001111110010" => data_out <= rom_array(9202);
		when "0010001111110011" => data_out <= rom_array(9203);
		when "0010001111110100" => data_out <= rom_array(9204);
		when "0010001111110101" => data_out <= rom_array(9205);
		when "0010001111110110" => data_out <= rom_array(9206);
		when "0010001111110111" => data_out <= rom_array(9207);
		when "0010001111111000" => data_out <= rom_array(9208);
		when "0010001111111001" => data_out <= rom_array(9209);
		when "0010001111111010" => data_out <= rom_array(9210);
		when "0010001111111011" => data_out <= rom_array(9211);
		when "0010001111111100" => data_out <= rom_array(9212);
		when "0010001111111101" => data_out <= rom_array(9213);
		when "0010001111111110" => data_out <= rom_array(9214);
		when "0010001111111111" => data_out <= rom_array(9215);
		when "0010010000000000" => data_out <= rom_array(9216);
		when "0010010000000001" => data_out <= rom_array(9217);
		when "0010010000000010" => data_out <= rom_array(9218);
		when "0010010000000011" => data_out <= rom_array(9219);
		when "0010010000000100" => data_out <= rom_array(9220);
		when "0010010000000101" => data_out <= rom_array(9221);
		when "0010010000000110" => data_out <= rom_array(9222);
		when "0010010000000111" => data_out <= rom_array(9223);
		when "0010010000001000" => data_out <= rom_array(9224);
		when "0010010000001001" => data_out <= rom_array(9225);
		when "0010010000001010" => data_out <= rom_array(9226);
		when "0010010000001011" => data_out <= rom_array(9227);
		when "0010010000001100" => data_out <= rom_array(9228);
		when "0010010000001101" => data_out <= rom_array(9229);
		when "0010010000001110" => data_out <= rom_array(9230);
		when "0010010000001111" => data_out <= rom_array(9231);
		when "0010010000010000" => data_out <= rom_array(9232);
		when "0010010000010001" => data_out <= rom_array(9233);
		when "0010010000010010" => data_out <= rom_array(9234);
		when "0010010000010011" => data_out <= rom_array(9235);
		when "0010010000010100" => data_out <= rom_array(9236);
		when "0010010000010101" => data_out <= rom_array(9237);
		when "0010010000010110" => data_out <= rom_array(9238);
		when "0010010000010111" => data_out <= rom_array(9239);
		when "0010010000011000" => data_out <= rom_array(9240);
		when "0010010000011001" => data_out <= rom_array(9241);
		when "0010010000011010" => data_out <= rom_array(9242);
		when "0010010000011011" => data_out <= rom_array(9243);
		when "0010010000011100" => data_out <= rom_array(9244);
		when "0010010000011101" => data_out <= rom_array(9245);
		when "0010010000011110" => data_out <= rom_array(9246);
		when "0010010000011111" => data_out <= rom_array(9247);
		when "0010010000100000" => data_out <= rom_array(9248);
		when "0010010000100001" => data_out <= rom_array(9249);
		when "0010010000100010" => data_out <= rom_array(9250);
		when "0010010000100011" => data_out <= rom_array(9251);
		when "0010010000100100" => data_out <= rom_array(9252);
		when "0010010000100101" => data_out <= rom_array(9253);
		when "0010010000100110" => data_out <= rom_array(9254);
		when "0010010000100111" => data_out <= rom_array(9255);
		when "0010010000101000" => data_out <= rom_array(9256);
		when "0010010000101001" => data_out <= rom_array(9257);
		when "0010010000101010" => data_out <= rom_array(9258);
		when "0010010000101011" => data_out <= rom_array(9259);
		when "0010010000101100" => data_out <= rom_array(9260);
		when "0010010000101101" => data_out <= rom_array(9261);
		when "0010010000101110" => data_out <= rom_array(9262);
		when "0010010000101111" => data_out <= rom_array(9263);
		when "0010010000110000" => data_out <= rom_array(9264);
		when "0010010000110001" => data_out <= rom_array(9265);
		when "0010010000110010" => data_out <= rom_array(9266);
		when "0010010000110011" => data_out <= rom_array(9267);
		when "0010010000110100" => data_out <= rom_array(9268);
		when "0010010000110101" => data_out <= rom_array(9269);
		when "0010010000110110" => data_out <= rom_array(9270);
		when "0010010000110111" => data_out <= rom_array(9271);
		when "0010010000111000" => data_out <= rom_array(9272);
		when "0010010000111001" => data_out <= rom_array(9273);
		when "0010010000111010" => data_out <= rom_array(9274);
		when "0010010000111011" => data_out <= rom_array(9275);
		when "0010010000111100" => data_out <= rom_array(9276);
		when "0010010000111101" => data_out <= rom_array(9277);
		when "0010010000111110" => data_out <= rom_array(9278);
		when "0010010000111111" => data_out <= rom_array(9279);
		when "0010010001000000" => data_out <= rom_array(9280);
		when "0010010001000001" => data_out <= rom_array(9281);
		when "0010010001000010" => data_out <= rom_array(9282);
		when "0010010001000011" => data_out <= rom_array(9283);
		when "0010010001000100" => data_out <= rom_array(9284);
		when "0010010001000101" => data_out <= rom_array(9285);
		when "0010010001000110" => data_out <= rom_array(9286);
		when "0010010001000111" => data_out <= rom_array(9287);
		when "0010010001001000" => data_out <= rom_array(9288);
		when "0010010001001001" => data_out <= rom_array(9289);
		when "0010010001001010" => data_out <= rom_array(9290);
		when "0010010001001011" => data_out <= rom_array(9291);
		when "0010010001001100" => data_out <= rom_array(9292);
		when "0010010001001101" => data_out <= rom_array(9293);
		when "0010010001001110" => data_out <= rom_array(9294);
		when "0010010001001111" => data_out <= rom_array(9295);
		when "0010010001010000" => data_out <= rom_array(9296);
		when "0010010001010001" => data_out <= rom_array(9297);
		when "0010010001010010" => data_out <= rom_array(9298);
		when "0010010001010011" => data_out <= rom_array(9299);
		when "0010010001010100" => data_out <= rom_array(9300);
		when "0010010001010101" => data_out <= rom_array(9301);
		when "0010010001010110" => data_out <= rom_array(9302);
		when "0010010001010111" => data_out <= rom_array(9303);
		when "0010010001011000" => data_out <= rom_array(9304);
		when "0010010001011001" => data_out <= rom_array(9305);
		when "0010010001011010" => data_out <= rom_array(9306);
		when "0010010001011011" => data_out <= rom_array(9307);
		when "0010010001011100" => data_out <= rom_array(9308);
		when "0010010001011101" => data_out <= rom_array(9309);
		when "0010010001011110" => data_out <= rom_array(9310);
		when "0010010001011111" => data_out <= rom_array(9311);
		when "0010010001100000" => data_out <= rom_array(9312);
		when "0010010001100001" => data_out <= rom_array(9313);
		when "0010010001100010" => data_out <= rom_array(9314);
		when "0010010001100011" => data_out <= rom_array(9315);
		when "0010010001100100" => data_out <= rom_array(9316);
		when "0010010001100101" => data_out <= rom_array(9317);
		when "0010010001100110" => data_out <= rom_array(9318);
		when "0010010001100111" => data_out <= rom_array(9319);
		when "0010010001101000" => data_out <= rom_array(9320);
		when "0010010001101001" => data_out <= rom_array(9321);
		when "0010010001101010" => data_out <= rom_array(9322);
		when "0010010001101011" => data_out <= rom_array(9323);
		when "0010010001101100" => data_out <= rom_array(9324);
		when "0010010001101101" => data_out <= rom_array(9325);
		when "0010010001101110" => data_out <= rom_array(9326);
		when "0010010001101111" => data_out <= rom_array(9327);
		when "0010010001110000" => data_out <= rom_array(9328);
		when "0010010001110001" => data_out <= rom_array(9329);
		when "0010010001110010" => data_out <= rom_array(9330);
		when "0010010001110011" => data_out <= rom_array(9331);
		when "0010010001110100" => data_out <= rom_array(9332);
		when "0010010001110101" => data_out <= rom_array(9333);
		when "0010010001110110" => data_out <= rom_array(9334);
		when "0010010001110111" => data_out <= rom_array(9335);
		when "0010010001111000" => data_out <= rom_array(9336);
		when "0010010001111001" => data_out <= rom_array(9337);
		when "0010010001111010" => data_out <= rom_array(9338);
		when "0010010001111011" => data_out <= rom_array(9339);
		when "0010010001111100" => data_out <= rom_array(9340);
		when "0010010001111101" => data_out <= rom_array(9341);
		when "0010010001111110" => data_out <= rom_array(9342);
		when "0010010001111111" => data_out <= rom_array(9343);
		when "0010010010000000" => data_out <= rom_array(9344);
		when "0010010010000001" => data_out <= rom_array(9345);
		when "0010010010000010" => data_out <= rom_array(9346);
		when "0010010010000011" => data_out <= rom_array(9347);
		when "0010010010000100" => data_out <= rom_array(9348);
		when "0010010010000101" => data_out <= rom_array(9349);
		when "0010010010000110" => data_out <= rom_array(9350);
		when "0010010010000111" => data_out <= rom_array(9351);
		when "0010010010001000" => data_out <= rom_array(9352);
		when "0010010010001001" => data_out <= rom_array(9353);
		when "0010010010001010" => data_out <= rom_array(9354);
		when "0010010010001011" => data_out <= rom_array(9355);
		when "0010010010001100" => data_out <= rom_array(9356);
		when "0010010010001101" => data_out <= rom_array(9357);
		when "0010010010001110" => data_out <= rom_array(9358);
		when "0010010010001111" => data_out <= rom_array(9359);
		when "0010010010010000" => data_out <= rom_array(9360);
		when "0010010010010001" => data_out <= rom_array(9361);
		when "0010010010010010" => data_out <= rom_array(9362);
		when "0010010010010011" => data_out <= rom_array(9363);
		when "0010010010010100" => data_out <= rom_array(9364);
		when "0010010010010101" => data_out <= rom_array(9365);
		when "0010010010010110" => data_out <= rom_array(9366);
		when "0010010010010111" => data_out <= rom_array(9367);
		when "0010010010011000" => data_out <= rom_array(9368);
		when "0010010010011001" => data_out <= rom_array(9369);
		when "0010010010011010" => data_out <= rom_array(9370);
		when "0010010010011011" => data_out <= rom_array(9371);
		when "0010010010011100" => data_out <= rom_array(9372);
		when "0010010010011101" => data_out <= rom_array(9373);
		when "0010010010011110" => data_out <= rom_array(9374);
		when "0010010010011111" => data_out <= rom_array(9375);
		when "0010010010100000" => data_out <= rom_array(9376);
		when "0010010010100001" => data_out <= rom_array(9377);
		when "0010010010100010" => data_out <= rom_array(9378);
		when "0010010010100011" => data_out <= rom_array(9379);
		when "0010010010100100" => data_out <= rom_array(9380);
		when "0010010010100101" => data_out <= rom_array(9381);
		when "0010010010100110" => data_out <= rom_array(9382);
		when "0010010010100111" => data_out <= rom_array(9383);
		when "0010010010101000" => data_out <= rom_array(9384);
		when "0010010010101001" => data_out <= rom_array(9385);
		when "0010010010101010" => data_out <= rom_array(9386);
		when "0010010010101011" => data_out <= rom_array(9387);
		when "0010010010101100" => data_out <= rom_array(9388);
		when "0010010010101101" => data_out <= rom_array(9389);
		when "0010010010101110" => data_out <= rom_array(9390);
		when "0010010010101111" => data_out <= rom_array(9391);
		when "0010010010110000" => data_out <= rom_array(9392);
		when "0010010010110001" => data_out <= rom_array(9393);
		when "0010010010110010" => data_out <= rom_array(9394);
		when "0010010010110011" => data_out <= rom_array(9395);
		when "0010010010110100" => data_out <= rom_array(9396);
		when "0010010010110101" => data_out <= rom_array(9397);
		when "0010010010110110" => data_out <= rom_array(9398);
		when "0010010010110111" => data_out <= rom_array(9399);
		when "0010010010111000" => data_out <= rom_array(9400);
		when "0010010010111001" => data_out <= rom_array(9401);
		when "0010010010111010" => data_out <= rom_array(9402);
		when "0010010010111011" => data_out <= rom_array(9403);
		when "0010010010111100" => data_out <= rom_array(9404);
		when "0010010010111101" => data_out <= rom_array(9405);
		when "0010010010111110" => data_out <= rom_array(9406);
		when "0010010010111111" => data_out <= rom_array(9407);
		when "0010010011000000" => data_out <= rom_array(9408);
		when "0010010011000001" => data_out <= rom_array(9409);
		when "0010010011000010" => data_out <= rom_array(9410);
		when "0010010011000011" => data_out <= rom_array(9411);
		when "0010010011000100" => data_out <= rom_array(9412);
		when "0010010011000101" => data_out <= rom_array(9413);
		when "0010010011000110" => data_out <= rom_array(9414);
		when "0010010011000111" => data_out <= rom_array(9415);
		when "0010010011001000" => data_out <= rom_array(9416);
		when "0010010011001001" => data_out <= rom_array(9417);
		when "0010010011001010" => data_out <= rom_array(9418);
		when "0010010011001011" => data_out <= rom_array(9419);
		when "0010010011001100" => data_out <= rom_array(9420);
		when "0010010011001101" => data_out <= rom_array(9421);
		when "0010010011001110" => data_out <= rom_array(9422);
		when "0010010011001111" => data_out <= rom_array(9423);
		when "0010010011010000" => data_out <= rom_array(9424);
		when "0010010011010001" => data_out <= rom_array(9425);
		when "0010010011010010" => data_out <= rom_array(9426);
		when "0010010011010011" => data_out <= rom_array(9427);
		when "0010010011010100" => data_out <= rom_array(9428);
		when "0010010011010101" => data_out <= rom_array(9429);
		when "0010010011010110" => data_out <= rom_array(9430);
		when "0010010011010111" => data_out <= rom_array(9431);
		when "0010010011011000" => data_out <= rom_array(9432);
		when "0010010011011001" => data_out <= rom_array(9433);
		when "0010010011011010" => data_out <= rom_array(9434);
		when "0010010011011011" => data_out <= rom_array(9435);
		when "0010010011011100" => data_out <= rom_array(9436);
		when "0010010011011101" => data_out <= rom_array(9437);
		when "0010010011011110" => data_out <= rom_array(9438);
		when "0010010011011111" => data_out <= rom_array(9439);
		when "0010010011100000" => data_out <= rom_array(9440);
		when "0010010011100001" => data_out <= rom_array(9441);
		when "0010010011100010" => data_out <= rom_array(9442);
		when "0010010011100011" => data_out <= rom_array(9443);
		when "0010010011100100" => data_out <= rom_array(9444);
		when "0010010011100101" => data_out <= rom_array(9445);
		when "0010010011100110" => data_out <= rom_array(9446);
		when "0010010011100111" => data_out <= rom_array(9447);
		when "0010010011101000" => data_out <= rom_array(9448);
		when "0010010011101001" => data_out <= rom_array(9449);
		when "0010010011101010" => data_out <= rom_array(9450);
		when "0010010011101011" => data_out <= rom_array(9451);
		when "0010010011101100" => data_out <= rom_array(9452);
		when "0010010011101101" => data_out <= rom_array(9453);
		when "0010010011101110" => data_out <= rom_array(9454);
		when "0010010011101111" => data_out <= rom_array(9455);
		when "0010010011110000" => data_out <= rom_array(9456);
		when "0010010011110001" => data_out <= rom_array(9457);
		when "0010010011110010" => data_out <= rom_array(9458);
		when "0010010011110011" => data_out <= rom_array(9459);
		when "0010010011110100" => data_out <= rom_array(9460);
		when "0010010011110101" => data_out <= rom_array(9461);
		when "0010010011110110" => data_out <= rom_array(9462);
		when "0010010011110111" => data_out <= rom_array(9463);
		when "0010010011111000" => data_out <= rom_array(9464);
		when "0010010011111001" => data_out <= rom_array(9465);
		when "0010010011111010" => data_out <= rom_array(9466);
		when "0010010011111011" => data_out <= rom_array(9467);
		when "0010010011111100" => data_out <= rom_array(9468);
		when "0010010011111101" => data_out <= rom_array(9469);
		when "0010010011111110" => data_out <= rom_array(9470);
		when "0010010011111111" => data_out <= rom_array(9471);
		when "0010010100000000" => data_out <= rom_array(9472);
		when "0010010100000001" => data_out <= rom_array(9473);
		when "0010010100000010" => data_out <= rom_array(9474);
		when "0010010100000011" => data_out <= rom_array(9475);
		when "0010010100000100" => data_out <= rom_array(9476);
		when "0010010100000101" => data_out <= rom_array(9477);
		when "0010010100000110" => data_out <= rom_array(9478);
		when "0010010100000111" => data_out <= rom_array(9479);
		when "0010010100001000" => data_out <= rom_array(9480);
		when "0010010100001001" => data_out <= rom_array(9481);
		when "0010010100001010" => data_out <= rom_array(9482);
		when "0010010100001011" => data_out <= rom_array(9483);
		when "0010010100001100" => data_out <= rom_array(9484);
		when "0010010100001101" => data_out <= rom_array(9485);
		when "0010010100001110" => data_out <= rom_array(9486);
		when "0010010100001111" => data_out <= rom_array(9487);
		when "0010010100010000" => data_out <= rom_array(9488);
		when "0010010100010001" => data_out <= rom_array(9489);
		when "0010010100010010" => data_out <= rom_array(9490);
		when "0010010100010011" => data_out <= rom_array(9491);
		when "0010010100010100" => data_out <= rom_array(9492);
		when "0010010100010101" => data_out <= rom_array(9493);
		when "0010010100010110" => data_out <= rom_array(9494);
		when "0010010100010111" => data_out <= rom_array(9495);
		when "0010010100011000" => data_out <= rom_array(9496);
		when "0010010100011001" => data_out <= rom_array(9497);
		when "0010010100011010" => data_out <= rom_array(9498);
		when "0010010100011011" => data_out <= rom_array(9499);
		when "0010010100011100" => data_out <= rom_array(9500);
		when "0010010100011101" => data_out <= rom_array(9501);
		when "0010010100011110" => data_out <= rom_array(9502);
		when "0010010100011111" => data_out <= rom_array(9503);
		when "0010010100100000" => data_out <= rom_array(9504);
		when "0010010100100001" => data_out <= rom_array(9505);
		when "0010010100100010" => data_out <= rom_array(9506);
		when "0010010100100011" => data_out <= rom_array(9507);
		when "0010010100100100" => data_out <= rom_array(9508);
		when "0010010100100101" => data_out <= rom_array(9509);
		when "0010010100100110" => data_out <= rom_array(9510);
		when "0010010100100111" => data_out <= rom_array(9511);
		when "0010010100101000" => data_out <= rom_array(9512);
		when "0010010100101001" => data_out <= rom_array(9513);
		when "0010010100101010" => data_out <= rom_array(9514);
		when "0010010100101011" => data_out <= rom_array(9515);
		when "0010010100101100" => data_out <= rom_array(9516);
		when "0010010100101101" => data_out <= rom_array(9517);
		when "0010010100101110" => data_out <= rom_array(9518);
		when "0010010100101111" => data_out <= rom_array(9519);
		when "0010010100110000" => data_out <= rom_array(9520);
		when "0010010100110001" => data_out <= rom_array(9521);
		when "0010010100110010" => data_out <= rom_array(9522);
		when "0010010100110011" => data_out <= rom_array(9523);
		when "0010010100110100" => data_out <= rom_array(9524);
		when "0010010100110101" => data_out <= rom_array(9525);
		when "0010010100110110" => data_out <= rom_array(9526);
		when "0010010100110111" => data_out <= rom_array(9527);
		when "0010010100111000" => data_out <= rom_array(9528);
		when "0010010100111001" => data_out <= rom_array(9529);
		when "0010010100111010" => data_out <= rom_array(9530);
		when "0010010100111011" => data_out <= rom_array(9531);
		when "0010010100111100" => data_out <= rom_array(9532);
		when "0010010100111101" => data_out <= rom_array(9533);
		when "0010010100111110" => data_out <= rom_array(9534);
		when "0010010100111111" => data_out <= rom_array(9535);
		when "0010010101000000" => data_out <= rom_array(9536);
		when "0010010101000001" => data_out <= rom_array(9537);
		when "0010010101000010" => data_out <= rom_array(9538);
		when "0010010101000011" => data_out <= rom_array(9539);
		when "0010010101000100" => data_out <= rom_array(9540);
		when "0010010101000101" => data_out <= rom_array(9541);
		when "0010010101000110" => data_out <= rom_array(9542);
		when "0010010101000111" => data_out <= rom_array(9543);
		when "0010010101001000" => data_out <= rom_array(9544);
		when "0010010101001001" => data_out <= rom_array(9545);
		when "0010010101001010" => data_out <= rom_array(9546);
		when "0010010101001011" => data_out <= rom_array(9547);
		when "0010010101001100" => data_out <= rom_array(9548);
		when "0010010101001101" => data_out <= rom_array(9549);
		when "0010010101001110" => data_out <= rom_array(9550);
		when "0010010101001111" => data_out <= rom_array(9551);
		when "0010010101010000" => data_out <= rom_array(9552);
		when "0010010101010001" => data_out <= rom_array(9553);
		when "0010010101010010" => data_out <= rom_array(9554);
		when "0010010101010011" => data_out <= rom_array(9555);
		when "0010010101010100" => data_out <= rom_array(9556);
		when "0010010101010101" => data_out <= rom_array(9557);
		when "0010010101010110" => data_out <= rom_array(9558);
		when "0010010101010111" => data_out <= rom_array(9559);
		when "0010010101011000" => data_out <= rom_array(9560);
		when "0010010101011001" => data_out <= rom_array(9561);
		when "0010010101011010" => data_out <= rom_array(9562);
		when "0010010101011011" => data_out <= rom_array(9563);
		when "0010010101011100" => data_out <= rom_array(9564);
		when "0010010101011101" => data_out <= rom_array(9565);
		when "0010010101011110" => data_out <= rom_array(9566);
		when "0010010101011111" => data_out <= rom_array(9567);
		when "0010010101100000" => data_out <= rom_array(9568);
		when "0010010101100001" => data_out <= rom_array(9569);
		when "0010010101100010" => data_out <= rom_array(9570);
		when "0010010101100011" => data_out <= rom_array(9571);
		when "0010010101100100" => data_out <= rom_array(9572);
		when "0010010101100101" => data_out <= rom_array(9573);
		when "0010010101100110" => data_out <= rom_array(9574);
		when "0010010101100111" => data_out <= rom_array(9575);
		when "0010010101101000" => data_out <= rom_array(9576);
		when "0010010101101001" => data_out <= rom_array(9577);
		when "0010010101101010" => data_out <= rom_array(9578);
		when "0010010101101011" => data_out <= rom_array(9579);
		when "0010010101101100" => data_out <= rom_array(9580);
		when "0010010101101101" => data_out <= rom_array(9581);
		when "0010010101101110" => data_out <= rom_array(9582);
		when "0010010101101111" => data_out <= rom_array(9583);
		when "0010010101110000" => data_out <= rom_array(9584);
		when "0010010101110001" => data_out <= rom_array(9585);
		when "0010010101110010" => data_out <= rom_array(9586);
		when "0010010101110011" => data_out <= rom_array(9587);
		when "0010010101110100" => data_out <= rom_array(9588);
		when "0010010101110101" => data_out <= rom_array(9589);
		when "0010010101110110" => data_out <= rom_array(9590);
		when "0010010101110111" => data_out <= rom_array(9591);
		when "0010010101111000" => data_out <= rom_array(9592);
		when "0010010101111001" => data_out <= rom_array(9593);
		when "0010010101111010" => data_out <= rom_array(9594);
		when "0010010101111011" => data_out <= rom_array(9595);
		when "0010010101111100" => data_out <= rom_array(9596);
		when "0010010101111101" => data_out <= rom_array(9597);
		when "0010010101111110" => data_out <= rom_array(9598);
		when "0010010101111111" => data_out <= rom_array(9599);
		when "0010010110000000" => data_out <= rom_array(9600);
		when "0010010110000001" => data_out <= rom_array(9601);
		when "0010010110000010" => data_out <= rom_array(9602);
		when "0010010110000011" => data_out <= rom_array(9603);
		when "0010010110000100" => data_out <= rom_array(9604);
		when "0010010110000101" => data_out <= rom_array(9605);
		when "0010010110000110" => data_out <= rom_array(9606);
		when "0010010110000111" => data_out <= rom_array(9607);
		when "0010010110001000" => data_out <= rom_array(9608);
		when "0010010110001001" => data_out <= rom_array(9609);
		when "0010010110001010" => data_out <= rom_array(9610);
		when "0010010110001011" => data_out <= rom_array(9611);
		when "0010010110001100" => data_out <= rom_array(9612);
		when "0010010110001101" => data_out <= rom_array(9613);
		when "0010010110001110" => data_out <= rom_array(9614);
		when "0010010110001111" => data_out <= rom_array(9615);
		when "0010010110010000" => data_out <= rom_array(9616);
		when "0010010110010001" => data_out <= rom_array(9617);
		when "0010010110010010" => data_out <= rom_array(9618);
		when "0010010110010011" => data_out <= rom_array(9619);
		when "0010010110010100" => data_out <= rom_array(9620);
		when "0010010110010101" => data_out <= rom_array(9621);
		when "0010010110010110" => data_out <= rom_array(9622);
		when "0010010110010111" => data_out <= rom_array(9623);
		when "0010010110011000" => data_out <= rom_array(9624);
		when "0010010110011001" => data_out <= rom_array(9625);
		when "0010010110011010" => data_out <= rom_array(9626);
		when "0010010110011011" => data_out <= rom_array(9627);
		when "0010010110011100" => data_out <= rom_array(9628);
		when "0010010110011101" => data_out <= rom_array(9629);
		when "0010010110011110" => data_out <= rom_array(9630);
		when "0010010110011111" => data_out <= rom_array(9631);
		when "0010010110100000" => data_out <= rom_array(9632);
		when "0010010110100001" => data_out <= rom_array(9633);
		when "0010010110100010" => data_out <= rom_array(9634);
		when "0010010110100011" => data_out <= rom_array(9635);
		when "0010010110100100" => data_out <= rom_array(9636);
		when "0010010110100101" => data_out <= rom_array(9637);
		when "0010010110100110" => data_out <= rom_array(9638);
		when "0010010110100111" => data_out <= rom_array(9639);
		when "0010010110101000" => data_out <= rom_array(9640);
		when "0010010110101001" => data_out <= rom_array(9641);
		when "0010010110101010" => data_out <= rom_array(9642);
		when "0010010110101011" => data_out <= rom_array(9643);
		when "0010010110101100" => data_out <= rom_array(9644);
		when "0010010110101101" => data_out <= rom_array(9645);
		when "0010010110101110" => data_out <= rom_array(9646);
		when "0010010110101111" => data_out <= rom_array(9647);
		when "0010010110110000" => data_out <= rom_array(9648);
		when "0010010110110001" => data_out <= rom_array(9649);
		when "0010010110110010" => data_out <= rom_array(9650);
		when "0010010110110011" => data_out <= rom_array(9651);
		when "0010010110110100" => data_out <= rom_array(9652);
		when "0010010110110101" => data_out <= rom_array(9653);
		when "0010010110110110" => data_out <= rom_array(9654);
		when "0010010110110111" => data_out <= rom_array(9655);
		when "0010010110111000" => data_out <= rom_array(9656);
		when "0010010110111001" => data_out <= rom_array(9657);
		when "0010010110111010" => data_out <= rom_array(9658);
		when "0010010110111011" => data_out <= rom_array(9659);
		when "0010010110111100" => data_out <= rom_array(9660);
		when "0010010110111101" => data_out <= rom_array(9661);
		when "0010010110111110" => data_out <= rom_array(9662);
		when "0010010110111111" => data_out <= rom_array(9663);
		when "0010010111000000" => data_out <= rom_array(9664);
		when "0010010111000001" => data_out <= rom_array(9665);
		when "0010010111000010" => data_out <= rom_array(9666);
		when "0010010111000011" => data_out <= rom_array(9667);
		when "0010010111000100" => data_out <= rom_array(9668);
		when "0010010111000101" => data_out <= rom_array(9669);
		when "0010010111000110" => data_out <= rom_array(9670);
		when "0010010111000111" => data_out <= rom_array(9671);
		when "0010010111001000" => data_out <= rom_array(9672);
		when "0010010111001001" => data_out <= rom_array(9673);
		when "0010010111001010" => data_out <= rom_array(9674);
		when "0010010111001011" => data_out <= rom_array(9675);
		when "0010010111001100" => data_out <= rom_array(9676);
		when "0010010111001101" => data_out <= rom_array(9677);
		when "0010010111001110" => data_out <= rom_array(9678);
		when "0010010111001111" => data_out <= rom_array(9679);
		when "0010010111010000" => data_out <= rom_array(9680);
		when "0010010111010001" => data_out <= rom_array(9681);
		when "0010010111010010" => data_out <= rom_array(9682);
		when "0010010111010011" => data_out <= rom_array(9683);
		when "0010010111010100" => data_out <= rom_array(9684);
		when "0010010111010101" => data_out <= rom_array(9685);
		when "0010010111010110" => data_out <= rom_array(9686);
		when "0010010111010111" => data_out <= rom_array(9687);
		when "0010010111011000" => data_out <= rom_array(9688);
		when "0010010111011001" => data_out <= rom_array(9689);
		when "0010010111011010" => data_out <= rom_array(9690);
		when "0010010111011011" => data_out <= rom_array(9691);
		when "0010010111011100" => data_out <= rom_array(9692);
		when "0010010111011101" => data_out <= rom_array(9693);
		when "0010010111011110" => data_out <= rom_array(9694);
		when "0010010111011111" => data_out <= rom_array(9695);
		when "0010010111100000" => data_out <= rom_array(9696);
		when "0010010111100001" => data_out <= rom_array(9697);
		when "0010010111100010" => data_out <= rom_array(9698);
		when "0010010111100011" => data_out <= rom_array(9699);
		when "0010010111100100" => data_out <= rom_array(9700);
		when "0010010111100101" => data_out <= rom_array(9701);
		when "0010010111100110" => data_out <= rom_array(9702);
		when "0010010111100111" => data_out <= rom_array(9703);
		when "0010010111101000" => data_out <= rom_array(9704);
		when "0010010111101001" => data_out <= rom_array(9705);
		when "0010010111101010" => data_out <= rom_array(9706);
		when "0010010111101011" => data_out <= rom_array(9707);
		when "0010010111101100" => data_out <= rom_array(9708);
		when "0010010111101101" => data_out <= rom_array(9709);
		when "0010010111101110" => data_out <= rom_array(9710);
		when "0010010111101111" => data_out <= rom_array(9711);
		when "0010010111110000" => data_out <= rom_array(9712);
		when "0010010111110001" => data_out <= rom_array(9713);
		when "0010010111110010" => data_out <= rom_array(9714);
		when "0010010111110011" => data_out <= rom_array(9715);
		when "0010010111110100" => data_out <= rom_array(9716);
		when "0010010111110101" => data_out <= rom_array(9717);
		when "0010010111110110" => data_out <= rom_array(9718);
		when "0010010111110111" => data_out <= rom_array(9719);
		when "0010010111111000" => data_out <= rom_array(9720);
		when "0010010111111001" => data_out <= rom_array(9721);
		when "0010010111111010" => data_out <= rom_array(9722);
		when "0010010111111011" => data_out <= rom_array(9723);
		when "0010010111111100" => data_out <= rom_array(9724);
		when "0010010111111101" => data_out <= rom_array(9725);
		when "0010010111111110" => data_out <= rom_array(9726);
		when "0010010111111111" => data_out <= rom_array(9727);
		when "0010011000000000" => data_out <= rom_array(9728);
		when "0010011000000001" => data_out <= rom_array(9729);
		when "0010011000000010" => data_out <= rom_array(9730);
		when "0010011000000011" => data_out <= rom_array(9731);
		when "0010011000000100" => data_out <= rom_array(9732);
		when "0010011000000101" => data_out <= rom_array(9733);
		when "0010011000000110" => data_out <= rom_array(9734);
		when "0010011000000111" => data_out <= rom_array(9735);
		when "0010011000001000" => data_out <= rom_array(9736);
		when "0010011000001001" => data_out <= rom_array(9737);
		when "0010011000001010" => data_out <= rom_array(9738);
		when "0010011000001011" => data_out <= rom_array(9739);
		when "0010011000001100" => data_out <= rom_array(9740);
		when "0010011000001101" => data_out <= rom_array(9741);
		when "0010011000001110" => data_out <= rom_array(9742);
		when "0010011000001111" => data_out <= rom_array(9743);
		when "0010011000010000" => data_out <= rom_array(9744);
		when "0010011000010001" => data_out <= rom_array(9745);
		when "0010011000010010" => data_out <= rom_array(9746);
		when "0010011000010011" => data_out <= rom_array(9747);
		when "0010011000010100" => data_out <= rom_array(9748);
		when "0010011000010101" => data_out <= rom_array(9749);
		when "0010011000010110" => data_out <= rom_array(9750);
		when "0010011000010111" => data_out <= rom_array(9751);
		when "0010011000011000" => data_out <= rom_array(9752);
		when "0010011000011001" => data_out <= rom_array(9753);
		when "0010011000011010" => data_out <= rom_array(9754);
		when "0010011000011011" => data_out <= rom_array(9755);
		when "0010011000011100" => data_out <= rom_array(9756);
		when "0010011000011101" => data_out <= rom_array(9757);
		when "0010011000011110" => data_out <= rom_array(9758);
		when "0010011000011111" => data_out <= rom_array(9759);
		when "0010011000100000" => data_out <= rom_array(9760);
		when "0010011000100001" => data_out <= rom_array(9761);
		when "0010011000100010" => data_out <= rom_array(9762);
		when "0010011000100011" => data_out <= rom_array(9763);
		when "0010011000100100" => data_out <= rom_array(9764);
		when "0010011000100101" => data_out <= rom_array(9765);
		when "0010011000100110" => data_out <= rom_array(9766);
		when "0010011000100111" => data_out <= rom_array(9767);
		when "0010011000101000" => data_out <= rom_array(9768);
		when "0010011000101001" => data_out <= rom_array(9769);
		when "0010011000101010" => data_out <= rom_array(9770);
		when "0010011000101011" => data_out <= rom_array(9771);
		when "0010011000101100" => data_out <= rom_array(9772);
		when "0010011000101101" => data_out <= rom_array(9773);
		when "0010011000101110" => data_out <= rom_array(9774);
		when "0010011000101111" => data_out <= rom_array(9775);
		when "0010011000110000" => data_out <= rom_array(9776);
		when "0010011000110001" => data_out <= rom_array(9777);
		when "0010011000110010" => data_out <= rom_array(9778);
		when "0010011000110011" => data_out <= rom_array(9779);
		when "0010011000110100" => data_out <= rom_array(9780);
		when "0010011000110101" => data_out <= rom_array(9781);
		when "0010011000110110" => data_out <= rom_array(9782);
		when "0010011000110111" => data_out <= rom_array(9783);
		when "0010011000111000" => data_out <= rom_array(9784);
		when "0010011000111001" => data_out <= rom_array(9785);
		when "0010011000111010" => data_out <= rom_array(9786);
		when "0010011000111011" => data_out <= rom_array(9787);
		when "0010011000111100" => data_out <= rom_array(9788);
		when "0010011000111101" => data_out <= rom_array(9789);
		when "0010011000111110" => data_out <= rom_array(9790);
		when "0010011000111111" => data_out <= rom_array(9791);
		when "0010011001000000" => data_out <= rom_array(9792);
		when "0010011001000001" => data_out <= rom_array(9793);
		when "0010011001000010" => data_out <= rom_array(9794);
		when "0010011001000011" => data_out <= rom_array(9795);
		when "0010011001000100" => data_out <= rom_array(9796);
		when "0010011001000101" => data_out <= rom_array(9797);
		when "0010011001000110" => data_out <= rom_array(9798);
		when "0010011001000111" => data_out <= rom_array(9799);
		when "0010011001001000" => data_out <= rom_array(9800);
		when "0010011001001001" => data_out <= rom_array(9801);
		when "0010011001001010" => data_out <= rom_array(9802);
		when "0010011001001011" => data_out <= rom_array(9803);
		when "0010011001001100" => data_out <= rom_array(9804);
		when "0010011001001101" => data_out <= rom_array(9805);
		when "0010011001001110" => data_out <= rom_array(9806);
		when "0010011001001111" => data_out <= rom_array(9807);
		when "0010011001010000" => data_out <= rom_array(9808);
		when "0010011001010001" => data_out <= rom_array(9809);
		when "0010011001010010" => data_out <= rom_array(9810);
		when "0010011001010011" => data_out <= rom_array(9811);
		when "0010011001010100" => data_out <= rom_array(9812);
		when "0010011001010101" => data_out <= rom_array(9813);
		when "0010011001010110" => data_out <= rom_array(9814);
		when "0010011001010111" => data_out <= rom_array(9815);
		when "0010011001011000" => data_out <= rom_array(9816);
		when "0010011001011001" => data_out <= rom_array(9817);
		when "0010011001011010" => data_out <= rom_array(9818);
		when "0010011001011011" => data_out <= rom_array(9819);
		when "0010011001011100" => data_out <= rom_array(9820);
		when "0010011001011101" => data_out <= rom_array(9821);
		when "0010011001011110" => data_out <= rom_array(9822);
		when "0010011001011111" => data_out <= rom_array(9823);
		when "0010011001100000" => data_out <= rom_array(9824);
		when "0010011001100001" => data_out <= rom_array(9825);
		when "0010011001100010" => data_out <= rom_array(9826);
		when "0010011001100011" => data_out <= rom_array(9827);
		when "0010011001100100" => data_out <= rom_array(9828);
		when "0010011001100101" => data_out <= rom_array(9829);
		when "0010011001100110" => data_out <= rom_array(9830);
		when "0010011001100111" => data_out <= rom_array(9831);
		when "0010011001101000" => data_out <= rom_array(9832);
		when "0010011001101001" => data_out <= rom_array(9833);
		when "0010011001101010" => data_out <= rom_array(9834);
		when "0010011001101011" => data_out <= rom_array(9835);
		when "0010011001101100" => data_out <= rom_array(9836);
		when "0010011001101101" => data_out <= rom_array(9837);
		when "0010011001101110" => data_out <= rom_array(9838);
		when "0010011001101111" => data_out <= rom_array(9839);
		when "0010011001110000" => data_out <= rom_array(9840);
		when "0010011001110001" => data_out <= rom_array(9841);
		when "0010011001110010" => data_out <= rom_array(9842);
		when "0010011001110011" => data_out <= rom_array(9843);
		when "0010011001110100" => data_out <= rom_array(9844);
		when "0010011001110101" => data_out <= rom_array(9845);
		when "0010011001110110" => data_out <= rom_array(9846);
		when "0010011001110111" => data_out <= rom_array(9847);
		when "0010011001111000" => data_out <= rom_array(9848);
		when "0010011001111001" => data_out <= rom_array(9849);
		when "0010011001111010" => data_out <= rom_array(9850);
		when "0010011001111011" => data_out <= rom_array(9851);
		when "0010011001111100" => data_out <= rom_array(9852);
		when "0010011001111101" => data_out <= rom_array(9853);
		when "0010011001111110" => data_out <= rom_array(9854);
		when "0010011001111111" => data_out <= rom_array(9855);
		when "0010011010000000" => data_out <= rom_array(9856);
		when "0010011010000001" => data_out <= rom_array(9857);
		when "0010011010000010" => data_out <= rom_array(9858);
		when "0010011010000011" => data_out <= rom_array(9859);
		when "0010011010000100" => data_out <= rom_array(9860);
		when "0010011010000101" => data_out <= rom_array(9861);
		when "0010011010000110" => data_out <= rom_array(9862);
		when "0010011010000111" => data_out <= rom_array(9863);
		when "0010011010001000" => data_out <= rom_array(9864);
		when "0010011010001001" => data_out <= rom_array(9865);
		when "0010011010001010" => data_out <= rom_array(9866);
		when "0010011010001011" => data_out <= rom_array(9867);
		when "0010011010001100" => data_out <= rom_array(9868);
		when "0010011010001101" => data_out <= rom_array(9869);
		when "0010011010001110" => data_out <= rom_array(9870);
		when "0010011010001111" => data_out <= rom_array(9871);
		when "0010011010010000" => data_out <= rom_array(9872);
		when "0010011010010001" => data_out <= rom_array(9873);
		when "0010011010010010" => data_out <= rom_array(9874);
		when "0010011010010011" => data_out <= rom_array(9875);
		when "0010011010010100" => data_out <= rom_array(9876);
		when "0010011010010101" => data_out <= rom_array(9877);
		when "0010011010010110" => data_out <= rom_array(9878);
		when "0010011010010111" => data_out <= rom_array(9879);
		when "0010011010011000" => data_out <= rom_array(9880);
		when "0010011010011001" => data_out <= rom_array(9881);
		when "0010011010011010" => data_out <= rom_array(9882);
		when "0010011010011011" => data_out <= rom_array(9883);
		when "0010011010011100" => data_out <= rom_array(9884);
		when "0010011010011101" => data_out <= rom_array(9885);
		when "0010011010011110" => data_out <= rom_array(9886);
		when "0010011010011111" => data_out <= rom_array(9887);
		when "0010011010100000" => data_out <= rom_array(9888);
		when "0010011010100001" => data_out <= rom_array(9889);
		when "0010011010100010" => data_out <= rom_array(9890);
		when "0010011010100011" => data_out <= rom_array(9891);
		when "0010011010100100" => data_out <= rom_array(9892);
		when "0010011010100101" => data_out <= rom_array(9893);
		when "0010011010100110" => data_out <= rom_array(9894);
		when "0010011010100111" => data_out <= rom_array(9895);
		when "0010011010101000" => data_out <= rom_array(9896);
		when "0010011010101001" => data_out <= rom_array(9897);
		when "0010011010101010" => data_out <= rom_array(9898);
		when "0010011010101011" => data_out <= rom_array(9899);
		when "0010011010101100" => data_out <= rom_array(9900);
		when "0010011010101101" => data_out <= rom_array(9901);
		when "0010011010101110" => data_out <= rom_array(9902);
		when "0010011010101111" => data_out <= rom_array(9903);
		when "0010011010110000" => data_out <= rom_array(9904);
		when "0010011010110001" => data_out <= rom_array(9905);
		when "0010011010110010" => data_out <= rom_array(9906);
		when "0010011010110011" => data_out <= rom_array(9907);
		when "0010011010110100" => data_out <= rom_array(9908);
		when "0010011010110101" => data_out <= rom_array(9909);
		when "0010011010110110" => data_out <= rom_array(9910);
		when "0010011010110111" => data_out <= rom_array(9911);
		when "0010011010111000" => data_out <= rom_array(9912);
		when "0010011010111001" => data_out <= rom_array(9913);
		when "0010011010111010" => data_out <= rom_array(9914);
		when "0010011010111011" => data_out <= rom_array(9915);
		when "0010011010111100" => data_out <= rom_array(9916);
		when "0010011010111101" => data_out <= rom_array(9917);
		when "0010011010111110" => data_out <= rom_array(9918);
		when "0010011010111111" => data_out <= rom_array(9919);
		when "0010011011000000" => data_out <= rom_array(9920);
		when "0010011011000001" => data_out <= rom_array(9921);
		when "0010011011000010" => data_out <= rom_array(9922);
		when "0010011011000011" => data_out <= rom_array(9923);
		when "0010011011000100" => data_out <= rom_array(9924);
		when "0010011011000101" => data_out <= rom_array(9925);
		when "0010011011000110" => data_out <= rom_array(9926);
		when "0010011011000111" => data_out <= rom_array(9927);
		when "0010011011001000" => data_out <= rom_array(9928);
		when "0010011011001001" => data_out <= rom_array(9929);
		when "0010011011001010" => data_out <= rom_array(9930);
		when "0010011011001011" => data_out <= rom_array(9931);
		when "0010011011001100" => data_out <= rom_array(9932);
		when "0010011011001101" => data_out <= rom_array(9933);
		when "0010011011001110" => data_out <= rom_array(9934);
		when "0010011011001111" => data_out <= rom_array(9935);
		when "0010011011010000" => data_out <= rom_array(9936);
		when "0010011011010001" => data_out <= rom_array(9937);
		when "0010011011010010" => data_out <= rom_array(9938);
		when "0010011011010011" => data_out <= rom_array(9939);
		when "0010011011010100" => data_out <= rom_array(9940);
		when "0010011011010101" => data_out <= rom_array(9941);
		when "0010011011010110" => data_out <= rom_array(9942);
		when "0010011011010111" => data_out <= rom_array(9943);
		when "0010011011011000" => data_out <= rom_array(9944);
		when "0010011011011001" => data_out <= rom_array(9945);
		when "0010011011011010" => data_out <= rom_array(9946);
		when "0010011011011011" => data_out <= rom_array(9947);
		when "0010011011011100" => data_out <= rom_array(9948);
		when "0010011011011101" => data_out <= rom_array(9949);
		when "0010011011011110" => data_out <= rom_array(9950);
		when "0010011011011111" => data_out <= rom_array(9951);
		when "0010011011100000" => data_out <= rom_array(9952);
		when "0010011011100001" => data_out <= rom_array(9953);
		when "0010011011100010" => data_out <= rom_array(9954);
		when "0010011011100011" => data_out <= rom_array(9955);
		when "0010011011100100" => data_out <= rom_array(9956);
		when "0010011011100101" => data_out <= rom_array(9957);
		when "0010011011100110" => data_out <= rom_array(9958);
		when "0010011011100111" => data_out <= rom_array(9959);
		when "0010011011101000" => data_out <= rom_array(9960);
		when "0010011011101001" => data_out <= rom_array(9961);
		when "0010011011101010" => data_out <= rom_array(9962);
		when "0010011011101011" => data_out <= rom_array(9963);
		when "0010011011101100" => data_out <= rom_array(9964);
		when "0010011011101101" => data_out <= rom_array(9965);
		when "0010011011101110" => data_out <= rom_array(9966);
		when "0010011011101111" => data_out <= rom_array(9967);
		when "0010011011110000" => data_out <= rom_array(9968);
		when "0010011011110001" => data_out <= rom_array(9969);
		when "0010011011110010" => data_out <= rom_array(9970);
		when "0010011011110011" => data_out <= rom_array(9971);
		when "0010011011110100" => data_out <= rom_array(9972);
		when "0010011011110101" => data_out <= rom_array(9973);
		when "0010011011110110" => data_out <= rom_array(9974);
		when "0010011011110111" => data_out <= rom_array(9975);
		when "0010011011111000" => data_out <= rom_array(9976);
		when "0010011011111001" => data_out <= rom_array(9977);
		when "0010011011111010" => data_out <= rom_array(9978);
		when "0010011011111011" => data_out <= rom_array(9979);
		when "0010011011111100" => data_out <= rom_array(9980);
		when "0010011011111101" => data_out <= rom_array(9981);
		when "0010011011111110" => data_out <= rom_array(9982);
		when "0010011011111111" => data_out <= rom_array(9983);
		when "0010011100000000" => data_out <= rom_array(9984);
		when "0010011100000001" => data_out <= rom_array(9985);
		when "0010011100000010" => data_out <= rom_array(9986);
		when "0010011100000011" => data_out <= rom_array(9987);
		when "0010011100000100" => data_out <= rom_array(9988);
		when "0010011100000101" => data_out <= rom_array(9989);
		when "0010011100000110" => data_out <= rom_array(9990);
		when "0010011100000111" => data_out <= rom_array(9991);
		when "0010011100001000" => data_out <= rom_array(9992);
		when "0010011100001001" => data_out <= rom_array(9993);
		when "0010011100001010" => data_out <= rom_array(9994);
		when "0010011100001011" => data_out <= rom_array(9995);
		when "0010011100001100" => data_out <= rom_array(9996);
		when "0010011100001101" => data_out <= rom_array(9997);
		when "0010011100001110" => data_out <= rom_array(9998);
		when "0010011100001111" => data_out <= rom_array(9999);
		when "0010011100010000" => data_out <= rom_array(10000);
		when "0010011100010001" => data_out <= rom_array(10001);
		when "0010011100010010" => data_out <= rom_array(10002);
		when "0010011100010011" => data_out <= rom_array(10003);
		when "0010011100010100" => data_out <= rom_array(10004);
		when "0010011100010101" => data_out <= rom_array(10005);
		when "0010011100010110" => data_out <= rom_array(10006);
		when "0010011100010111" => data_out <= rom_array(10007);
		when "0010011100011000" => data_out <= rom_array(10008);
		when "0010011100011001" => data_out <= rom_array(10009);
		when "0010011100011010" => data_out <= rom_array(10010);
		when "0010011100011011" => data_out <= rom_array(10011);
		when "0010011100011100" => data_out <= rom_array(10012);
		when "0010011100011101" => data_out <= rom_array(10013);
		when "0010011100011110" => data_out <= rom_array(10014);
		when "0010011100011111" => data_out <= rom_array(10015);
		when "0010011100100000" => data_out <= rom_array(10016);
		when "0010011100100001" => data_out <= rom_array(10017);
		when "0010011100100010" => data_out <= rom_array(10018);
		when "0010011100100011" => data_out <= rom_array(10019);
		when "0010011100100100" => data_out <= rom_array(10020);
		when "0010011100100101" => data_out <= rom_array(10021);
		when "0010011100100110" => data_out <= rom_array(10022);
		when "0010011100100111" => data_out <= rom_array(10023);
		when "0010011100101000" => data_out <= rom_array(10024);
		when "0010011100101001" => data_out <= rom_array(10025);
		when "0010011100101010" => data_out <= rom_array(10026);
		when "0010011100101011" => data_out <= rom_array(10027);
		when "0010011100101100" => data_out <= rom_array(10028);
		when "0010011100101101" => data_out <= rom_array(10029);
		when "0010011100101110" => data_out <= rom_array(10030);
		when "0010011100101111" => data_out <= rom_array(10031);
		when "0010011100110000" => data_out <= rom_array(10032);
		when "0010011100110001" => data_out <= rom_array(10033);
		when "0010011100110010" => data_out <= rom_array(10034);
		when "0010011100110011" => data_out <= rom_array(10035);
		when "0010011100110100" => data_out <= rom_array(10036);
		when "0010011100110101" => data_out <= rom_array(10037);
		when "0010011100110110" => data_out <= rom_array(10038);
		when "0010011100110111" => data_out <= rom_array(10039);
		when "0010011100111000" => data_out <= rom_array(10040);
		when "0010011100111001" => data_out <= rom_array(10041);
		when "0010011100111010" => data_out <= rom_array(10042);
		when "0010011100111011" => data_out <= rom_array(10043);
		when "0010011100111100" => data_out <= rom_array(10044);
		when "0010011100111101" => data_out <= rom_array(10045);
		when "0010011100111110" => data_out <= rom_array(10046);
		when "0010011100111111" => data_out <= rom_array(10047);
		when "0010011101000000" => data_out <= rom_array(10048);
		when "0010011101000001" => data_out <= rom_array(10049);
		when "0010011101000010" => data_out <= rom_array(10050);
		when "0010011101000011" => data_out <= rom_array(10051);
		when "0010011101000100" => data_out <= rom_array(10052);
		when "0010011101000101" => data_out <= rom_array(10053);
		when "0010011101000110" => data_out <= rom_array(10054);
		when "0010011101000111" => data_out <= rom_array(10055);
		when "0010011101001000" => data_out <= rom_array(10056);
		when "0010011101001001" => data_out <= rom_array(10057);
		when "0010011101001010" => data_out <= rom_array(10058);
		when "0010011101001011" => data_out <= rom_array(10059);
		when "0010011101001100" => data_out <= rom_array(10060);
		when "0010011101001101" => data_out <= rom_array(10061);
		when "0010011101001110" => data_out <= rom_array(10062);
		when "0010011101001111" => data_out <= rom_array(10063);
		when "0010011101010000" => data_out <= rom_array(10064);
		when "0010011101010001" => data_out <= rom_array(10065);
		when "0010011101010010" => data_out <= rom_array(10066);
		when "0010011101010011" => data_out <= rom_array(10067);
		when "0010011101010100" => data_out <= rom_array(10068);
		when "0010011101010101" => data_out <= rom_array(10069);
		when "0010011101010110" => data_out <= rom_array(10070);
		when "0010011101010111" => data_out <= rom_array(10071);
		when "0010011101011000" => data_out <= rom_array(10072);
		when "0010011101011001" => data_out <= rom_array(10073);
		when "0010011101011010" => data_out <= rom_array(10074);
		when "0010011101011011" => data_out <= rom_array(10075);
		when "0010011101011100" => data_out <= rom_array(10076);
		when "0010011101011101" => data_out <= rom_array(10077);
		when "0010011101011110" => data_out <= rom_array(10078);
		when "0010011101011111" => data_out <= rom_array(10079);
		when "0010011101100000" => data_out <= rom_array(10080);
		when "0010011101100001" => data_out <= rom_array(10081);
		when "0010011101100010" => data_out <= rom_array(10082);
		when "0010011101100011" => data_out <= rom_array(10083);
		when "0010011101100100" => data_out <= rom_array(10084);
		when "0010011101100101" => data_out <= rom_array(10085);
		when "0010011101100110" => data_out <= rom_array(10086);
		when "0010011101100111" => data_out <= rom_array(10087);
		when "0010011101101000" => data_out <= rom_array(10088);
		when "0010011101101001" => data_out <= rom_array(10089);
		when "0010011101101010" => data_out <= rom_array(10090);
		when "0010011101101011" => data_out <= rom_array(10091);
		when "0010011101101100" => data_out <= rom_array(10092);
		when "0010011101101101" => data_out <= rom_array(10093);
		when "0010011101101110" => data_out <= rom_array(10094);
		when "0010011101101111" => data_out <= rom_array(10095);
		when "0010011101110000" => data_out <= rom_array(10096);
		when "0010011101110001" => data_out <= rom_array(10097);
		when "0010011101110010" => data_out <= rom_array(10098);
		when "0010011101110011" => data_out <= rom_array(10099);
		when "0010011101110100" => data_out <= rom_array(10100);
		when "0010011101110101" => data_out <= rom_array(10101);
		when "0010011101110110" => data_out <= rom_array(10102);
		when "0010011101110111" => data_out <= rom_array(10103);
		when "0010011101111000" => data_out <= rom_array(10104);
		when "0010011101111001" => data_out <= rom_array(10105);
		when "0010011101111010" => data_out <= rom_array(10106);
		when "0010011101111011" => data_out <= rom_array(10107);
		when "0010011101111100" => data_out <= rom_array(10108);
		when "0010011101111101" => data_out <= rom_array(10109);
		when "0010011101111110" => data_out <= rom_array(10110);
		when "0010011101111111" => data_out <= rom_array(10111);
		when "0010011110000000" => data_out <= rom_array(10112);
		when "0010011110000001" => data_out <= rom_array(10113);
		when "0010011110000010" => data_out <= rom_array(10114);
		when "0010011110000011" => data_out <= rom_array(10115);
		when "0010011110000100" => data_out <= rom_array(10116);
		when "0010011110000101" => data_out <= rom_array(10117);
		when "0010011110000110" => data_out <= rom_array(10118);
		when "0010011110000111" => data_out <= rom_array(10119);
		when "0010011110001000" => data_out <= rom_array(10120);
		when "0010011110001001" => data_out <= rom_array(10121);
		when "0010011110001010" => data_out <= rom_array(10122);
		when "0010011110001011" => data_out <= rom_array(10123);
		when "0010011110001100" => data_out <= rom_array(10124);
		when "0010011110001101" => data_out <= rom_array(10125);
		when "0010011110001110" => data_out <= rom_array(10126);
		when "0010011110001111" => data_out <= rom_array(10127);
		when "0010011110010000" => data_out <= rom_array(10128);
		when "0010011110010001" => data_out <= rom_array(10129);
		when "0010011110010010" => data_out <= rom_array(10130);
		when "0010011110010011" => data_out <= rom_array(10131);
		when "0010011110010100" => data_out <= rom_array(10132);
		when "0010011110010101" => data_out <= rom_array(10133);
		when "0010011110010110" => data_out <= rom_array(10134);
		when "0010011110010111" => data_out <= rom_array(10135);
		when "0010011110011000" => data_out <= rom_array(10136);
		when "0010011110011001" => data_out <= rom_array(10137);
		when "0010011110011010" => data_out <= rom_array(10138);
		when "0010011110011011" => data_out <= rom_array(10139);
		when "0010011110011100" => data_out <= rom_array(10140);
		when "0010011110011101" => data_out <= rom_array(10141);
		when "0010011110011110" => data_out <= rom_array(10142);
		when "0010011110011111" => data_out <= rom_array(10143);
		when "0010011110100000" => data_out <= rom_array(10144);
		when "0010011110100001" => data_out <= rom_array(10145);
		when "0010011110100010" => data_out <= rom_array(10146);
		when "0010011110100011" => data_out <= rom_array(10147);
		when "0010011110100100" => data_out <= rom_array(10148);
		when "0010011110100101" => data_out <= rom_array(10149);
		when "0010011110100110" => data_out <= rom_array(10150);
		when "0010011110100111" => data_out <= rom_array(10151);
		when "0010011110101000" => data_out <= rom_array(10152);
		when "0010011110101001" => data_out <= rom_array(10153);
		when "0010011110101010" => data_out <= rom_array(10154);
		when "0010011110101011" => data_out <= rom_array(10155);
		when "0010011110101100" => data_out <= rom_array(10156);
		when "0010011110101101" => data_out <= rom_array(10157);
		when "0010011110101110" => data_out <= rom_array(10158);
		when "0010011110101111" => data_out <= rom_array(10159);
		when "0010011110110000" => data_out <= rom_array(10160);
		when "0010011110110001" => data_out <= rom_array(10161);
		when "0010011110110010" => data_out <= rom_array(10162);
		when "0010011110110011" => data_out <= rom_array(10163);
		when "0010011110110100" => data_out <= rom_array(10164);
		when "0010011110110101" => data_out <= rom_array(10165);
		when "0010011110110110" => data_out <= rom_array(10166);
		when "0010011110110111" => data_out <= rom_array(10167);
		when "0010011110111000" => data_out <= rom_array(10168);
		when "0010011110111001" => data_out <= rom_array(10169);
		when "0010011110111010" => data_out <= rom_array(10170);
		when "0010011110111011" => data_out <= rom_array(10171);
		when "0010011110111100" => data_out <= rom_array(10172);
		when "0010011110111101" => data_out <= rom_array(10173);
		when "0010011110111110" => data_out <= rom_array(10174);
		when "0010011110111111" => data_out <= rom_array(10175);
		when "0010011111000000" => data_out <= rom_array(10176);
		when "0010011111000001" => data_out <= rom_array(10177);
		when "0010011111000010" => data_out <= rom_array(10178);
		when "0010011111000011" => data_out <= rom_array(10179);
		when "0010011111000100" => data_out <= rom_array(10180);
		when "0010011111000101" => data_out <= rom_array(10181);
		when "0010011111000110" => data_out <= rom_array(10182);
		when "0010011111000111" => data_out <= rom_array(10183);
		when "0010011111001000" => data_out <= rom_array(10184);
		when "0010011111001001" => data_out <= rom_array(10185);
		when "0010011111001010" => data_out <= rom_array(10186);
		when "0010011111001011" => data_out <= rom_array(10187);
		when "0010011111001100" => data_out <= rom_array(10188);
		when "0010011111001101" => data_out <= rom_array(10189);
		when "0010011111001110" => data_out <= rom_array(10190);
		when "0010011111001111" => data_out <= rom_array(10191);
		when "0010011111010000" => data_out <= rom_array(10192);
		when "0010011111010001" => data_out <= rom_array(10193);
		when "0010011111010010" => data_out <= rom_array(10194);
		when "0010011111010011" => data_out <= rom_array(10195);
		when "0010011111010100" => data_out <= rom_array(10196);
		when "0010011111010101" => data_out <= rom_array(10197);
		when "0010011111010110" => data_out <= rom_array(10198);
		when "0010011111010111" => data_out <= rom_array(10199);
		when "0010011111011000" => data_out <= rom_array(10200);
		when "0010011111011001" => data_out <= rom_array(10201);
		when "0010011111011010" => data_out <= rom_array(10202);
		when "0010011111011011" => data_out <= rom_array(10203);
		when "0010011111011100" => data_out <= rom_array(10204);
		when "0010011111011101" => data_out <= rom_array(10205);
		when "0010011111011110" => data_out <= rom_array(10206);
		when "0010011111011111" => data_out <= rom_array(10207);
		when "0010011111100000" => data_out <= rom_array(10208);
		when "0010011111100001" => data_out <= rom_array(10209);
		when "0010011111100010" => data_out <= rom_array(10210);
		when "0010011111100011" => data_out <= rom_array(10211);
		when "0010011111100100" => data_out <= rom_array(10212);
		when "0010011111100101" => data_out <= rom_array(10213);
		when "0010011111100110" => data_out <= rom_array(10214);
		when "0010011111100111" => data_out <= rom_array(10215);
		when "0010011111101000" => data_out <= rom_array(10216);
		when "0010011111101001" => data_out <= rom_array(10217);
		when "0010011111101010" => data_out <= rom_array(10218);
		when "0010011111101011" => data_out <= rom_array(10219);
		when "0010011111101100" => data_out <= rom_array(10220);
		when "0010011111101101" => data_out <= rom_array(10221);
		when "0010011111101110" => data_out <= rom_array(10222);
		when "0010011111101111" => data_out <= rom_array(10223);
		when "0010011111110000" => data_out <= rom_array(10224);
		when "0010011111110001" => data_out <= rom_array(10225);
		when "0010011111110010" => data_out <= rom_array(10226);
		when "0010011111110011" => data_out <= rom_array(10227);
		when "0010011111110100" => data_out <= rom_array(10228);
		when "0010011111110101" => data_out <= rom_array(10229);
		when "0010011111110110" => data_out <= rom_array(10230);
		when "0010011111110111" => data_out <= rom_array(10231);
		when "0010011111111000" => data_out <= rom_array(10232);
		when "0010011111111001" => data_out <= rom_array(10233);
		when "0010011111111010" => data_out <= rom_array(10234);
		when "0010011111111011" => data_out <= rom_array(10235);
		when "0010011111111100" => data_out <= rom_array(10236);
		when "0010011111111101" => data_out <= rom_array(10237);
		when "0010011111111110" => data_out <= rom_array(10238);
		when "0010011111111111" => data_out <= rom_array(10239);
		when "0010100000000000" => data_out <= rom_array(10240);
		when "0010100000000001" => data_out <= rom_array(10241);
		when "0010100000000010" => data_out <= rom_array(10242);
		when "0010100000000011" => data_out <= rom_array(10243);
		when "0010100000000100" => data_out <= rom_array(10244);
		when "0010100000000101" => data_out <= rom_array(10245);
		when "0010100000000110" => data_out <= rom_array(10246);
		when "0010100000000111" => data_out <= rom_array(10247);
		when "0010100000001000" => data_out <= rom_array(10248);
		when "0010100000001001" => data_out <= rom_array(10249);
		when "0010100000001010" => data_out <= rom_array(10250);
		when "0010100000001011" => data_out <= rom_array(10251);
		when "0010100000001100" => data_out <= rom_array(10252);
		when "0010100000001101" => data_out <= rom_array(10253);
		when "0010100000001110" => data_out <= rom_array(10254);
		when "0010100000001111" => data_out <= rom_array(10255);
		when "0010100000010000" => data_out <= rom_array(10256);
		when "0010100000010001" => data_out <= rom_array(10257);
		when "0010100000010010" => data_out <= rom_array(10258);
		when "0010100000010011" => data_out <= rom_array(10259);
		when "0010100000010100" => data_out <= rom_array(10260);
		when "0010100000010101" => data_out <= rom_array(10261);
		when "0010100000010110" => data_out <= rom_array(10262);
		when "0010100000010111" => data_out <= rom_array(10263);
		when "0010100000011000" => data_out <= rom_array(10264);
		when "0010100000011001" => data_out <= rom_array(10265);
		when "0010100000011010" => data_out <= rom_array(10266);
		when "0010100000011011" => data_out <= rom_array(10267);
		when "0010100000011100" => data_out <= rom_array(10268);
		when "0010100000011101" => data_out <= rom_array(10269);
		when "0010100000011110" => data_out <= rom_array(10270);
		when "0010100000011111" => data_out <= rom_array(10271);
		when "0010100000100000" => data_out <= rom_array(10272);
		when "0010100000100001" => data_out <= rom_array(10273);
		when "0010100000100010" => data_out <= rom_array(10274);
		when "0010100000100011" => data_out <= rom_array(10275);
		when "0010100000100100" => data_out <= rom_array(10276);
		when "0010100000100101" => data_out <= rom_array(10277);
		when "0010100000100110" => data_out <= rom_array(10278);
		when "0010100000100111" => data_out <= rom_array(10279);
		when "0010100000101000" => data_out <= rom_array(10280);
		when "0010100000101001" => data_out <= rom_array(10281);
		when "0010100000101010" => data_out <= rom_array(10282);
		when "0010100000101011" => data_out <= rom_array(10283);
		when "0010100000101100" => data_out <= rom_array(10284);
		when "0010100000101101" => data_out <= rom_array(10285);
		when "0010100000101110" => data_out <= rom_array(10286);
		when "0010100000101111" => data_out <= rom_array(10287);
		when "0010100000110000" => data_out <= rom_array(10288);
		when "0010100000110001" => data_out <= rom_array(10289);
		when "0010100000110010" => data_out <= rom_array(10290);
		when "0010100000110011" => data_out <= rom_array(10291);
		when "0010100000110100" => data_out <= rom_array(10292);
		when "0010100000110101" => data_out <= rom_array(10293);
		when "0010100000110110" => data_out <= rom_array(10294);
		when "0010100000110111" => data_out <= rom_array(10295);
		when "0010100000111000" => data_out <= rom_array(10296);
		when "0010100000111001" => data_out <= rom_array(10297);
		when "0010100000111010" => data_out <= rom_array(10298);
		when "0010100000111011" => data_out <= rom_array(10299);
		when "0010100000111100" => data_out <= rom_array(10300);
		when "0010100000111101" => data_out <= rom_array(10301);
		when "0010100000111110" => data_out <= rom_array(10302);
		when "0010100000111111" => data_out <= rom_array(10303);
		when "0010100001000000" => data_out <= rom_array(10304);
		when "0010100001000001" => data_out <= rom_array(10305);
		when "0010100001000010" => data_out <= rom_array(10306);
		when "0010100001000011" => data_out <= rom_array(10307);
		when "0010100001000100" => data_out <= rom_array(10308);
		when "0010100001000101" => data_out <= rom_array(10309);
		when "0010100001000110" => data_out <= rom_array(10310);
		when "0010100001000111" => data_out <= rom_array(10311);
		when "0010100001001000" => data_out <= rom_array(10312);
		when "0010100001001001" => data_out <= rom_array(10313);
		when "0010100001001010" => data_out <= rom_array(10314);
		when "0010100001001011" => data_out <= rom_array(10315);
		when "0010100001001100" => data_out <= rom_array(10316);
		when "0010100001001101" => data_out <= rom_array(10317);
		when "0010100001001110" => data_out <= rom_array(10318);
		when "0010100001001111" => data_out <= rom_array(10319);
		when "0010100001010000" => data_out <= rom_array(10320);
		when "0010100001010001" => data_out <= rom_array(10321);
		when "0010100001010010" => data_out <= rom_array(10322);
		when "0010100001010011" => data_out <= rom_array(10323);
		when "0010100001010100" => data_out <= rom_array(10324);
		when "0010100001010101" => data_out <= rom_array(10325);
		when "0010100001010110" => data_out <= rom_array(10326);
		when "0010100001010111" => data_out <= rom_array(10327);
		when "0010100001011000" => data_out <= rom_array(10328);
		when "0010100001011001" => data_out <= rom_array(10329);
		when "0010100001011010" => data_out <= rom_array(10330);
		when "0010100001011011" => data_out <= rom_array(10331);
		when "0010100001011100" => data_out <= rom_array(10332);
		when "0010100001011101" => data_out <= rom_array(10333);
		when "0010100001011110" => data_out <= rom_array(10334);
		when "0010100001011111" => data_out <= rom_array(10335);
		when "0010100001100000" => data_out <= rom_array(10336);
		when "0010100001100001" => data_out <= rom_array(10337);
		when "0010100001100010" => data_out <= rom_array(10338);
		when "0010100001100011" => data_out <= rom_array(10339);
		when "0010100001100100" => data_out <= rom_array(10340);
		when "0010100001100101" => data_out <= rom_array(10341);
		when "0010100001100110" => data_out <= rom_array(10342);
		when "0010100001100111" => data_out <= rom_array(10343);
		when "0010100001101000" => data_out <= rom_array(10344);
		when "0010100001101001" => data_out <= rom_array(10345);
		when "0010100001101010" => data_out <= rom_array(10346);
		when "0010100001101011" => data_out <= rom_array(10347);
		when "0010100001101100" => data_out <= rom_array(10348);
		when "0010100001101101" => data_out <= rom_array(10349);
		when "0010100001101110" => data_out <= rom_array(10350);
		when "0010100001101111" => data_out <= rom_array(10351);
		when "0010100001110000" => data_out <= rom_array(10352);
		when "0010100001110001" => data_out <= rom_array(10353);
		when "0010100001110010" => data_out <= rom_array(10354);
		when "0010100001110011" => data_out <= rom_array(10355);
		when "0010100001110100" => data_out <= rom_array(10356);
		when "0010100001110101" => data_out <= rom_array(10357);
		when "0010100001110110" => data_out <= rom_array(10358);
		when "0010100001110111" => data_out <= rom_array(10359);
		when "0010100001111000" => data_out <= rom_array(10360);
		when "0010100001111001" => data_out <= rom_array(10361);
		when "0010100001111010" => data_out <= rom_array(10362);
		when "0010100001111011" => data_out <= rom_array(10363);
		when "0010100001111100" => data_out <= rom_array(10364);
		when "0010100001111101" => data_out <= rom_array(10365);
		when "0010100001111110" => data_out <= rom_array(10366);
		when "0010100001111111" => data_out <= rom_array(10367);
		when "0010100010000000" => data_out <= rom_array(10368);
		when "0010100010000001" => data_out <= rom_array(10369);
		when "0010100010000010" => data_out <= rom_array(10370);
		when "0010100010000011" => data_out <= rom_array(10371);
		when "0010100010000100" => data_out <= rom_array(10372);
		when "0010100010000101" => data_out <= rom_array(10373);
		when "0010100010000110" => data_out <= rom_array(10374);
		when "0010100010000111" => data_out <= rom_array(10375);
		when "0010100010001000" => data_out <= rom_array(10376);
		when "0010100010001001" => data_out <= rom_array(10377);
		when "0010100010001010" => data_out <= rom_array(10378);
		when "0010100010001011" => data_out <= rom_array(10379);
		when "0010100010001100" => data_out <= rom_array(10380);
		when "0010100010001101" => data_out <= rom_array(10381);
		when "0010100010001110" => data_out <= rom_array(10382);
		when "0010100010001111" => data_out <= rom_array(10383);
		when "0010100010010000" => data_out <= rom_array(10384);
		when "0010100010010001" => data_out <= rom_array(10385);
		when "0010100010010010" => data_out <= rom_array(10386);
		when "0010100010010011" => data_out <= rom_array(10387);
		when "0010100010010100" => data_out <= rom_array(10388);
		when "0010100010010101" => data_out <= rom_array(10389);
		when "0010100010010110" => data_out <= rom_array(10390);
		when "0010100010010111" => data_out <= rom_array(10391);
		when "0010100010011000" => data_out <= rom_array(10392);
		when "0010100010011001" => data_out <= rom_array(10393);
		when "0010100010011010" => data_out <= rom_array(10394);
		when "0010100010011011" => data_out <= rom_array(10395);
		when "0010100010011100" => data_out <= rom_array(10396);
		when "0010100010011101" => data_out <= rom_array(10397);
		when "0010100010011110" => data_out <= rom_array(10398);
		when "0010100010011111" => data_out <= rom_array(10399);
		when "0010100010100000" => data_out <= rom_array(10400);
		when "0010100010100001" => data_out <= rom_array(10401);
		when "0010100010100010" => data_out <= rom_array(10402);
		when "0010100010100011" => data_out <= rom_array(10403);
		when "0010100010100100" => data_out <= rom_array(10404);
		when "0010100010100101" => data_out <= rom_array(10405);
		when "0010100010100110" => data_out <= rom_array(10406);
		when "0010100010100111" => data_out <= rom_array(10407);
		when "0010100010101000" => data_out <= rom_array(10408);
		when "0010100010101001" => data_out <= rom_array(10409);
		when "0010100010101010" => data_out <= rom_array(10410);
		when "0010100010101011" => data_out <= rom_array(10411);
		when "0010100010101100" => data_out <= rom_array(10412);
		when "0010100010101101" => data_out <= rom_array(10413);
		when "0010100010101110" => data_out <= rom_array(10414);
		when "0010100010101111" => data_out <= rom_array(10415);
		when "0010100010110000" => data_out <= rom_array(10416);
		when "0010100010110001" => data_out <= rom_array(10417);
		when "0010100010110010" => data_out <= rom_array(10418);
		when "0010100010110011" => data_out <= rom_array(10419);
		when "0010100010110100" => data_out <= rom_array(10420);
		when "0010100010110101" => data_out <= rom_array(10421);
		when "0010100010110110" => data_out <= rom_array(10422);
		when "0010100010110111" => data_out <= rom_array(10423);
		when "0010100010111000" => data_out <= rom_array(10424);
		when "0010100010111001" => data_out <= rom_array(10425);
		when "0010100010111010" => data_out <= rom_array(10426);
		when "0010100010111011" => data_out <= rom_array(10427);
		when "0010100010111100" => data_out <= rom_array(10428);
		when "0010100010111101" => data_out <= rom_array(10429);
		when "0010100010111110" => data_out <= rom_array(10430);
		when "0010100010111111" => data_out <= rom_array(10431);
		when "0010100011000000" => data_out <= rom_array(10432);
		when "0010100011000001" => data_out <= rom_array(10433);
		when "0010100011000010" => data_out <= rom_array(10434);
		when "0010100011000011" => data_out <= rom_array(10435);
		when "0010100011000100" => data_out <= rom_array(10436);
		when "0010100011000101" => data_out <= rom_array(10437);
		when "0010100011000110" => data_out <= rom_array(10438);
		when "0010100011000111" => data_out <= rom_array(10439);
		when "0010100011001000" => data_out <= rom_array(10440);
		when "0010100011001001" => data_out <= rom_array(10441);
		when "0010100011001010" => data_out <= rom_array(10442);
		when "0010100011001011" => data_out <= rom_array(10443);
		when "0010100011001100" => data_out <= rom_array(10444);
		when "0010100011001101" => data_out <= rom_array(10445);
		when "0010100011001110" => data_out <= rom_array(10446);
		when "0010100011001111" => data_out <= rom_array(10447);
		when "0010100011010000" => data_out <= rom_array(10448);
		when "0010100011010001" => data_out <= rom_array(10449);
		when "0010100011010010" => data_out <= rom_array(10450);
		when "0010100011010011" => data_out <= rom_array(10451);
		when "0010100011010100" => data_out <= rom_array(10452);
		when "0010100011010101" => data_out <= rom_array(10453);
		when "0010100011010110" => data_out <= rom_array(10454);
		when "0010100011010111" => data_out <= rom_array(10455);
		when "0010100011011000" => data_out <= rom_array(10456);
		when "0010100011011001" => data_out <= rom_array(10457);
		when "0010100011011010" => data_out <= rom_array(10458);
		when "0010100011011011" => data_out <= rom_array(10459);
		when "0010100011011100" => data_out <= rom_array(10460);
		when "0010100011011101" => data_out <= rom_array(10461);
		when "0010100011011110" => data_out <= rom_array(10462);
		when "0010100011011111" => data_out <= rom_array(10463);
		when "0010100011100000" => data_out <= rom_array(10464);
		when "0010100011100001" => data_out <= rom_array(10465);
		when "0010100011100010" => data_out <= rom_array(10466);
		when "0010100011100011" => data_out <= rom_array(10467);
		when "0010100011100100" => data_out <= rom_array(10468);
		when "0010100011100101" => data_out <= rom_array(10469);
		when "0010100011100110" => data_out <= rom_array(10470);
		when "0010100011100111" => data_out <= rom_array(10471);
		when "0010100011101000" => data_out <= rom_array(10472);
		when "0010100011101001" => data_out <= rom_array(10473);
		when "0010100011101010" => data_out <= rom_array(10474);
		when "0010100011101011" => data_out <= rom_array(10475);
		when "0010100011101100" => data_out <= rom_array(10476);
		when "0010100011101101" => data_out <= rom_array(10477);
		when "0010100011101110" => data_out <= rom_array(10478);
		when "0010100011101111" => data_out <= rom_array(10479);
		when "0010100011110000" => data_out <= rom_array(10480);
		when "0010100011110001" => data_out <= rom_array(10481);
		when "0010100011110010" => data_out <= rom_array(10482);
		when "0010100011110011" => data_out <= rom_array(10483);
		when "0010100011110100" => data_out <= rom_array(10484);
		when "0010100011110101" => data_out <= rom_array(10485);
		when "0010100011110110" => data_out <= rom_array(10486);
		when "0010100011110111" => data_out <= rom_array(10487);
		when "0010100011111000" => data_out <= rom_array(10488);
		when "0010100011111001" => data_out <= rom_array(10489);
		when "0010100011111010" => data_out <= rom_array(10490);
		when "0010100011111011" => data_out <= rom_array(10491);
		when "0010100011111100" => data_out <= rom_array(10492);
		when "0010100011111101" => data_out <= rom_array(10493);
		when "0010100011111110" => data_out <= rom_array(10494);
		when "0010100011111111" => data_out <= rom_array(10495);
		when "0010100100000000" => data_out <= rom_array(10496);
		when "0010100100000001" => data_out <= rom_array(10497);
		when "0010100100000010" => data_out <= rom_array(10498);
		when "0010100100000011" => data_out <= rom_array(10499);
		when "0010100100000100" => data_out <= rom_array(10500);
		when "0010100100000101" => data_out <= rom_array(10501);
		when "0010100100000110" => data_out <= rom_array(10502);
		when "0010100100000111" => data_out <= rom_array(10503);
		when "0010100100001000" => data_out <= rom_array(10504);
		when "0010100100001001" => data_out <= rom_array(10505);
		when "0010100100001010" => data_out <= rom_array(10506);
		when "0010100100001011" => data_out <= rom_array(10507);
		when "0010100100001100" => data_out <= rom_array(10508);
		when "0010100100001101" => data_out <= rom_array(10509);
		when "0010100100001110" => data_out <= rom_array(10510);
		when "0010100100001111" => data_out <= rom_array(10511);
		when "0010100100010000" => data_out <= rom_array(10512);
		when "0010100100010001" => data_out <= rom_array(10513);
		when "0010100100010010" => data_out <= rom_array(10514);
		when "0010100100010011" => data_out <= rom_array(10515);
		when "0010100100010100" => data_out <= rom_array(10516);
		when "0010100100010101" => data_out <= rom_array(10517);
		when "0010100100010110" => data_out <= rom_array(10518);
		when "0010100100010111" => data_out <= rom_array(10519);
		when "0010100100011000" => data_out <= rom_array(10520);
		when "0010100100011001" => data_out <= rom_array(10521);
		when "0010100100011010" => data_out <= rom_array(10522);
		when "0010100100011011" => data_out <= rom_array(10523);
		when "0010100100011100" => data_out <= rom_array(10524);
		when "0010100100011101" => data_out <= rom_array(10525);
		when "0010100100011110" => data_out <= rom_array(10526);
		when "0010100100011111" => data_out <= rom_array(10527);
		when "0010100100100000" => data_out <= rom_array(10528);
		when "0010100100100001" => data_out <= rom_array(10529);
		when "0010100100100010" => data_out <= rom_array(10530);
		when "0010100100100011" => data_out <= rom_array(10531);
		when "0010100100100100" => data_out <= rom_array(10532);
		when "0010100100100101" => data_out <= rom_array(10533);
		when "0010100100100110" => data_out <= rom_array(10534);
		when "0010100100100111" => data_out <= rom_array(10535);
		when "0010100100101000" => data_out <= rom_array(10536);
		when "0010100100101001" => data_out <= rom_array(10537);
		when "0010100100101010" => data_out <= rom_array(10538);
		when "0010100100101011" => data_out <= rom_array(10539);
		when "0010100100101100" => data_out <= rom_array(10540);
		when "0010100100101101" => data_out <= rom_array(10541);
		when "0010100100101110" => data_out <= rom_array(10542);
		when "0010100100101111" => data_out <= rom_array(10543);
		when "0010100100110000" => data_out <= rom_array(10544);
		when "0010100100110001" => data_out <= rom_array(10545);
		when "0010100100110010" => data_out <= rom_array(10546);
		when "0010100100110011" => data_out <= rom_array(10547);
		when "0010100100110100" => data_out <= rom_array(10548);
		when "0010100100110101" => data_out <= rom_array(10549);
		when "0010100100110110" => data_out <= rom_array(10550);
		when "0010100100110111" => data_out <= rom_array(10551);
		when "0010100100111000" => data_out <= rom_array(10552);
		when "0010100100111001" => data_out <= rom_array(10553);
		when "0010100100111010" => data_out <= rom_array(10554);
		when "0010100100111011" => data_out <= rom_array(10555);
		when "0010100100111100" => data_out <= rom_array(10556);
		when "0010100100111101" => data_out <= rom_array(10557);
		when "0010100100111110" => data_out <= rom_array(10558);
		when "0010100100111111" => data_out <= rom_array(10559);
		when "0010100101000000" => data_out <= rom_array(10560);
		when "0010100101000001" => data_out <= rom_array(10561);
		when "0010100101000010" => data_out <= rom_array(10562);
		when "0010100101000011" => data_out <= rom_array(10563);
		when "0010100101000100" => data_out <= rom_array(10564);
		when "0010100101000101" => data_out <= rom_array(10565);
		when "0010100101000110" => data_out <= rom_array(10566);
		when "0010100101000111" => data_out <= rom_array(10567);
		when "0010100101001000" => data_out <= rom_array(10568);
		when "0010100101001001" => data_out <= rom_array(10569);
		when "0010100101001010" => data_out <= rom_array(10570);
		when "0010100101001011" => data_out <= rom_array(10571);
		when "0010100101001100" => data_out <= rom_array(10572);
		when "0010100101001101" => data_out <= rom_array(10573);
		when "0010100101001110" => data_out <= rom_array(10574);
		when "0010100101001111" => data_out <= rom_array(10575);
		when "0010100101010000" => data_out <= rom_array(10576);
		when "0010100101010001" => data_out <= rom_array(10577);
		when "0010100101010010" => data_out <= rom_array(10578);
		when "0010100101010011" => data_out <= rom_array(10579);
		when "0010100101010100" => data_out <= rom_array(10580);
		when "0010100101010101" => data_out <= rom_array(10581);
		when "0010100101010110" => data_out <= rom_array(10582);
		when "0010100101010111" => data_out <= rom_array(10583);
		when "0010100101011000" => data_out <= rom_array(10584);
		when "0010100101011001" => data_out <= rom_array(10585);
		when "0010100101011010" => data_out <= rom_array(10586);
		when "0010100101011011" => data_out <= rom_array(10587);
		when "0010100101011100" => data_out <= rom_array(10588);
		when "0010100101011101" => data_out <= rom_array(10589);
		when "0010100101011110" => data_out <= rom_array(10590);
		when "0010100101011111" => data_out <= rom_array(10591);
		when "0010100101100000" => data_out <= rom_array(10592);
		when "0010100101100001" => data_out <= rom_array(10593);
		when "0010100101100010" => data_out <= rom_array(10594);
		when "0010100101100011" => data_out <= rom_array(10595);
		when "0010100101100100" => data_out <= rom_array(10596);
		when "0010100101100101" => data_out <= rom_array(10597);
		when "0010100101100110" => data_out <= rom_array(10598);
		when "0010100101100111" => data_out <= rom_array(10599);
		when "0010100101101000" => data_out <= rom_array(10600);
		when "0010100101101001" => data_out <= rom_array(10601);
		when "0010100101101010" => data_out <= rom_array(10602);
		when "0010100101101011" => data_out <= rom_array(10603);
		when "0010100101101100" => data_out <= rom_array(10604);
		when "0010100101101101" => data_out <= rom_array(10605);
		when "0010100101101110" => data_out <= rom_array(10606);
		when "0010100101101111" => data_out <= rom_array(10607);
		when "0010100101110000" => data_out <= rom_array(10608);
		when "0010100101110001" => data_out <= rom_array(10609);
		when "0010100101110010" => data_out <= rom_array(10610);
		when "0010100101110011" => data_out <= rom_array(10611);
		when "0010100101110100" => data_out <= rom_array(10612);
		when "0010100101110101" => data_out <= rom_array(10613);
		when "0010100101110110" => data_out <= rom_array(10614);
		when "0010100101110111" => data_out <= rom_array(10615);
		when "0010100101111000" => data_out <= rom_array(10616);
		when "0010100101111001" => data_out <= rom_array(10617);
		when "0010100101111010" => data_out <= rom_array(10618);
		when "0010100101111011" => data_out <= rom_array(10619);
		when "0010100101111100" => data_out <= rom_array(10620);
		when "0010100101111101" => data_out <= rom_array(10621);
		when "0010100101111110" => data_out <= rom_array(10622);
		when "0010100101111111" => data_out <= rom_array(10623);
		when "0010100110000000" => data_out <= rom_array(10624);
		when "0010100110000001" => data_out <= rom_array(10625);
		when "0010100110000010" => data_out <= rom_array(10626);
		when "0010100110000011" => data_out <= rom_array(10627);
		when "0010100110000100" => data_out <= rom_array(10628);
		when "0010100110000101" => data_out <= rom_array(10629);
		when "0010100110000110" => data_out <= rom_array(10630);
		when "0010100110000111" => data_out <= rom_array(10631);
		when "0010100110001000" => data_out <= rom_array(10632);
		when "0010100110001001" => data_out <= rom_array(10633);
		when "0010100110001010" => data_out <= rom_array(10634);
		when "0010100110001011" => data_out <= rom_array(10635);
		when "0010100110001100" => data_out <= rom_array(10636);
		when "0010100110001101" => data_out <= rom_array(10637);
		when "0010100110001110" => data_out <= rom_array(10638);
		when "0010100110001111" => data_out <= rom_array(10639);
		when "0010100110010000" => data_out <= rom_array(10640);
		when "0010100110010001" => data_out <= rom_array(10641);
		when "0010100110010010" => data_out <= rom_array(10642);
		when "0010100110010011" => data_out <= rom_array(10643);
		when "0010100110010100" => data_out <= rom_array(10644);
		when "0010100110010101" => data_out <= rom_array(10645);
		when "0010100110010110" => data_out <= rom_array(10646);
		when "0010100110010111" => data_out <= rom_array(10647);
		when "0010100110011000" => data_out <= rom_array(10648);
		when "0010100110011001" => data_out <= rom_array(10649);
		when "0010100110011010" => data_out <= rom_array(10650);
		when "0010100110011011" => data_out <= rom_array(10651);
		when "0010100110011100" => data_out <= rom_array(10652);
		when "0010100110011101" => data_out <= rom_array(10653);
		when "0010100110011110" => data_out <= rom_array(10654);
		when "0010100110011111" => data_out <= rom_array(10655);
		when "0010100110100000" => data_out <= rom_array(10656);
		when "0010100110100001" => data_out <= rom_array(10657);
		when "0010100110100010" => data_out <= rom_array(10658);
		when "0010100110100011" => data_out <= rom_array(10659);
		when "0010100110100100" => data_out <= rom_array(10660);
		when "0010100110100101" => data_out <= rom_array(10661);
		when "0010100110100110" => data_out <= rom_array(10662);
		when "0010100110100111" => data_out <= rom_array(10663);
		when "0010100110101000" => data_out <= rom_array(10664);
		when "0010100110101001" => data_out <= rom_array(10665);
		when "0010100110101010" => data_out <= rom_array(10666);
		when "0010100110101011" => data_out <= rom_array(10667);
		when "0010100110101100" => data_out <= rom_array(10668);
		when "0010100110101101" => data_out <= rom_array(10669);
		when "0010100110101110" => data_out <= rom_array(10670);
		when "0010100110101111" => data_out <= rom_array(10671);
		when "0010100110110000" => data_out <= rom_array(10672);
		when "0010100110110001" => data_out <= rom_array(10673);
		when "0010100110110010" => data_out <= rom_array(10674);
		when "0010100110110011" => data_out <= rom_array(10675);
		when "0010100110110100" => data_out <= rom_array(10676);
		when "0010100110110101" => data_out <= rom_array(10677);
		when "0010100110110110" => data_out <= rom_array(10678);
		when "0010100110110111" => data_out <= rom_array(10679);
		when "0010100110111000" => data_out <= rom_array(10680);
		when "0010100110111001" => data_out <= rom_array(10681);
		when "0010100110111010" => data_out <= rom_array(10682);
		when "0010100110111011" => data_out <= rom_array(10683);
		when "0010100110111100" => data_out <= rom_array(10684);
		when "0010100110111101" => data_out <= rom_array(10685);
		when "0010100110111110" => data_out <= rom_array(10686);
		when "0010100110111111" => data_out <= rom_array(10687);
		when "0010100111000000" => data_out <= rom_array(10688);
		when "0010100111000001" => data_out <= rom_array(10689);
		when "0010100111000010" => data_out <= rom_array(10690);
		when "0010100111000011" => data_out <= rom_array(10691);
		when "0010100111000100" => data_out <= rom_array(10692);
		when "0010100111000101" => data_out <= rom_array(10693);
		when "0010100111000110" => data_out <= rom_array(10694);
		when "0010100111000111" => data_out <= rom_array(10695);
		when "0010100111001000" => data_out <= rom_array(10696);
		when "0010100111001001" => data_out <= rom_array(10697);
		when "0010100111001010" => data_out <= rom_array(10698);
		when "0010100111001011" => data_out <= rom_array(10699);
		when "0010100111001100" => data_out <= rom_array(10700);
		when "0010100111001101" => data_out <= rom_array(10701);
		when "0010100111001110" => data_out <= rom_array(10702);
		when "0010100111001111" => data_out <= rom_array(10703);
		when "0010100111010000" => data_out <= rom_array(10704);
		when "0010100111010001" => data_out <= rom_array(10705);
		when "0010100111010010" => data_out <= rom_array(10706);
		when "0010100111010011" => data_out <= rom_array(10707);
		when "0010100111010100" => data_out <= rom_array(10708);
		when "0010100111010101" => data_out <= rom_array(10709);
		when "0010100111010110" => data_out <= rom_array(10710);
		when "0010100111010111" => data_out <= rom_array(10711);
		when "0010100111011000" => data_out <= rom_array(10712);
		when "0010100111011001" => data_out <= rom_array(10713);
		when "0010100111011010" => data_out <= rom_array(10714);
		when "0010100111011011" => data_out <= rom_array(10715);
		when "0010100111011100" => data_out <= rom_array(10716);
		when "0010100111011101" => data_out <= rom_array(10717);
		when "0010100111011110" => data_out <= rom_array(10718);
		when "0010100111011111" => data_out <= rom_array(10719);
		when "0010100111100000" => data_out <= rom_array(10720);
		when "0010100111100001" => data_out <= rom_array(10721);
		when "0010100111100010" => data_out <= rom_array(10722);
		when "0010100111100011" => data_out <= rom_array(10723);
		when "0010100111100100" => data_out <= rom_array(10724);
		when "0010100111100101" => data_out <= rom_array(10725);
		when "0010100111100110" => data_out <= rom_array(10726);
		when "0010100111100111" => data_out <= rom_array(10727);
		when "0010100111101000" => data_out <= rom_array(10728);
		when "0010100111101001" => data_out <= rom_array(10729);
		when "0010100111101010" => data_out <= rom_array(10730);
		when "0010100111101011" => data_out <= rom_array(10731);
		when "0010100111101100" => data_out <= rom_array(10732);
		when "0010100111101101" => data_out <= rom_array(10733);
		when "0010100111101110" => data_out <= rom_array(10734);
		when "0010100111101111" => data_out <= rom_array(10735);
		when "0010100111110000" => data_out <= rom_array(10736);
		when "0010100111110001" => data_out <= rom_array(10737);
		when "0010100111110010" => data_out <= rom_array(10738);
		when "0010100111110011" => data_out <= rom_array(10739);
		when "0010100111110100" => data_out <= rom_array(10740);
		when "0010100111110101" => data_out <= rom_array(10741);
		when "0010100111110110" => data_out <= rom_array(10742);
		when "0010100111110111" => data_out <= rom_array(10743);
		when "0010100111111000" => data_out <= rom_array(10744);
		when "0010100111111001" => data_out <= rom_array(10745);
		when "0010100111111010" => data_out <= rom_array(10746);
		when "0010100111111011" => data_out <= rom_array(10747);
		when "0010100111111100" => data_out <= rom_array(10748);
		when "0010100111111101" => data_out <= rom_array(10749);
		when "0010100111111110" => data_out <= rom_array(10750);
		when "0010100111111111" => data_out <= rom_array(10751);
		when "0010101000000000" => data_out <= rom_array(10752);
		when "0010101000000001" => data_out <= rom_array(10753);
		when "0010101000000010" => data_out <= rom_array(10754);
		when "0010101000000011" => data_out <= rom_array(10755);
		when "0010101000000100" => data_out <= rom_array(10756);
		when "0010101000000101" => data_out <= rom_array(10757);
		when "0010101000000110" => data_out <= rom_array(10758);
		when "0010101000000111" => data_out <= rom_array(10759);
		when "0010101000001000" => data_out <= rom_array(10760);
		when "0010101000001001" => data_out <= rom_array(10761);
		when "0010101000001010" => data_out <= rom_array(10762);
		when "0010101000001011" => data_out <= rom_array(10763);
		when "0010101000001100" => data_out <= rom_array(10764);
		when "0010101000001101" => data_out <= rom_array(10765);
		when "0010101000001110" => data_out <= rom_array(10766);
		when "0010101000001111" => data_out <= rom_array(10767);
		when "0010101000010000" => data_out <= rom_array(10768);
		when "0010101000010001" => data_out <= rom_array(10769);
		when "0010101000010010" => data_out <= rom_array(10770);
		when "0010101000010011" => data_out <= rom_array(10771);
		when "0010101000010100" => data_out <= rom_array(10772);
		when "0010101000010101" => data_out <= rom_array(10773);
		when "0010101000010110" => data_out <= rom_array(10774);
		when "0010101000010111" => data_out <= rom_array(10775);
		when "0010101000011000" => data_out <= rom_array(10776);
		when "0010101000011001" => data_out <= rom_array(10777);
		when "0010101000011010" => data_out <= rom_array(10778);
		when "0010101000011011" => data_out <= rom_array(10779);
		when "0010101000011100" => data_out <= rom_array(10780);
		when "0010101000011101" => data_out <= rom_array(10781);
		when "0010101000011110" => data_out <= rom_array(10782);
		when "0010101000011111" => data_out <= rom_array(10783);
		when "0010101000100000" => data_out <= rom_array(10784);
		when "0010101000100001" => data_out <= rom_array(10785);
		when "0010101000100010" => data_out <= rom_array(10786);
		when "0010101000100011" => data_out <= rom_array(10787);
		when "0010101000100100" => data_out <= rom_array(10788);
		when "0010101000100101" => data_out <= rom_array(10789);
		when "0010101000100110" => data_out <= rom_array(10790);
		when "0010101000100111" => data_out <= rom_array(10791);
		when "0010101000101000" => data_out <= rom_array(10792);
		when "0010101000101001" => data_out <= rom_array(10793);
		when "0010101000101010" => data_out <= rom_array(10794);
		when "0010101000101011" => data_out <= rom_array(10795);
		when "0010101000101100" => data_out <= rom_array(10796);
		when "0010101000101101" => data_out <= rom_array(10797);
		when "0010101000101110" => data_out <= rom_array(10798);
		when "0010101000101111" => data_out <= rom_array(10799);
		when "0010101000110000" => data_out <= rom_array(10800);
		when "0010101000110001" => data_out <= rom_array(10801);
		when "0010101000110010" => data_out <= rom_array(10802);
		when "0010101000110011" => data_out <= rom_array(10803);
		when "0010101000110100" => data_out <= rom_array(10804);
		when "0010101000110101" => data_out <= rom_array(10805);
		when "0010101000110110" => data_out <= rom_array(10806);
		when "0010101000110111" => data_out <= rom_array(10807);
		when "0010101000111000" => data_out <= rom_array(10808);
		when "0010101000111001" => data_out <= rom_array(10809);
		when "0010101000111010" => data_out <= rom_array(10810);
		when "0010101000111011" => data_out <= rom_array(10811);
		when "0010101000111100" => data_out <= rom_array(10812);
		when "0010101000111101" => data_out <= rom_array(10813);
		when "0010101000111110" => data_out <= rom_array(10814);
		when "0010101000111111" => data_out <= rom_array(10815);
		when "0010101001000000" => data_out <= rom_array(10816);
		when "0010101001000001" => data_out <= rom_array(10817);
		when "0010101001000010" => data_out <= rom_array(10818);
		when "0010101001000011" => data_out <= rom_array(10819);
		when "0010101001000100" => data_out <= rom_array(10820);
		when "0010101001000101" => data_out <= rom_array(10821);
		when "0010101001000110" => data_out <= rom_array(10822);
		when "0010101001000111" => data_out <= rom_array(10823);
		when "0010101001001000" => data_out <= rom_array(10824);
		when "0010101001001001" => data_out <= rom_array(10825);
		when "0010101001001010" => data_out <= rom_array(10826);
		when "0010101001001011" => data_out <= rom_array(10827);
		when "0010101001001100" => data_out <= rom_array(10828);
		when "0010101001001101" => data_out <= rom_array(10829);
		when "0010101001001110" => data_out <= rom_array(10830);
		when "0010101001001111" => data_out <= rom_array(10831);
		when "0010101001010000" => data_out <= rom_array(10832);
		when "0010101001010001" => data_out <= rom_array(10833);
		when "0010101001010010" => data_out <= rom_array(10834);
		when "0010101001010011" => data_out <= rom_array(10835);
		when "0010101001010100" => data_out <= rom_array(10836);
		when "0010101001010101" => data_out <= rom_array(10837);
		when "0010101001010110" => data_out <= rom_array(10838);
		when "0010101001010111" => data_out <= rom_array(10839);
		when "0010101001011000" => data_out <= rom_array(10840);
		when "0010101001011001" => data_out <= rom_array(10841);
		when "0010101001011010" => data_out <= rom_array(10842);
		when "0010101001011011" => data_out <= rom_array(10843);
		when "0010101001011100" => data_out <= rom_array(10844);
		when "0010101001011101" => data_out <= rom_array(10845);
		when "0010101001011110" => data_out <= rom_array(10846);
		when "0010101001011111" => data_out <= rom_array(10847);
		when "0010101001100000" => data_out <= rom_array(10848);
		when "0010101001100001" => data_out <= rom_array(10849);
		when "0010101001100010" => data_out <= rom_array(10850);
		when "0010101001100011" => data_out <= rom_array(10851);
		when "0010101001100100" => data_out <= rom_array(10852);
		when "0010101001100101" => data_out <= rom_array(10853);
		when "0010101001100110" => data_out <= rom_array(10854);
		when "0010101001100111" => data_out <= rom_array(10855);
		when "0010101001101000" => data_out <= rom_array(10856);
		when "0010101001101001" => data_out <= rom_array(10857);
		when "0010101001101010" => data_out <= rom_array(10858);
		when "0010101001101011" => data_out <= rom_array(10859);
		when "0010101001101100" => data_out <= rom_array(10860);
		when "0010101001101101" => data_out <= rom_array(10861);
		when "0010101001101110" => data_out <= rom_array(10862);
		when "0010101001101111" => data_out <= rom_array(10863);
		when "0010101001110000" => data_out <= rom_array(10864);
		when "0010101001110001" => data_out <= rom_array(10865);
		when "0010101001110010" => data_out <= rom_array(10866);
		when "0010101001110011" => data_out <= rom_array(10867);
		when "0010101001110100" => data_out <= rom_array(10868);
		when "0010101001110101" => data_out <= rom_array(10869);
		when "0010101001110110" => data_out <= rom_array(10870);
		when "0010101001110111" => data_out <= rom_array(10871);
		when "0010101001111000" => data_out <= rom_array(10872);
		when "0010101001111001" => data_out <= rom_array(10873);
		when "0010101001111010" => data_out <= rom_array(10874);
		when "0010101001111011" => data_out <= rom_array(10875);
		when "0010101001111100" => data_out <= rom_array(10876);
		when "0010101001111101" => data_out <= rom_array(10877);
		when "0010101001111110" => data_out <= rom_array(10878);
		when "0010101001111111" => data_out <= rom_array(10879);
		when "0010101010000000" => data_out <= rom_array(10880);
		when "0010101010000001" => data_out <= rom_array(10881);
		when "0010101010000010" => data_out <= rom_array(10882);
		when "0010101010000011" => data_out <= rom_array(10883);
		when "0010101010000100" => data_out <= rom_array(10884);
		when "0010101010000101" => data_out <= rom_array(10885);
		when "0010101010000110" => data_out <= rom_array(10886);
		when "0010101010000111" => data_out <= rom_array(10887);
		when "0010101010001000" => data_out <= rom_array(10888);
		when "0010101010001001" => data_out <= rom_array(10889);
		when "0010101010001010" => data_out <= rom_array(10890);
		when "0010101010001011" => data_out <= rom_array(10891);
		when "0010101010001100" => data_out <= rom_array(10892);
		when "0010101010001101" => data_out <= rom_array(10893);
		when "0010101010001110" => data_out <= rom_array(10894);
		when "0010101010001111" => data_out <= rom_array(10895);
		when "0010101010010000" => data_out <= rom_array(10896);
		when "0010101010010001" => data_out <= rom_array(10897);
		when "0010101010010010" => data_out <= rom_array(10898);
		when "0010101010010011" => data_out <= rom_array(10899);
		when "0010101010010100" => data_out <= rom_array(10900);
		when "0010101010010101" => data_out <= rom_array(10901);
		when "0010101010010110" => data_out <= rom_array(10902);
		when "0010101010010111" => data_out <= rom_array(10903);
		when "0010101010011000" => data_out <= rom_array(10904);
		when "0010101010011001" => data_out <= rom_array(10905);
		when "0010101010011010" => data_out <= rom_array(10906);
		when "0010101010011011" => data_out <= rom_array(10907);
		when "0010101010011100" => data_out <= rom_array(10908);
		when "0010101010011101" => data_out <= rom_array(10909);
		when "0010101010011110" => data_out <= rom_array(10910);
		when "0010101010011111" => data_out <= rom_array(10911);
		when "0010101010100000" => data_out <= rom_array(10912);
		when "0010101010100001" => data_out <= rom_array(10913);
		when "0010101010100010" => data_out <= rom_array(10914);
		when "0010101010100011" => data_out <= rom_array(10915);
		when "0010101010100100" => data_out <= rom_array(10916);
		when "0010101010100101" => data_out <= rom_array(10917);
		when "0010101010100110" => data_out <= rom_array(10918);
		when "0010101010100111" => data_out <= rom_array(10919);
		when "0010101010101000" => data_out <= rom_array(10920);
		when "0010101010101001" => data_out <= rom_array(10921);
		when "0010101010101010" => data_out <= rom_array(10922);
		when "0010101010101011" => data_out <= rom_array(10923);
		when "0010101010101100" => data_out <= rom_array(10924);
		when "0010101010101101" => data_out <= rom_array(10925);
		when "0010101010101110" => data_out <= rom_array(10926);
		when "0010101010101111" => data_out <= rom_array(10927);
		when "0010101010110000" => data_out <= rom_array(10928);
		when "0010101010110001" => data_out <= rom_array(10929);
		when "0010101010110010" => data_out <= rom_array(10930);
		when "0010101010110011" => data_out <= rom_array(10931);
		when "0010101010110100" => data_out <= rom_array(10932);
		when "0010101010110101" => data_out <= rom_array(10933);
		when "0010101010110110" => data_out <= rom_array(10934);
		when "0010101010110111" => data_out <= rom_array(10935);
		when "0010101010111000" => data_out <= rom_array(10936);
		when "0010101010111001" => data_out <= rom_array(10937);
		when "0010101010111010" => data_out <= rom_array(10938);
		when "0010101010111011" => data_out <= rom_array(10939);
		when "0010101010111100" => data_out <= rom_array(10940);
		when "0010101010111101" => data_out <= rom_array(10941);
		when "0010101010111110" => data_out <= rom_array(10942);
		when "0010101010111111" => data_out <= rom_array(10943);
		when "0010101011000000" => data_out <= rom_array(10944);
		when "0010101011000001" => data_out <= rom_array(10945);
		when "0010101011000010" => data_out <= rom_array(10946);
		when "0010101011000011" => data_out <= rom_array(10947);
		when "0010101011000100" => data_out <= rom_array(10948);
		when "0010101011000101" => data_out <= rom_array(10949);
		when "0010101011000110" => data_out <= rom_array(10950);
		when "0010101011000111" => data_out <= rom_array(10951);
		when "0010101011001000" => data_out <= rom_array(10952);
		when "0010101011001001" => data_out <= rom_array(10953);
		when "0010101011001010" => data_out <= rom_array(10954);
		when "0010101011001011" => data_out <= rom_array(10955);
		when "0010101011001100" => data_out <= rom_array(10956);
		when "0010101011001101" => data_out <= rom_array(10957);
		when "0010101011001110" => data_out <= rom_array(10958);
		when "0010101011001111" => data_out <= rom_array(10959);
		when "0010101011010000" => data_out <= rom_array(10960);
		when "0010101011010001" => data_out <= rom_array(10961);
		when "0010101011010010" => data_out <= rom_array(10962);
		when "0010101011010011" => data_out <= rom_array(10963);
		when "0010101011010100" => data_out <= rom_array(10964);
		when "0010101011010101" => data_out <= rom_array(10965);
		when "0010101011010110" => data_out <= rom_array(10966);
		when "0010101011010111" => data_out <= rom_array(10967);
		when "0010101011011000" => data_out <= rom_array(10968);
		when "0010101011011001" => data_out <= rom_array(10969);
		when "0010101011011010" => data_out <= rom_array(10970);
		when "0010101011011011" => data_out <= rom_array(10971);
		when "0010101011011100" => data_out <= rom_array(10972);
		when "0010101011011101" => data_out <= rom_array(10973);
		when "0010101011011110" => data_out <= rom_array(10974);
		when "0010101011011111" => data_out <= rom_array(10975);
		when "0010101011100000" => data_out <= rom_array(10976);
		when "0010101011100001" => data_out <= rom_array(10977);
		when "0010101011100010" => data_out <= rom_array(10978);
		when "0010101011100011" => data_out <= rom_array(10979);
		when "0010101011100100" => data_out <= rom_array(10980);
		when "0010101011100101" => data_out <= rom_array(10981);
		when "0010101011100110" => data_out <= rom_array(10982);
		when "0010101011100111" => data_out <= rom_array(10983);
		when "0010101011101000" => data_out <= rom_array(10984);
		when "0010101011101001" => data_out <= rom_array(10985);
		when "0010101011101010" => data_out <= rom_array(10986);
		when "0010101011101011" => data_out <= rom_array(10987);
		when "0010101011101100" => data_out <= rom_array(10988);
		when "0010101011101101" => data_out <= rom_array(10989);
		when "0010101011101110" => data_out <= rom_array(10990);
		when "0010101011101111" => data_out <= rom_array(10991);
		when "0010101011110000" => data_out <= rom_array(10992);
		when "0010101011110001" => data_out <= rom_array(10993);
		when "0010101011110010" => data_out <= rom_array(10994);
		when "0010101011110011" => data_out <= rom_array(10995);
		when "0010101011110100" => data_out <= rom_array(10996);
		when "0010101011110101" => data_out <= rom_array(10997);
		when "0010101011110110" => data_out <= rom_array(10998);
		when "0010101011110111" => data_out <= rom_array(10999);
		when "0010101011111000" => data_out <= rom_array(11000);
		when "0010101011111001" => data_out <= rom_array(11001);
		when "0010101011111010" => data_out <= rom_array(11002);
		when "0010101011111011" => data_out <= rom_array(11003);
		when "0010101011111100" => data_out <= rom_array(11004);
		when "0010101011111101" => data_out <= rom_array(11005);
		when "0010101011111110" => data_out <= rom_array(11006);
		when "0010101011111111" => data_out <= rom_array(11007);
		when "0010101100000000" => data_out <= rom_array(11008);
		when "0010101100000001" => data_out <= rom_array(11009);
		when "0010101100000010" => data_out <= rom_array(11010);
		when "0010101100000011" => data_out <= rom_array(11011);
		when "0010101100000100" => data_out <= rom_array(11012);
		when "0010101100000101" => data_out <= rom_array(11013);
		when "0010101100000110" => data_out <= rom_array(11014);
		when "0010101100000111" => data_out <= rom_array(11015);
		when "0010101100001000" => data_out <= rom_array(11016);
		when "0010101100001001" => data_out <= rom_array(11017);
		when "0010101100001010" => data_out <= rom_array(11018);
		when "0010101100001011" => data_out <= rom_array(11019);
		when "0010101100001100" => data_out <= rom_array(11020);
		when "0010101100001101" => data_out <= rom_array(11021);
		when "0010101100001110" => data_out <= rom_array(11022);
		when "0010101100001111" => data_out <= rom_array(11023);
		when "0010101100010000" => data_out <= rom_array(11024);
		when "0010101100010001" => data_out <= rom_array(11025);
		when "0010101100010010" => data_out <= rom_array(11026);
		when "0010101100010011" => data_out <= rom_array(11027);
		when "0010101100010100" => data_out <= rom_array(11028);
		when "0010101100010101" => data_out <= rom_array(11029);
		when "0010101100010110" => data_out <= rom_array(11030);
		when "0010101100010111" => data_out <= rom_array(11031);
		when "0010101100011000" => data_out <= rom_array(11032);
		when "0010101100011001" => data_out <= rom_array(11033);
		when "0010101100011010" => data_out <= rom_array(11034);
		when "0010101100011011" => data_out <= rom_array(11035);
		when "0010101100011100" => data_out <= rom_array(11036);
		when "0010101100011101" => data_out <= rom_array(11037);
		when "0010101100011110" => data_out <= rom_array(11038);
		when "0010101100011111" => data_out <= rom_array(11039);
		when "0010101100100000" => data_out <= rom_array(11040);
		when "0010101100100001" => data_out <= rom_array(11041);
		when "0010101100100010" => data_out <= rom_array(11042);
		when "0010101100100011" => data_out <= rom_array(11043);
		when "0010101100100100" => data_out <= rom_array(11044);
		when "0010101100100101" => data_out <= rom_array(11045);
		when "0010101100100110" => data_out <= rom_array(11046);
		when "0010101100100111" => data_out <= rom_array(11047);
		when "0010101100101000" => data_out <= rom_array(11048);
		when "0010101100101001" => data_out <= rom_array(11049);
		when "0010101100101010" => data_out <= rom_array(11050);
		when "0010101100101011" => data_out <= rom_array(11051);
		when "0010101100101100" => data_out <= rom_array(11052);
		when "0010101100101101" => data_out <= rom_array(11053);
		when "0010101100101110" => data_out <= rom_array(11054);
		when "0010101100101111" => data_out <= rom_array(11055);
		when "0010101100110000" => data_out <= rom_array(11056);
		when "0010101100110001" => data_out <= rom_array(11057);
		when "0010101100110010" => data_out <= rom_array(11058);
		when "0010101100110011" => data_out <= rom_array(11059);
		when "0010101100110100" => data_out <= rom_array(11060);
		when "0010101100110101" => data_out <= rom_array(11061);
		when "0010101100110110" => data_out <= rom_array(11062);
		when "0010101100110111" => data_out <= rom_array(11063);
		when "0010101100111000" => data_out <= rom_array(11064);
		when "0010101100111001" => data_out <= rom_array(11065);
		when "0010101100111010" => data_out <= rom_array(11066);
		when "0010101100111011" => data_out <= rom_array(11067);
		when "0010101100111100" => data_out <= rom_array(11068);
		when "0010101100111101" => data_out <= rom_array(11069);
		when "0010101100111110" => data_out <= rom_array(11070);
		when "0010101100111111" => data_out <= rom_array(11071);
		when "0010101101000000" => data_out <= rom_array(11072);
		when "0010101101000001" => data_out <= rom_array(11073);
		when "0010101101000010" => data_out <= rom_array(11074);
		when "0010101101000011" => data_out <= rom_array(11075);
		when "0010101101000100" => data_out <= rom_array(11076);
		when "0010101101000101" => data_out <= rom_array(11077);
		when "0010101101000110" => data_out <= rom_array(11078);
		when "0010101101000111" => data_out <= rom_array(11079);
		when "0010101101001000" => data_out <= rom_array(11080);
		when "0010101101001001" => data_out <= rom_array(11081);
		when "0010101101001010" => data_out <= rom_array(11082);
		when "0010101101001011" => data_out <= rom_array(11083);
		when "0010101101001100" => data_out <= rom_array(11084);
		when "0010101101001101" => data_out <= rom_array(11085);
		when "0010101101001110" => data_out <= rom_array(11086);
		when "0010101101001111" => data_out <= rom_array(11087);
		when "0010101101010000" => data_out <= rom_array(11088);
		when "0010101101010001" => data_out <= rom_array(11089);
		when "0010101101010010" => data_out <= rom_array(11090);
		when "0010101101010011" => data_out <= rom_array(11091);
		when "0010101101010100" => data_out <= rom_array(11092);
		when "0010101101010101" => data_out <= rom_array(11093);
		when "0010101101010110" => data_out <= rom_array(11094);
		when "0010101101010111" => data_out <= rom_array(11095);
		when "0010101101011000" => data_out <= rom_array(11096);
		when "0010101101011001" => data_out <= rom_array(11097);
		when "0010101101011010" => data_out <= rom_array(11098);
		when "0010101101011011" => data_out <= rom_array(11099);
		when "0010101101011100" => data_out <= rom_array(11100);
		when "0010101101011101" => data_out <= rom_array(11101);
		when "0010101101011110" => data_out <= rom_array(11102);
		when "0010101101011111" => data_out <= rom_array(11103);
		when "0010101101100000" => data_out <= rom_array(11104);
		when "0010101101100001" => data_out <= rom_array(11105);
		when "0010101101100010" => data_out <= rom_array(11106);
		when "0010101101100011" => data_out <= rom_array(11107);
		when "0010101101100100" => data_out <= rom_array(11108);
		when "0010101101100101" => data_out <= rom_array(11109);
		when "0010101101100110" => data_out <= rom_array(11110);
		when "0010101101100111" => data_out <= rom_array(11111);
		when "0010101101101000" => data_out <= rom_array(11112);
		when "0010101101101001" => data_out <= rom_array(11113);
		when "0010101101101010" => data_out <= rom_array(11114);
		when "0010101101101011" => data_out <= rom_array(11115);
		when "0010101101101100" => data_out <= rom_array(11116);
		when "0010101101101101" => data_out <= rom_array(11117);
		when "0010101101101110" => data_out <= rom_array(11118);
		when "0010101101101111" => data_out <= rom_array(11119);
		when "0010101101110000" => data_out <= rom_array(11120);
		when "0010101101110001" => data_out <= rom_array(11121);
		when "0010101101110010" => data_out <= rom_array(11122);
		when "0010101101110011" => data_out <= rom_array(11123);
		when "0010101101110100" => data_out <= rom_array(11124);
		when "0010101101110101" => data_out <= rom_array(11125);
		when "0010101101110110" => data_out <= rom_array(11126);
		when "0010101101110111" => data_out <= rom_array(11127);
		when "0010101101111000" => data_out <= rom_array(11128);
		when "0010101101111001" => data_out <= rom_array(11129);
		when "0010101101111010" => data_out <= rom_array(11130);
		when "0010101101111011" => data_out <= rom_array(11131);
		when "0010101101111100" => data_out <= rom_array(11132);
		when "0010101101111101" => data_out <= rom_array(11133);
		when "0010101101111110" => data_out <= rom_array(11134);
		when "0010101101111111" => data_out <= rom_array(11135);
		when "0010101110000000" => data_out <= rom_array(11136);
		when "0010101110000001" => data_out <= rom_array(11137);
		when "0010101110000010" => data_out <= rom_array(11138);
		when "0010101110000011" => data_out <= rom_array(11139);
		when "0010101110000100" => data_out <= rom_array(11140);
		when "0010101110000101" => data_out <= rom_array(11141);
		when "0010101110000110" => data_out <= rom_array(11142);
		when "0010101110000111" => data_out <= rom_array(11143);
		when "0010101110001000" => data_out <= rom_array(11144);
		when "0010101110001001" => data_out <= rom_array(11145);
		when "0010101110001010" => data_out <= rom_array(11146);
		when "0010101110001011" => data_out <= rom_array(11147);
		when "0010101110001100" => data_out <= rom_array(11148);
		when "0010101110001101" => data_out <= rom_array(11149);
		when "0010101110001110" => data_out <= rom_array(11150);
		when "0010101110001111" => data_out <= rom_array(11151);
		when "0010101110010000" => data_out <= rom_array(11152);
		when "0010101110010001" => data_out <= rom_array(11153);
		when "0010101110010010" => data_out <= rom_array(11154);
		when "0010101110010011" => data_out <= rom_array(11155);
		when "0010101110010100" => data_out <= rom_array(11156);
		when "0010101110010101" => data_out <= rom_array(11157);
		when "0010101110010110" => data_out <= rom_array(11158);
		when "0010101110010111" => data_out <= rom_array(11159);
		when "0010101110011000" => data_out <= rom_array(11160);
		when "0010101110011001" => data_out <= rom_array(11161);
		when "0010101110011010" => data_out <= rom_array(11162);
		when "0010101110011011" => data_out <= rom_array(11163);
		when "0010101110011100" => data_out <= rom_array(11164);
		when "0010101110011101" => data_out <= rom_array(11165);
		when "0010101110011110" => data_out <= rom_array(11166);
		when "0010101110011111" => data_out <= rom_array(11167);
		when "0010101110100000" => data_out <= rom_array(11168);
		when "0010101110100001" => data_out <= rom_array(11169);
		when "0010101110100010" => data_out <= rom_array(11170);
		when "0010101110100011" => data_out <= rom_array(11171);
		when "0010101110100100" => data_out <= rom_array(11172);
		when "0010101110100101" => data_out <= rom_array(11173);
		when "0010101110100110" => data_out <= rom_array(11174);
		when "0010101110100111" => data_out <= rom_array(11175);
		when "0010101110101000" => data_out <= rom_array(11176);
		when "0010101110101001" => data_out <= rom_array(11177);
		when "0010101110101010" => data_out <= rom_array(11178);
		when "0010101110101011" => data_out <= rom_array(11179);
		when "0010101110101100" => data_out <= rom_array(11180);
		when "0010101110101101" => data_out <= rom_array(11181);
		when "0010101110101110" => data_out <= rom_array(11182);
		when "0010101110101111" => data_out <= rom_array(11183);
		when "0010101110110000" => data_out <= rom_array(11184);
		when "0010101110110001" => data_out <= rom_array(11185);
		when "0010101110110010" => data_out <= rom_array(11186);
		when "0010101110110011" => data_out <= rom_array(11187);
		when "0010101110110100" => data_out <= rom_array(11188);
		when "0010101110110101" => data_out <= rom_array(11189);
		when "0010101110110110" => data_out <= rom_array(11190);
		when "0010101110110111" => data_out <= rom_array(11191);
		when "0010101110111000" => data_out <= rom_array(11192);
		when "0010101110111001" => data_out <= rom_array(11193);
		when "0010101110111010" => data_out <= rom_array(11194);
		when "0010101110111011" => data_out <= rom_array(11195);
		when "0010101110111100" => data_out <= rom_array(11196);
		when "0010101110111101" => data_out <= rom_array(11197);
		when "0010101110111110" => data_out <= rom_array(11198);
		when "0010101110111111" => data_out <= rom_array(11199);
		when "0010101111000000" => data_out <= rom_array(11200);
		when "0010101111000001" => data_out <= rom_array(11201);
		when "0010101111000010" => data_out <= rom_array(11202);
		when "0010101111000011" => data_out <= rom_array(11203);
		when "0010101111000100" => data_out <= rom_array(11204);
		when "0010101111000101" => data_out <= rom_array(11205);
		when "0010101111000110" => data_out <= rom_array(11206);
		when "0010101111000111" => data_out <= rom_array(11207);
		when "0010101111001000" => data_out <= rom_array(11208);
		when "0010101111001001" => data_out <= rom_array(11209);
		when "0010101111001010" => data_out <= rom_array(11210);
		when "0010101111001011" => data_out <= rom_array(11211);
		when "0010101111001100" => data_out <= rom_array(11212);
		when "0010101111001101" => data_out <= rom_array(11213);
		when "0010101111001110" => data_out <= rom_array(11214);
		when "0010101111001111" => data_out <= rom_array(11215);
		when "0010101111010000" => data_out <= rom_array(11216);
		when "0010101111010001" => data_out <= rom_array(11217);
		when "0010101111010010" => data_out <= rom_array(11218);
		when "0010101111010011" => data_out <= rom_array(11219);
		when "0010101111010100" => data_out <= rom_array(11220);
		when "0010101111010101" => data_out <= rom_array(11221);
		when "0010101111010110" => data_out <= rom_array(11222);
		when "0010101111010111" => data_out <= rom_array(11223);
		when "0010101111011000" => data_out <= rom_array(11224);
		when "0010101111011001" => data_out <= rom_array(11225);
		when "0010101111011010" => data_out <= rom_array(11226);
		when "0010101111011011" => data_out <= rom_array(11227);
		when "0010101111011100" => data_out <= rom_array(11228);
		when "0010101111011101" => data_out <= rom_array(11229);
		when "0010101111011110" => data_out <= rom_array(11230);
		when "0010101111011111" => data_out <= rom_array(11231);
		when "0010101111100000" => data_out <= rom_array(11232);
		when "0010101111100001" => data_out <= rom_array(11233);
		when "0010101111100010" => data_out <= rom_array(11234);
		when "0010101111100011" => data_out <= rom_array(11235);
		when "0010101111100100" => data_out <= rom_array(11236);
		when "0010101111100101" => data_out <= rom_array(11237);
		when "0010101111100110" => data_out <= rom_array(11238);
		when "0010101111100111" => data_out <= rom_array(11239);
		when "0010101111101000" => data_out <= rom_array(11240);
		when "0010101111101001" => data_out <= rom_array(11241);
		when "0010101111101010" => data_out <= rom_array(11242);
		when "0010101111101011" => data_out <= rom_array(11243);
		when "0010101111101100" => data_out <= rom_array(11244);
		when "0010101111101101" => data_out <= rom_array(11245);
		when "0010101111101110" => data_out <= rom_array(11246);
		when "0010101111101111" => data_out <= rom_array(11247);
		when "0010101111110000" => data_out <= rom_array(11248);
		when "0010101111110001" => data_out <= rom_array(11249);
		when "0010101111110010" => data_out <= rom_array(11250);
		when "0010101111110011" => data_out <= rom_array(11251);
		when "0010101111110100" => data_out <= rom_array(11252);
		when "0010101111110101" => data_out <= rom_array(11253);
		when "0010101111110110" => data_out <= rom_array(11254);
		when "0010101111110111" => data_out <= rom_array(11255);
		when "0010101111111000" => data_out <= rom_array(11256);
		when "0010101111111001" => data_out <= rom_array(11257);
		when "0010101111111010" => data_out <= rom_array(11258);
		when "0010101111111011" => data_out <= rom_array(11259);
		when "0010101111111100" => data_out <= rom_array(11260);
		when "0010101111111101" => data_out <= rom_array(11261);
		when "0010101111111110" => data_out <= rom_array(11262);
		when "0010101111111111" => data_out <= rom_array(11263);
		when "0010110000000000" => data_out <= rom_array(11264);
		when "0010110000000001" => data_out <= rom_array(11265);
		when "0010110000000010" => data_out <= rom_array(11266);
		when "0010110000000011" => data_out <= rom_array(11267);
		when "0010110000000100" => data_out <= rom_array(11268);
		when "0010110000000101" => data_out <= rom_array(11269);
		when "0010110000000110" => data_out <= rom_array(11270);
		when "0010110000000111" => data_out <= rom_array(11271);
		when "0010110000001000" => data_out <= rom_array(11272);
		when "0010110000001001" => data_out <= rom_array(11273);
		when "0010110000001010" => data_out <= rom_array(11274);
		when "0010110000001011" => data_out <= rom_array(11275);
		when "0010110000001100" => data_out <= rom_array(11276);
		when "0010110000001101" => data_out <= rom_array(11277);
		when "0010110000001110" => data_out <= rom_array(11278);
		when "0010110000001111" => data_out <= rom_array(11279);
		when "0010110000010000" => data_out <= rom_array(11280);
		when "0010110000010001" => data_out <= rom_array(11281);
		when "0010110000010010" => data_out <= rom_array(11282);
		when "0010110000010011" => data_out <= rom_array(11283);
		when "0010110000010100" => data_out <= rom_array(11284);
		when "0010110000010101" => data_out <= rom_array(11285);
		when "0010110000010110" => data_out <= rom_array(11286);
		when "0010110000010111" => data_out <= rom_array(11287);
		when "0010110000011000" => data_out <= rom_array(11288);
		when "0010110000011001" => data_out <= rom_array(11289);
		when "0010110000011010" => data_out <= rom_array(11290);
		when "0010110000011011" => data_out <= rom_array(11291);
		when "0010110000011100" => data_out <= rom_array(11292);
		when "0010110000011101" => data_out <= rom_array(11293);
		when "0010110000011110" => data_out <= rom_array(11294);
		when "0010110000011111" => data_out <= rom_array(11295);
		when "0010110000100000" => data_out <= rom_array(11296);
		when "0010110000100001" => data_out <= rom_array(11297);
		when "0010110000100010" => data_out <= rom_array(11298);
		when "0010110000100011" => data_out <= rom_array(11299);
		when "0010110000100100" => data_out <= rom_array(11300);
		when "0010110000100101" => data_out <= rom_array(11301);
		when "0010110000100110" => data_out <= rom_array(11302);
		when "0010110000100111" => data_out <= rom_array(11303);
		when "0010110000101000" => data_out <= rom_array(11304);
		when "0010110000101001" => data_out <= rom_array(11305);
		when "0010110000101010" => data_out <= rom_array(11306);
		when "0010110000101011" => data_out <= rom_array(11307);
		when "0010110000101100" => data_out <= rom_array(11308);
		when "0010110000101101" => data_out <= rom_array(11309);
		when "0010110000101110" => data_out <= rom_array(11310);
		when "0010110000101111" => data_out <= rom_array(11311);
		when "0010110000110000" => data_out <= rom_array(11312);
		when "0010110000110001" => data_out <= rom_array(11313);
		when "0010110000110010" => data_out <= rom_array(11314);
		when "0010110000110011" => data_out <= rom_array(11315);
		when "0010110000110100" => data_out <= rom_array(11316);
		when "0010110000110101" => data_out <= rom_array(11317);
		when "0010110000110110" => data_out <= rom_array(11318);
		when "0010110000110111" => data_out <= rom_array(11319);
		when "0010110000111000" => data_out <= rom_array(11320);
		when "0010110000111001" => data_out <= rom_array(11321);
		when "0010110000111010" => data_out <= rom_array(11322);
		when "0010110000111011" => data_out <= rom_array(11323);
		when "0010110000111100" => data_out <= rom_array(11324);
		when "0010110000111101" => data_out <= rom_array(11325);
		when "0010110000111110" => data_out <= rom_array(11326);
		when "0010110000111111" => data_out <= rom_array(11327);
		when "0010110001000000" => data_out <= rom_array(11328);
		when "0010110001000001" => data_out <= rom_array(11329);
		when "0010110001000010" => data_out <= rom_array(11330);
		when "0010110001000011" => data_out <= rom_array(11331);
		when "0010110001000100" => data_out <= rom_array(11332);
		when "0010110001000101" => data_out <= rom_array(11333);
		when "0010110001000110" => data_out <= rom_array(11334);
		when "0010110001000111" => data_out <= rom_array(11335);
		when "0010110001001000" => data_out <= rom_array(11336);
		when "0010110001001001" => data_out <= rom_array(11337);
		when "0010110001001010" => data_out <= rom_array(11338);
		when "0010110001001011" => data_out <= rom_array(11339);
		when "0010110001001100" => data_out <= rom_array(11340);
		when "0010110001001101" => data_out <= rom_array(11341);
		when "0010110001001110" => data_out <= rom_array(11342);
		when "0010110001001111" => data_out <= rom_array(11343);
		when "0010110001010000" => data_out <= rom_array(11344);
		when "0010110001010001" => data_out <= rom_array(11345);
		when "0010110001010010" => data_out <= rom_array(11346);
		when "0010110001010011" => data_out <= rom_array(11347);
		when "0010110001010100" => data_out <= rom_array(11348);
		when "0010110001010101" => data_out <= rom_array(11349);
		when "0010110001010110" => data_out <= rom_array(11350);
		when "0010110001010111" => data_out <= rom_array(11351);
		when "0010110001011000" => data_out <= rom_array(11352);
		when "0010110001011001" => data_out <= rom_array(11353);
		when "0010110001011010" => data_out <= rom_array(11354);
		when "0010110001011011" => data_out <= rom_array(11355);
		when "0010110001011100" => data_out <= rom_array(11356);
		when "0010110001011101" => data_out <= rom_array(11357);
		when "0010110001011110" => data_out <= rom_array(11358);
		when "0010110001011111" => data_out <= rom_array(11359);
		when "0010110001100000" => data_out <= rom_array(11360);
		when "0010110001100001" => data_out <= rom_array(11361);
		when "0010110001100010" => data_out <= rom_array(11362);
		when "0010110001100011" => data_out <= rom_array(11363);
		when "0010110001100100" => data_out <= rom_array(11364);
		when "0010110001100101" => data_out <= rom_array(11365);
		when "0010110001100110" => data_out <= rom_array(11366);
		when "0010110001100111" => data_out <= rom_array(11367);
		when "0010110001101000" => data_out <= rom_array(11368);
		when "0010110001101001" => data_out <= rom_array(11369);
		when "0010110001101010" => data_out <= rom_array(11370);
		when "0010110001101011" => data_out <= rom_array(11371);
		when "0010110001101100" => data_out <= rom_array(11372);
		when "0010110001101101" => data_out <= rom_array(11373);
		when "0010110001101110" => data_out <= rom_array(11374);
		when "0010110001101111" => data_out <= rom_array(11375);
		when "0010110001110000" => data_out <= rom_array(11376);
		when "0010110001110001" => data_out <= rom_array(11377);
		when "0010110001110010" => data_out <= rom_array(11378);
		when "0010110001110011" => data_out <= rom_array(11379);
		when "0010110001110100" => data_out <= rom_array(11380);
		when "0010110001110101" => data_out <= rom_array(11381);
		when "0010110001110110" => data_out <= rom_array(11382);
		when "0010110001110111" => data_out <= rom_array(11383);
		when "0010110001111000" => data_out <= rom_array(11384);
		when "0010110001111001" => data_out <= rom_array(11385);
		when "0010110001111010" => data_out <= rom_array(11386);
		when "0010110001111011" => data_out <= rom_array(11387);
		when "0010110001111100" => data_out <= rom_array(11388);
		when "0010110001111101" => data_out <= rom_array(11389);
		when "0010110001111110" => data_out <= rom_array(11390);
		when "0010110001111111" => data_out <= rom_array(11391);
		when "0010110010000000" => data_out <= rom_array(11392);
		when "0010110010000001" => data_out <= rom_array(11393);
		when "0010110010000010" => data_out <= rom_array(11394);
		when "0010110010000011" => data_out <= rom_array(11395);
		when "0010110010000100" => data_out <= rom_array(11396);
		when "0010110010000101" => data_out <= rom_array(11397);
		when "0010110010000110" => data_out <= rom_array(11398);
		when "0010110010000111" => data_out <= rom_array(11399);
		when "0010110010001000" => data_out <= rom_array(11400);
		when "0010110010001001" => data_out <= rom_array(11401);
		when "0010110010001010" => data_out <= rom_array(11402);
		when "0010110010001011" => data_out <= rom_array(11403);
		when "0010110010001100" => data_out <= rom_array(11404);
		when "0010110010001101" => data_out <= rom_array(11405);
		when "0010110010001110" => data_out <= rom_array(11406);
		when "0010110010001111" => data_out <= rom_array(11407);
		when "0010110010010000" => data_out <= rom_array(11408);
		when "0010110010010001" => data_out <= rom_array(11409);
		when "0010110010010010" => data_out <= rom_array(11410);
		when "0010110010010011" => data_out <= rom_array(11411);
		when "0010110010010100" => data_out <= rom_array(11412);
		when "0010110010010101" => data_out <= rom_array(11413);
		when "0010110010010110" => data_out <= rom_array(11414);
		when "0010110010010111" => data_out <= rom_array(11415);
		when "0010110010011000" => data_out <= rom_array(11416);
		when "0010110010011001" => data_out <= rom_array(11417);
		when "0010110010011010" => data_out <= rom_array(11418);
		when "0010110010011011" => data_out <= rom_array(11419);
		when "0010110010011100" => data_out <= rom_array(11420);
		when "0010110010011101" => data_out <= rom_array(11421);
		when "0010110010011110" => data_out <= rom_array(11422);
		when "0010110010011111" => data_out <= rom_array(11423);
		when "0010110010100000" => data_out <= rom_array(11424);
		when "0010110010100001" => data_out <= rom_array(11425);
		when "0010110010100010" => data_out <= rom_array(11426);
		when "0010110010100011" => data_out <= rom_array(11427);
		when "0010110010100100" => data_out <= rom_array(11428);
		when "0010110010100101" => data_out <= rom_array(11429);
		when "0010110010100110" => data_out <= rom_array(11430);
		when "0010110010100111" => data_out <= rom_array(11431);
		when "0010110010101000" => data_out <= rom_array(11432);
		when "0010110010101001" => data_out <= rom_array(11433);
		when "0010110010101010" => data_out <= rom_array(11434);
		when "0010110010101011" => data_out <= rom_array(11435);
		when "0010110010101100" => data_out <= rom_array(11436);
		when "0010110010101101" => data_out <= rom_array(11437);
		when "0010110010101110" => data_out <= rom_array(11438);
		when "0010110010101111" => data_out <= rom_array(11439);
		when "0010110010110000" => data_out <= rom_array(11440);
		when "0010110010110001" => data_out <= rom_array(11441);
		when "0010110010110010" => data_out <= rom_array(11442);
		when "0010110010110011" => data_out <= rom_array(11443);
		when "0010110010110100" => data_out <= rom_array(11444);
		when "0010110010110101" => data_out <= rom_array(11445);
		when "0010110010110110" => data_out <= rom_array(11446);
		when "0010110010110111" => data_out <= rom_array(11447);
		when "0010110010111000" => data_out <= rom_array(11448);
		when "0010110010111001" => data_out <= rom_array(11449);
		when "0010110010111010" => data_out <= rom_array(11450);
		when "0010110010111011" => data_out <= rom_array(11451);
		when "0010110010111100" => data_out <= rom_array(11452);
		when "0010110010111101" => data_out <= rom_array(11453);
		when "0010110010111110" => data_out <= rom_array(11454);
		when "0010110010111111" => data_out <= rom_array(11455);
		when "0010110011000000" => data_out <= rom_array(11456);
		when "0010110011000001" => data_out <= rom_array(11457);
		when "0010110011000010" => data_out <= rom_array(11458);
		when "0010110011000011" => data_out <= rom_array(11459);
		when "0010110011000100" => data_out <= rom_array(11460);
		when "0010110011000101" => data_out <= rom_array(11461);
		when "0010110011000110" => data_out <= rom_array(11462);
		when "0010110011000111" => data_out <= rom_array(11463);
		when "0010110011001000" => data_out <= rom_array(11464);
		when "0010110011001001" => data_out <= rom_array(11465);
		when "0010110011001010" => data_out <= rom_array(11466);
		when "0010110011001011" => data_out <= rom_array(11467);
		when "0010110011001100" => data_out <= rom_array(11468);
		when "0010110011001101" => data_out <= rom_array(11469);
		when "0010110011001110" => data_out <= rom_array(11470);
		when "0010110011001111" => data_out <= rom_array(11471);
		when "0010110011010000" => data_out <= rom_array(11472);
		when "0010110011010001" => data_out <= rom_array(11473);
		when "0010110011010010" => data_out <= rom_array(11474);
		when "0010110011010011" => data_out <= rom_array(11475);
		when "0010110011010100" => data_out <= rom_array(11476);
		when "0010110011010101" => data_out <= rom_array(11477);
		when "0010110011010110" => data_out <= rom_array(11478);
		when "0010110011010111" => data_out <= rom_array(11479);
		when "0010110011011000" => data_out <= rom_array(11480);
		when "0010110011011001" => data_out <= rom_array(11481);
		when "0010110011011010" => data_out <= rom_array(11482);
		when "0010110011011011" => data_out <= rom_array(11483);
		when "0010110011011100" => data_out <= rom_array(11484);
		when "0010110011011101" => data_out <= rom_array(11485);
		when "0010110011011110" => data_out <= rom_array(11486);
		when "0010110011011111" => data_out <= rom_array(11487);
		when "0010110011100000" => data_out <= rom_array(11488);
		when "0010110011100001" => data_out <= rom_array(11489);
		when "0010110011100010" => data_out <= rom_array(11490);
		when "0010110011100011" => data_out <= rom_array(11491);
		when "0010110011100100" => data_out <= rom_array(11492);
		when "0010110011100101" => data_out <= rom_array(11493);
		when "0010110011100110" => data_out <= rom_array(11494);
		when "0010110011100111" => data_out <= rom_array(11495);
		when "0010110011101000" => data_out <= rom_array(11496);
		when "0010110011101001" => data_out <= rom_array(11497);
		when "0010110011101010" => data_out <= rom_array(11498);
		when "0010110011101011" => data_out <= rom_array(11499);
		when "0010110011101100" => data_out <= rom_array(11500);
		when "0010110011101101" => data_out <= rom_array(11501);
		when "0010110011101110" => data_out <= rom_array(11502);
		when "0010110011101111" => data_out <= rom_array(11503);
		when "0010110011110000" => data_out <= rom_array(11504);
		when "0010110011110001" => data_out <= rom_array(11505);
		when "0010110011110010" => data_out <= rom_array(11506);
		when "0010110011110011" => data_out <= rom_array(11507);
		when "0010110011110100" => data_out <= rom_array(11508);
		when "0010110011110101" => data_out <= rom_array(11509);
		when "0010110011110110" => data_out <= rom_array(11510);
		when "0010110011110111" => data_out <= rom_array(11511);
		when "0010110011111000" => data_out <= rom_array(11512);
		when "0010110011111001" => data_out <= rom_array(11513);
		when "0010110011111010" => data_out <= rom_array(11514);
		when "0010110011111011" => data_out <= rom_array(11515);
		when "0010110011111100" => data_out <= rom_array(11516);
		when "0010110011111101" => data_out <= rom_array(11517);
		when "0010110011111110" => data_out <= rom_array(11518);
		when "0010110011111111" => data_out <= rom_array(11519);
		when "0010110100000000" => data_out <= rom_array(11520);
		when "0010110100000001" => data_out <= rom_array(11521);
		when "0010110100000010" => data_out <= rom_array(11522);
		when "0010110100000011" => data_out <= rom_array(11523);
		when "0010110100000100" => data_out <= rom_array(11524);
		when "0010110100000101" => data_out <= rom_array(11525);
		when "0010110100000110" => data_out <= rom_array(11526);
		when "0010110100000111" => data_out <= rom_array(11527);
		when "0010110100001000" => data_out <= rom_array(11528);
		when "0010110100001001" => data_out <= rom_array(11529);
		when "0010110100001010" => data_out <= rom_array(11530);
		when "0010110100001011" => data_out <= rom_array(11531);
		when "0010110100001100" => data_out <= rom_array(11532);
		when "0010110100001101" => data_out <= rom_array(11533);
		when "0010110100001110" => data_out <= rom_array(11534);
		when "0010110100001111" => data_out <= rom_array(11535);
		when "0010110100010000" => data_out <= rom_array(11536);
		when "0010110100010001" => data_out <= rom_array(11537);
		when "0010110100010010" => data_out <= rom_array(11538);
		when "0010110100010011" => data_out <= rom_array(11539);
		when "0010110100010100" => data_out <= rom_array(11540);
		when "0010110100010101" => data_out <= rom_array(11541);
		when "0010110100010110" => data_out <= rom_array(11542);
		when "0010110100010111" => data_out <= rom_array(11543);
		when "0010110100011000" => data_out <= rom_array(11544);
		when "0010110100011001" => data_out <= rom_array(11545);
		when "0010110100011010" => data_out <= rom_array(11546);
		when "0010110100011011" => data_out <= rom_array(11547);
		when "0010110100011100" => data_out <= rom_array(11548);
		when "0010110100011101" => data_out <= rom_array(11549);
		when "0010110100011110" => data_out <= rom_array(11550);
		when "0010110100011111" => data_out <= rom_array(11551);
		when "0010110100100000" => data_out <= rom_array(11552);
		when "0010110100100001" => data_out <= rom_array(11553);
		when "0010110100100010" => data_out <= rom_array(11554);
		when "0010110100100011" => data_out <= rom_array(11555);
		when "0010110100100100" => data_out <= rom_array(11556);
		when "0010110100100101" => data_out <= rom_array(11557);
		when "0010110100100110" => data_out <= rom_array(11558);
		when "0010110100100111" => data_out <= rom_array(11559);
		when "0010110100101000" => data_out <= rom_array(11560);
		when "0010110100101001" => data_out <= rom_array(11561);
		when "0010110100101010" => data_out <= rom_array(11562);
		when "0010110100101011" => data_out <= rom_array(11563);
		when "0010110100101100" => data_out <= rom_array(11564);
		when "0010110100101101" => data_out <= rom_array(11565);
		when "0010110100101110" => data_out <= rom_array(11566);
		when "0010110100101111" => data_out <= rom_array(11567);
		when "0010110100110000" => data_out <= rom_array(11568);
		when "0010110100110001" => data_out <= rom_array(11569);
		when "0010110100110010" => data_out <= rom_array(11570);
		when "0010110100110011" => data_out <= rom_array(11571);
		when "0010110100110100" => data_out <= rom_array(11572);
		when "0010110100110101" => data_out <= rom_array(11573);
		when "0010110100110110" => data_out <= rom_array(11574);
		when "0010110100110111" => data_out <= rom_array(11575);
		when "0010110100111000" => data_out <= rom_array(11576);
		when "0010110100111001" => data_out <= rom_array(11577);
		when "0010110100111010" => data_out <= rom_array(11578);
		when "0010110100111011" => data_out <= rom_array(11579);
		when "0010110100111100" => data_out <= rom_array(11580);
		when "0010110100111101" => data_out <= rom_array(11581);
		when "0010110100111110" => data_out <= rom_array(11582);
		when "0010110100111111" => data_out <= rom_array(11583);
		when "0010110101000000" => data_out <= rom_array(11584);
		when "0010110101000001" => data_out <= rom_array(11585);
		when "0010110101000010" => data_out <= rom_array(11586);
		when "0010110101000011" => data_out <= rom_array(11587);
		when "0010110101000100" => data_out <= rom_array(11588);
		when "0010110101000101" => data_out <= rom_array(11589);
		when "0010110101000110" => data_out <= rom_array(11590);
		when "0010110101000111" => data_out <= rom_array(11591);
		when "0010110101001000" => data_out <= rom_array(11592);
		when "0010110101001001" => data_out <= rom_array(11593);
		when "0010110101001010" => data_out <= rom_array(11594);
		when "0010110101001011" => data_out <= rom_array(11595);
		when "0010110101001100" => data_out <= rom_array(11596);
		when "0010110101001101" => data_out <= rom_array(11597);
		when "0010110101001110" => data_out <= rom_array(11598);
		when "0010110101001111" => data_out <= rom_array(11599);
		when "0010110101010000" => data_out <= rom_array(11600);
		when "0010110101010001" => data_out <= rom_array(11601);
		when "0010110101010010" => data_out <= rom_array(11602);
		when "0010110101010011" => data_out <= rom_array(11603);
		when "0010110101010100" => data_out <= rom_array(11604);
		when "0010110101010101" => data_out <= rom_array(11605);
		when "0010110101010110" => data_out <= rom_array(11606);
		when "0010110101010111" => data_out <= rom_array(11607);
		when "0010110101011000" => data_out <= rom_array(11608);
		when "0010110101011001" => data_out <= rom_array(11609);
		when "0010110101011010" => data_out <= rom_array(11610);
		when "0010110101011011" => data_out <= rom_array(11611);
		when "0010110101011100" => data_out <= rom_array(11612);
		when "0010110101011101" => data_out <= rom_array(11613);
		when "0010110101011110" => data_out <= rom_array(11614);
		when "0010110101011111" => data_out <= rom_array(11615);
		when "0010110101100000" => data_out <= rom_array(11616);
		when "0010110101100001" => data_out <= rom_array(11617);
		when "0010110101100010" => data_out <= rom_array(11618);
		when "0010110101100011" => data_out <= rom_array(11619);
		when "0010110101100100" => data_out <= rom_array(11620);
		when "0010110101100101" => data_out <= rom_array(11621);
		when "0010110101100110" => data_out <= rom_array(11622);
		when "0010110101100111" => data_out <= rom_array(11623);
		when "0010110101101000" => data_out <= rom_array(11624);
		when "0010110101101001" => data_out <= rom_array(11625);
		when "0010110101101010" => data_out <= rom_array(11626);
		when "0010110101101011" => data_out <= rom_array(11627);
		when "0010110101101100" => data_out <= rom_array(11628);
		when "0010110101101101" => data_out <= rom_array(11629);
		when "0010110101101110" => data_out <= rom_array(11630);
		when "0010110101101111" => data_out <= rom_array(11631);
		when "0010110101110000" => data_out <= rom_array(11632);
		when "0010110101110001" => data_out <= rom_array(11633);
		when "0010110101110010" => data_out <= rom_array(11634);
		when "0010110101110011" => data_out <= rom_array(11635);
		when "0010110101110100" => data_out <= rom_array(11636);
		when "0010110101110101" => data_out <= rom_array(11637);
		when "0010110101110110" => data_out <= rom_array(11638);
		when "0010110101110111" => data_out <= rom_array(11639);
		when "0010110101111000" => data_out <= rom_array(11640);
		when "0010110101111001" => data_out <= rom_array(11641);
		when "0010110101111010" => data_out <= rom_array(11642);
		when "0010110101111011" => data_out <= rom_array(11643);
		when "0010110101111100" => data_out <= rom_array(11644);
		when "0010110101111101" => data_out <= rom_array(11645);
		when "0010110101111110" => data_out <= rom_array(11646);
		when "0010110101111111" => data_out <= rom_array(11647);
		when "0010110110000000" => data_out <= rom_array(11648);
		when "0010110110000001" => data_out <= rom_array(11649);
		when "0010110110000010" => data_out <= rom_array(11650);
		when "0010110110000011" => data_out <= rom_array(11651);
		when "0010110110000100" => data_out <= rom_array(11652);
		when "0010110110000101" => data_out <= rom_array(11653);
		when "0010110110000110" => data_out <= rom_array(11654);
		when "0010110110000111" => data_out <= rom_array(11655);
		when "0010110110001000" => data_out <= rom_array(11656);
		when "0010110110001001" => data_out <= rom_array(11657);
		when "0010110110001010" => data_out <= rom_array(11658);
		when "0010110110001011" => data_out <= rom_array(11659);
		when "0010110110001100" => data_out <= rom_array(11660);
		when "0010110110001101" => data_out <= rom_array(11661);
		when "0010110110001110" => data_out <= rom_array(11662);
		when "0010110110001111" => data_out <= rom_array(11663);
		when "0010110110010000" => data_out <= rom_array(11664);
		when "0010110110010001" => data_out <= rom_array(11665);
		when "0010110110010010" => data_out <= rom_array(11666);
		when "0010110110010011" => data_out <= rom_array(11667);
		when "0010110110010100" => data_out <= rom_array(11668);
		when "0010110110010101" => data_out <= rom_array(11669);
		when "0010110110010110" => data_out <= rom_array(11670);
		when "0010110110010111" => data_out <= rom_array(11671);
		when "0010110110011000" => data_out <= rom_array(11672);
		when "0010110110011001" => data_out <= rom_array(11673);
		when "0010110110011010" => data_out <= rom_array(11674);
		when "0010110110011011" => data_out <= rom_array(11675);
		when "0010110110011100" => data_out <= rom_array(11676);
		when "0010110110011101" => data_out <= rom_array(11677);
		when "0010110110011110" => data_out <= rom_array(11678);
		when "0010110110011111" => data_out <= rom_array(11679);
		when "0010110110100000" => data_out <= rom_array(11680);
		when "0010110110100001" => data_out <= rom_array(11681);
		when "0010110110100010" => data_out <= rom_array(11682);
		when "0010110110100011" => data_out <= rom_array(11683);
		when "0010110110100100" => data_out <= rom_array(11684);
		when "0010110110100101" => data_out <= rom_array(11685);
		when "0010110110100110" => data_out <= rom_array(11686);
		when "0010110110100111" => data_out <= rom_array(11687);
		when "0010110110101000" => data_out <= rom_array(11688);
		when "0010110110101001" => data_out <= rom_array(11689);
		when "0010110110101010" => data_out <= rom_array(11690);
		when "0010110110101011" => data_out <= rom_array(11691);
		when "0010110110101100" => data_out <= rom_array(11692);
		when "0010110110101101" => data_out <= rom_array(11693);
		when "0010110110101110" => data_out <= rom_array(11694);
		when "0010110110101111" => data_out <= rom_array(11695);
		when "0010110110110000" => data_out <= rom_array(11696);
		when "0010110110110001" => data_out <= rom_array(11697);
		when "0010110110110010" => data_out <= rom_array(11698);
		when "0010110110110011" => data_out <= rom_array(11699);
		when "0010110110110100" => data_out <= rom_array(11700);
		when "0010110110110101" => data_out <= rom_array(11701);
		when "0010110110110110" => data_out <= rom_array(11702);
		when "0010110110110111" => data_out <= rom_array(11703);
		when "0010110110111000" => data_out <= rom_array(11704);
		when "0010110110111001" => data_out <= rom_array(11705);
		when "0010110110111010" => data_out <= rom_array(11706);
		when "0010110110111011" => data_out <= rom_array(11707);
		when "0010110110111100" => data_out <= rom_array(11708);
		when "0010110110111101" => data_out <= rom_array(11709);
		when "0010110110111110" => data_out <= rom_array(11710);
		when "0010110110111111" => data_out <= rom_array(11711);
		when "0010110111000000" => data_out <= rom_array(11712);
		when "0010110111000001" => data_out <= rom_array(11713);
		when "0010110111000010" => data_out <= rom_array(11714);
		when "0010110111000011" => data_out <= rom_array(11715);
		when "0010110111000100" => data_out <= rom_array(11716);
		when "0010110111000101" => data_out <= rom_array(11717);
		when "0010110111000110" => data_out <= rom_array(11718);
		when "0010110111000111" => data_out <= rom_array(11719);
		when "0010110111001000" => data_out <= rom_array(11720);
		when "0010110111001001" => data_out <= rom_array(11721);
		when "0010110111001010" => data_out <= rom_array(11722);
		when "0010110111001011" => data_out <= rom_array(11723);
		when "0010110111001100" => data_out <= rom_array(11724);
		when "0010110111001101" => data_out <= rom_array(11725);
		when "0010110111001110" => data_out <= rom_array(11726);
		when "0010110111001111" => data_out <= rom_array(11727);
		when "0010110111010000" => data_out <= rom_array(11728);
		when "0010110111010001" => data_out <= rom_array(11729);
		when "0010110111010010" => data_out <= rom_array(11730);
		when "0010110111010011" => data_out <= rom_array(11731);
		when "0010110111010100" => data_out <= rom_array(11732);
		when "0010110111010101" => data_out <= rom_array(11733);
		when "0010110111010110" => data_out <= rom_array(11734);
		when "0010110111010111" => data_out <= rom_array(11735);
		when "0010110111011000" => data_out <= rom_array(11736);
		when "0010110111011001" => data_out <= rom_array(11737);
		when "0010110111011010" => data_out <= rom_array(11738);
		when "0010110111011011" => data_out <= rom_array(11739);
		when "0010110111011100" => data_out <= rom_array(11740);
		when "0010110111011101" => data_out <= rom_array(11741);
		when "0010110111011110" => data_out <= rom_array(11742);
		when "0010110111011111" => data_out <= rom_array(11743);
		when "0010110111100000" => data_out <= rom_array(11744);
		when "0010110111100001" => data_out <= rom_array(11745);
		when "0010110111100010" => data_out <= rom_array(11746);
		when "0010110111100011" => data_out <= rom_array(11747);
		when "0010110111100100" => data_out <= rom_array(11748);
		when "0010110111100101" => data_out <= rom_array(11749);
		when "0010110111100110" => data_out <= rom_array(11750);
		when "0010110111100111" => data_out <= rom_array(11751);
		when "0010110111101000" => data_out <= rom_array(11752);
		when "0010110111101001" => data_out <= rom_array(11753);
		when "0010110111101010" => data_out <= rom_array(11754);
		when "0010110111101011" => data_out <= rom_array(11755);
		when "0010110111101100" => data_out <= rom_array(11756);
		when "0010110111101101" => data_out <= rom_array(11757);
		when "0010110111101110" => data_out <= rom_array(11758);
		when "0010110111101111" => data_out <= rom_array(11759);
		when "0010110111110000" => data_out <= rom_array(11760);
		when "0010110111110001" => data_out <= rom_array(11761);
		when "0010110111110010" => data_out <= rom_array(11762);
		when "0010110111110011" => data_out <= rom_array(11763);
		when "0010110111110100" => data_out <= rom_array(11764);
		when "0010110111110101" => data_out <= rom_array(11765);
		when "0010110111110110" => data_out <= rom_array(11766);
		when "0010110111110111" => data_out <= rom_array(11767);
		when "0010110111111000" => data_out <= rom_array(11768);
		when "0010110111111001" => data_out <= rom_array(11769);
		when "0010110111111010" => data_out <= rom_array(11770);
		when "0010110111111011" => data_out <= rom_array(11771);
		when "0010110111111100" => data_out <= rom_array(11772);
		when "0010110111111101" => data_out <= rom_array(11773);
		when "0010110111111110" => data_out <= rom_array(11774);
		when "0010110111111111" => data_out <= rom_array(11775);
		when "0010111000000000" => data_out <= rom_array(11776);
		when "0010111000000001" => data_out <= rom_array(11777);
		when "0010111000000010" => data_out <= rom_array(11778);
		when "0010111000000011" => data_out <= rom_array(11779);
		when "0010111000000100" => data_out <= rom_array(11780);
		when "0010111000000101" => data_out <= rom_array(11781);
		when "0010111000000110" => data_out <= rom_array(11782);
		when "0010111000000111" => data_out <= rom_array(11783);
		when "0010111000001000" => data_out <= rom_array(11784);
		when "0010111000001001" => data_out <= rom_array(11785);
		when "0010111000001010" => data_out <= rom_array(11786);
		when "0010111000001011" => data_out <= rom_array(11787);
		when "0010111000001100" => data_out <= rom_array(11788);
		when "0010111000001101" => data_out <= rom_array(11789);
		when "0010111000001110" => data_out <= rom_array(11790);
		when "0010111000001111" => data_out <= rom_array(11791);
		when "0010111000010000" => data_out <= rom_array(11792);
		when "0010111000010001" => data_out <= rom_array(11793);
		when "0010111000010010" => data_out <= rom_array(11794);
		when "0010111000010011" => data_out <= rom_array(11795);
		when "0010111000010100" => data_out <= rom_array(11796);
		when "0010111000010101" => data_out <= rom_array(11797);
		when "0010111000010110" => data_out <= rom_array(11798);
		when "0010111000010111" => data_out <= rom_array(11799);
		when "0010111000011000" => data_out <= rom_array(11800);
		when "0010111000011001" => data_out <= rom_array(11801);
		when "0010111000011010" => data_out <= rom_array(11802);
		when "0010111000011011" => data_out <= rom_array(11803);
		when "0010111000011100" => data_out <= rom_array(11804);
		when "0010111000011101" => data_out <= rom_array(11805);
		when "0010111000011110" => data_out <= rom_array(11806);
		when "0010111000011111" => data_out <= rom_array(11807);
		when "0010111000100000" => data_out <= rom_array(11808);
		when "0010111000100001" => data_out <= rom_array(11809);
		when "0010111000100010" => data_out <= rom_array(11810);
		when "0010111000100011" => data_out <= rom_array(11811);
		when "0010111000100100" => data_out <= rom_array(11812);
		when "0010111000100101" => data_out <= rom_array(11813);
		when "0010111000100110" => data_out <= rom_array(11814);
		when "0010111000100111" => data_out <= rom_array(11815);
		when "0010111000101000" => data_out <= rom_array(11816);
		when "0010111000101001" => data_out <= rom_array(11817);
		when "0010111000101010" => data_out <= rom_array(11818);
		when "0010111000101011" => data_out <= rom_array(11819);
		when "0010111000101100" => data_out <= rom_array(11820);
		when "0010111000101101" => data_out <= rom_array(11821);
		when "0010111000101110" => data_out <= rom_array(11822);
		when "0010111000101111" => data_out <= rom_array(11823);
		when "0010111000110000" => data_out <= rom_array(11824);
		when "0010111000110001" => data_out <= rom_array(11825);
		when "0010111000110010" => data_out <= rom_array(11826);
		when "0010111000110011" => data_out <= rom_array(11827);
		when "0010111000110100" => data_out <= rom_array(11828);
		when "0010111000110101" => data_out <= rom_array(11829);
		when "0010111000110110" => data_out <= rom_array(11830);
		when "0010111000110111" => data_out <= rom_array(11831);
		when "0010111000111000" => data_out <= rom_array(11832);
		when "0010111000111001" => data_out <= rom_array(11833);
		when "0010111000111010" => data_out <= rom_array(11834);
		when "0010111000111011" => data_out <= rom_array(11835);
		when "0010111000111100" => data_out <= rom_array(11836);
		when "0010111000111101" => data_out <= rom_array(11837);
		when "0010111000111110" => data_out <= rom_array(11838);
		when "0010111000111111" => data_out <= rom_array(11839);
		when "0010111001000000" => data_out <= rom_array(11840);
		when "0010111001000001" => data_out <= rom_array(11841);
		when "0010111001000010" => data_out <= rom_array(11842);
		when "0010111001000011" => data_out <= rom_array(11843);
		when "0010111001000100" => data_out <= rom_array(11844);
		when "0010111001000101" => data_out <= rom_array(11845);
		when "0010111001000110" => data_out <= rom_array(11846);
		when "0010111001000111" => data_out <= rom_array(11847);
		when "0010111001001000" => data_out <= rom_array(11848);
		when "0010111001001001" => data_out <= rom_array(11849);
		when "0010111001001010" => data_out <= rom_array(11850);
		when "0010111001001011" => data_out <= rom_array(11851);
		when "0010111001001100" => data_out <= rom_array(11852);
		when "0010111001001101" => data_out <= rom_array(11853);
		when "0010111001001110" => data_out <= rom_array(11854);
		when "0010111001001111" => data_out <= rom_array(11855);
		when "0010111001010000" => data_out <= rom_array(11856);
		when "0010111001010001" => data_out <= rom_array(11857);
		when "0010111001010010" => data_out <= rom_array(11858);
		when "0010111001010011" => data_out <= rom_array(11859);
		when "0010111001010100" => data_out <= rom_array(11860);
		when "0010111001010101" => data_out <= rom_array(11861);
		when "0010111001010110" => data_out <= rom_array(11862);
		when "0010111001010111" => data_out <= rom_array(11863);
		when "0010111001011000" => data_out <= rom_array(11864);
		when "0010111001011001" => data_out <= rom_array(11865);
		when "0010111001011010" => data_out <= rom_array(11866);
		when "0010111001011011" => data_out <= rom_array(11867);
		when "0010111001011100" => data_out <= rom_array(11868);
		when "0010111001011101" => data_out <= rom_array(11869);
		when "0010111001011110" => data_out <= rom_array(11870);
		when "0010111001011111" => data_out <= rom_array(11871);
		when "0010111001100000" => data_out <= rom_array(11872);
		when "0010111001100001" => data_out <= rom_array(11873);
		when "0010111001100010" => data_out <= rom_array(11874);
		when "0010111001100011" => data_out <= rom_array(11875);
		when "0010111001100100" => data_out <= rom_array(11876);
		when "0010111001100101" => data_out <= rom_array(11877);
		when "0010111001100110" => data_out <= rom_array(11878);
		when "0010111001100111" => data_out <= rom_array(11879);
		when "0010111001101000" => data_out <= rom_array(11880);
		when "0010111001101001" => data_out <= rom_array(11881);
		when "0010111001101010" => data_out <= rom_array(11882);
		when "0010111001101011" => data_out <= rom_array(11883);
		when "0010111001101100" => data_out <= rom_array(11884);
		when "0010111001101101" => data_out <= rom_array(11885);
		when "0010111001101110" => data_out <= rom_array(11886);
		when "0010111001101111" => data_out <= rom_array(11887);
		when "0010111001110000" => data_out <= rom_array(11888);
		when "0010111001110001" => data_out <= rom_array(11889);
		when "0010111001110010" => data_out <= rom_array(11890);
		when "0010111001110011" => data_out <= rom_array(11891);
		when "0010111001110100" => data_out <= rom_array(11892);
		when "0010111001110101" => data_out <= rom_array(11893);
		when "0010111001110110" => data_out <= rom_array(11894);
		when "0010111001110111" => data_out <= rom_array(11895);
		when "0010111001111000" => data_out <= rom_array(11896);
		when "0010111001111001" => data_out <= rom_array(11897);
		when "0010111001111010" => data_out <= rom_array(11898);
		when "0010111001111011" => data_out <= rom_array(11899);
		when "0010111001111100" => data_out <= rom_array(11900);
		when "0010111001111101" => data_out <= rom_array(11901);
		when "0010111001111110" => data_out <= rom_array(11902);
		when "0010111001111111" => data_out <= rom_array(11903);
		when "0010111010000000" => data_out <= rom_array(11904);
		when "0010111010000001" => data_out <= rom_array(11905);
		when "0010111010000010" => data_out <= rom_array(11906);
		when "0010111010000011" => data_out <= rom_array(11907);
		when "0010111010000100" => data_out <= rom_array(11908);
		when "0010111010000101" => data_out <= rom_array(11909);
		when "0010111010000110" => data_out <= rom_array(11910);
		when "0010111010000111" => data_out <= rom_array(11911);
		when "0010111010001000" => data_out <= rom_array(11912);
		when "0010111010001001" => data_out <= rom_array(11913);
		when "0010111010001010" => data_out <= rom_array(11914);
		when "0010111010001011" => data_out <= rom_array(11915);
		when "0010111010001100" => data_out <= rom_array(11916);
		when "0010111010001101" => data_out <= rom_array(11917);
		when "0010111010001110" => data_out <= rom_array(11918);
		when "0010111010001111" => data_out <= rom_array(11919);
		when "0010111010010000" => data_out <= rom_array(11920);
		when "0010111010010001" => data_out <= rom_array(11921);
		when "0010111010010010" => data_out <= rom_array(11922);
		when "0010111010010011" => data_out <= rom_array(11923);
		when "0010111010010100" => data_out <= rom_array(11924);
		when "0010111010010101" => data_out <= rom_array(11925);
		when "0010111010010110" => data_out <= rom_array(11926);
		when "0010111010010111" => data_out <= rom_array(11927);
		when "0010111010011000" => data_out <= rom_array(11928);
		when "0010111010011001" => data_out <= rom_array(11929);
		when "0010111010011010" => data_out <= rom_array(11930);
		when "0010111010011011" => data_out <= rom_array(11931);
		when "0010111010011100" => data_out <= rom_array(11932);
		when "0010111010011101" => data_out <= rom_array(11933);
		when "0010111010011110" => data_out <= rom_array(11934);
		when "0010111010011111" => data_out <= rom_array(11935);
		when "0010111010100000" => data_out <= rom_array(11936);
		when "0010111010100001" => data_out <= rom_array(11937);
		when "0010111010100010" => data_out <= rom_array(11938);
		when "0010111010100011" => data_out <= rom_array(11939);
		when "0010111010100100" => data_out <= rom_array(11940);
		when "0010111010100101" => data_out <= rom_array(11941);
		when "0010111010100110" => data_out <= rom_array(11942);
		when "0010111010100111" => data_out <= rom_array(11943);
		when "0010111010101000" => data_out <= rom_array(11944);
		when "0010111010101001" => data_out <= rom_array(11945);
		when "0010111010101010" => data_out <= rom_array(11946);
		when "0010111010101011" => data_out <= rom_array(11947);
		when "0010111010101100" => data_out <= rom_array(11948);
		when "0010111010101101" => data_out <= rom_array(11949);
		when "0010111010101110" => data_out <= rom_array(11950);
		when "0010111010101111" => data_out <= rom_array(11951);
		when "0010111010110000" => data_out <= rom_array(11952);
		when "0010111010110001" => data_out <= rom_array(11953);
		when "0010111010110010" => data_out <= rom_array(11954);
		when "0010111010110011" => data_out <= rom_array(11955);
		when "0010111010110100" => data_out <= rom_array(11956);
		when "0010111010110101" => data_out <= rom_array(11957);
		when "0010111010110110" => data_out <= rom_array(11958);
		when "0010111010110111" => data_out <= rom_array(11959);
		when "0010111010111000" => data_out <= rom_array(11960);
		when "0010111010111001" => data_out <= rom_array(11961);
		when "0010111010111010" => data_out <= rom_array(11962);
		when "0010111010111011" => data_out <= rom_array(11963);
		when "0010111010111100" => data_out <= rom_array(11964);
		when "0010111010111101" => data_out <= rom_array(11965);
		when "0010111010111110" => data_out <= rom_array(11966);
		when "0010111010111111" => data_out <= rom_array(11967);
		when "0010111011000000" => data_out <= rom_array(11968);
		when "0010111011000001" => data_out <= rom_array(11969);
		when "0010111011000010" => data_out <= rom_array(11970);
		when "0010111011000011" => data_out <= rom_array(11971);
		when "0010111011000100" => data_out <= rom_array(11972);
		when "0010111011000101" => data_out <= rom_array(11973);
		when "0010111011000110" => data_out <= rom_array(11974);
		when "0010111011000111" => data_out <= rom_array(11975);
		when "0010111011001000" => data_out <= rom_array(11976);
		when "0010111011001001" => data_out <= rom_array(11977);
		when "0010111011001010" => data_out <= rom_array(11978);
		when "0010111011001011" => data_out <= rom_array(11979);
		when "0010111011001100" => data_out <= rom_array(11980);
		when "0010111011001101" => data_out <= rom_array(11981);
		when "0010111011001110" => data_out <= rom_array(11982);
		when "0010111011001111" => data_out <= rom_array(11983);
		when "0010111011010000" => data_out <= rom_array(11984);
		when "0010111011010001" => data_out <= rom_array(11985);
		when "0010111011010010" => data_out <= rom_array(11986);
		when "0010111011010011" => data_out <= rom_array(11987);
		when "0010111011010100" => data_out <= rom_array(11988);
		when "0010111011010101" => data_out <= rom_array(11989);
		when "0010111011010110" => data_out <= rom_array(11990);
		when "0010111011010111" => data_out <= rom_array(11991);
		when "0010111011011000" => data_out <= rom_array(11992);
		when "0010111011011001" => data_out <= rom_array(11993);
		when "0010111011011010" => data_out <= rom_array(11994);
		when "0010111011011011" => data_out <= rom_array(11995);
		when "0010111011011100" => data_out <= rom_array(11996);
		when "0010111011011101" => data_out <= rom_array(11997);
		when "0010111011011110" => data_out <= rom_array(11998);
		when "0010111011011111" => data_out <= rom_array(11999);
		when "0010111011100000" => data_out <= rom_array(12000);
		when "0010111011100001" => data_out <= rom_array(12001);
		when "0010111011100010" => data_out <= rom_array(12002);
		when "0010111011100011" => data_out <= rom_array(12003);
		when "0010111011100100" => data_out <= rom_array(12004);
		when "0010111011100101" => data_out <= rom_array(12005);
		when "0010111011100110" => data_out <= rom_array(12006);
		when "0010111011100111" => data_out <= rom_array(12007);
		when "0010111011101000" => data_out <= rom_array(12008);
		when "0010111011101001" => data_out <= rom_array(12009);
		when "0010111011101010" => data_out <= rom_array(12010);
		when "0010111011101011" => data_out <= rom_array(12011);
		when "0010111011101100" => data_out <= rom_array(12012);
		when "0010111011101101" => data_out <= rom_array(12013);
		when "0010111011101110" => data_out <= rom_array(12014);
		when "0010111011101111" => data_out <= rom_array(12015);
		when "0010111011110000" => data_out <= rom_array(12016);
		when "0010111011110001" => data_out <= rom_array(12017);
		when "0010111011110010" => data_out <= rom_array(12018);
		when "0010111011110011" => data_out <= rom_array(12019);
		when "0010111011110100" => data_out <= rom_array(12020);
		when "0010111011110101" => data_out <= rom_array(12021);
		when "0010111011110110" => data_out <= rom_array(12022);
		when "0010111011110111" => data_out <= rom_array(12023);
		when "0010111011111000" => data_out <= rom_array(12024);
		when "0010111011111001" => data_out <= rom_array(12025);
		when "0010111011111010" => data_out <= rom_array(12026);
		when "0010111011111011" => data_out <= rom_array(12027);
		when "0010111011111100" => data_out <= rom_array(12028);
		when "0010111011111101" => data_out <= rom_array(12029);
		when "0010111011111110" => data_out <= rom_array(12030);
		when "0010111011111111" => data_out <= rom_array(12031);
		when "0010111100000000" => data_out <= rom_array(12032);
		when "0010111100000001" => data_out <= rom_array(12033);
		when "0010111100000010" => data_out <= rom_array(12034);
		when "0010111100000011" => data_out <= rom_array(12035);
		when "0010111100000100" => data_out <= rom_array(12036);
		when "0010111100000101" => data_out <= rom_array(12037);
		when "0010111100000110" => data_out <= rom_array(12038);
		when "0010111100000111" => data_out <= rom_array(12039);
		when "0010111100001000" => data_out <= rom_array(12040);
		when "0010111100001001" => data_out <= rom_array(12041);
		when "0010111100001010" => data_out <= rom_array(12042);
		when "0010111100001011" => data_out <= rom_array(12043);
		when "0010111100001100" => data_out <= rom_array(12044);
		when "0010111100001101" => data_out <= rom_array(12045);
		when "0010111100001110" => data_out <= rom_array(12046);
		when "0010111100001111" => data_out <= rom_array(12047);
		when "0010111100010000" => data_out <= rom_array(12048);
		when "0010111100010001" => data_out <= rom_array(12049);
		when "0010111100010010" => data_out <= rom_array(12050);
		when "0010111100010011" => data_out <= rom_array(12051);
		when "0010111100010100" => data_out <= rom_array(12052);
		when "0010111100010101" => data_out <= rom_array(12053);
		when "0010111100010110" => data_out <= rom_array(12054);
		when "0010111100010111" => data_out <= rom_array(12055);
		when "0010111100011000" => data_out <= rom_array(12056);
		when "0010111100011001" => data_out <= rom_array(12057);
		when "0010111100011010" => data_out <= rom_array(12058);
		when "0010111100011011" => data_out <= rom_array(12059);
		when "0010111100011100" => data_out <= rom_array(12060);
		when "0010111100011101" => data_out <= rom_array(12061);
		when "0010111100011110" => data_out <= rom_array(12062);
		when "0010111100011111" => data_out <= rom_array(12063);
		when "0010111100100000" => data_out <= rom_array(12064);
		when "0010111100100001" => data_out <= rom_array(12065);
		when "0010111100100010" => data_out <= rom_array(12066);
		when "0010111100100011" => data_out <= rom_array(12067);
		when "0010111100100100" => data_out <= rom_array(12068);
		when "0010111100100101" => data_out <= rom_array(12069);
		when "0010111100100110" => data_out <= rom_array(12070);
		when "0010111100100111" => data_out <= rom_array(12071);
		when "0010111100101000" => data_out <= rom_array(12072);
		when "0010111100101001" => data_out <= rom_array(12073);
		when "0010111100101010" => data_out <= rom_array(12074);
		when "0010111100101011" => data_out <= rom_array(12075);
		when "0010111100101100" => data_out <= rom_array(12076);
		when "0010111100101101" => data_out <= rom_array(12077);
		when "0010111100101110" => data_out <= rom_array(12078);
		when "0010111100101111" => data_out <= rom_array(12079);
		when "0010111100110000" => data_out <= rom_array(12080);
		when "0010111100110001" => data_out <= rom_array(12081);
		when "0010111100110010" => data_out <= rom_array(12082);
		when "0010111100110011" => data_out <= rom_array(12083);
		when "0010111100110100" => data_out <= rom_array(12084);
		when "0010111100110101" => data_out <= rom_array(12085);
		when "0010111100110110" => data_out <= rom_array(12086);
		when "0010111100110111" => data_out <= rom_array(12087);
		when "0010111100111000" => data_out <= rom_array(12088);
		when "0010111100111001" => data_out <= rom_array(12089);
		when "0010111100111010" => data_out <= rom_array(12090);
		when "0010111100111011" => data_out <= rom_array(12091);
		when "0010111100111100" => data_out <= rom_array(12092);
		when "0010111100111101" => data_out <= rom_array(12093);
		when "0010111100111110" => data_out <= rom_array(12094);
		when "0010111100111111" => data_out <= rom_array(12095);
		when "0010111101000000" => data_out <= rom_array(12096);
		when "0010111101000001" => data_out <= rom_array(12097);
		when "0010111101000010" => data_out <= rom_array(12098);
		when "0010111101000011" => data_out <= rom_array(12099);
		when "0010111101000100" => data_out <= rom_array(12100);
		when "0010111101000101" => data_out <= rom_array(12101);
		when "0010111101000110" => data_out <= rom_array(12102);
		when "0010111101000111" => data_out <= rom_array(12103);
		when "0010111101001000" => data_out <= rom_array(12104);
		when "0010111101001001" => data_out <= rom_array(12105);
		when "0010111101001010" => data_out <= rom_array(12106);
		when "0010111101001011" => data_out <= rom_array(12107);
		when "0010111101001100" => data_out <= rom_array(12108);
		when "0010111101001101" => data_out <= rom_array(12109);
		when "0010111101001110" => data_out <= rom_array(12110);
		when "0010111101001111" => data_out <= rom_array(12111);
		when "0010111101010000" => data_out <= rom_array(12112);
		when "0010111101010001" => data_out <= rom_array(12113);
		when "0010111101010010" => data_out <= rom_array(12114);
		when "0010111101010011" => data_out <= rom_array(12115);
		when "0010111101010100" => data_out <= rom_array(12116);
		when "0010111101010101" => data_out <= rom_array(12117);
		when "0010111101010110" => data_out <= rom_array(12118);
		when "0010111101010111" => data_out <= rom_array(12119);
		when "0010111101011000" => data_out <= rom_array(12120);
		when "0010111101011001" => data_out <= rom_array(12121);
		when "0010111101011010" => data_out <= rom_array(12122);
		when "0010111101011011" => data_out <= rom_array(12123);
		when "0010111101011100" => data_out <= rom_array(12124);
		when "0010111101011101" => data_out <= rom_array(12125);
		when "0010111101011110" => data_out <= rom_array(12126);
		when "0010111101011111" => data_out <= rom_array(12127);
		when "0010111101100000" => data_out <= rom_array(12128);
		when "0010111101100001" => data_out <= rom_array(12129);
		when "0010111101100010" => data_out <= rom_array(12130);
		when "0010111101100011" => data_out <= rom_array(12131);
		when "0010111101100100" => data_out <= rom_array(12132);
		when "0010111101100101" => data_out <= rom_array(12133);
		when "0010111101100110" => data_out <= rom_array(12134);
		when "0010111101100111" => data_out <= rom_array(12135);
		when "0010111101101000" => data_out <= rom_array(12136);
		when "0010111101101001" => data_out <= rom_array(12137);
		when "0010111101101010" => data_out <= rom_array(12138);
		when "0010111101101011" => data_out <= rom_array(12139);
		when "0010111101101100" => data_out <= rom_array(12140);
		when "0010111101101101" => data_out <= rom_array(12141);
		when "0010111101101110" => data_out <= rom_array(12142);
		when "0010111101101111" => data_out <= rom_array(12143);
		when "0010111101110000" => data_out <= rom_array(12144);
		when "0010111101110001" => data_out <= rom_array(12145);
		when "0010111101110010" => data_out <= rom_array(12146);
		when "0010111101110011" => data_out <= rom_array(12147);
		when "0010111101110100" => data_out <= rom_array(12148);
		when "0010111101110101" => data_out <= rom_array(12149);
		when "0010111101110110" => data_out <= rom_array(12150);
		when "0010111101110111" => data_out <= rom_array(12151);
		when "0010111101111000" => data_out <= rom_array(12152);
		when "0010111101111001" => data_out <= rom_array(12153);
		when "0010111101111010" => data_out <= rom_array(12154);
		when "0010111101111011" => data_out <= rom_array(12155);
		when "0010111101111100" => data_out <= rom_array(12156);
		when "0010111101111101" => data_out <= rom_array(12157);
		when "0010111101111110" => data_out <= rom_array(12158);
		when "0010111101111111" => data_out <= rom_array(12159);
		when "0010111110000000" => data_out <= rom_array(12160);
		when "0010111110000001" => data_out <= rom_array(12161);
		when "0010111110000010" => data_out <= rom_array(12162);
		when "0010111110000011" => data_out <= rom_array(12163);
		when "0010111110000100" => data_out <= rom_array(12164);
		when "0010111110000101" => data_out <= rom_array(12165);
		when "0010111110000110" => data_out <= rom_array(12166);
		when "0010111110000111" => data_out <= rom_array(12167);
		when "0010111110001000" => data_out <= rom_array(12168);
		when "0010111110001001" => data_out <= rom_array(12169);
		when "0010111110001010" => data_out <= rom_array(12170);
		when "0010111110001011" => data_out <= rom_array(12171);
		when "0010111110001100" => data_out <= rom_array(12172);
		when "0010111110001101" => data_out <= rom_array(12173);
		when "0010111110001110" => data_out <= rom_array(12174);
		when "0010111110001111" => data_out <= rom_array(12175);
		when "0010111110010000" => data_out <= rom_array(12176);
		when "0010111110010001" => data_out <= rom_array(12177);
		when "0010111110010010" => data_out <= rom_array(12178);
		when "0010111110010011" => data_out <= rom_array(12179);
		when "0010111110010100" => data_out <= rom_array(12180);
		when "0010111110010101" => data_out <= rom_array(12181);
		when "0010111110010110" => data_out <= rom_array(12182);
		when "0010111110010111" => data_out <= rom_array(12183);
		when "0010111110011000" => data_out <= rom_array(12184);
		when "0010111110011001" => data_out <= rom_array(12185);
		when "0010111110011010" => data_out <= rom_array(12186);
		when "0010111110011011" => data_out <= rom_array(12187);
		when "0010111110011100" => data_out <= rom_array(12188);
		when "0010111110011101" => data_out <= rom_array(12189);
		when "0010111110011110" => data_out <= rom_array(12190);
		when "0010111110011111" => data_out <= rom_array(12191);
		when "0010111110100000" => data_out <= rom_array(12192);
		when "0010111110100001" => data_out <= rom_array(12193);
		when "0010111110100010" => data_out <= rom_array(12194);
		when "0010111110100011" => data_out <= rom_array(12195);
		when "0010111110100100" => data_out <= rom_array(12196);
		when "0010111110100101" => data_out <= rom_array(12197);
		when "0010111110100110" => data_out <= rom_array(12198);
		when "0010111110100111" => data_out <= rom_array(12199);
		when "0010111110101000" => data_out <= rom_array(12200);
		when "0010111110101001" => data_out <= rom_array(12201);
		when "0010111110101010" => data_out <= rom_array(12202);
		when "0010111110101011" => data_out <= rom_array(12203);
		when "0010111110101100" => data_out <= rom_array(12204);
		when "0010111110101101" => data_out <= rom_array(12205);
		when "0010111110101110" => data_out <= rom_array(12206);
		when "0010111110101111" => data_out <= rom_array(12207);
		when "0010111110110000" => data_out <= rom_array(12208);
		when "0010111110110001" => data_out <= rom_array(12209);
		when "0010111110110010" => data_out <= rom_array(12210);
		when "0010111110110011" => data_out <= rom_array(12211);
		when "0010111110110100" => data_out <= rom_array(12212);
		when "0010111110110101" => data_out <= rom_array(12213);
		when "0010111110110110" => data_out <= rom_array(12214);
		when "0010111110110111" => data_out <= rom_array(12215);
		when "0010111110111000" => data_out <= rom_array(12216);
		when "0010111110111001" => data_out <= rom_array(12217);
		when "0010111110111010" => data_out <= rom_array(12218);
		when "0010111110111011" => data_out <= rom_array(12219);
		when "0010111110111100" => data_out <= rom_array(12220);
		when "0010111110111101" => data_out <= rom_array(12221);
		when "0010111110111110" => data_out <= rom_array(12222);
		when "0010111110111111" => data_out <= rom_array(12223);
		when "0010111111000000" => data_out <= rom_array(12224);
		when "0010111111000001" => data_out <= rom_array(12225);
		when "0010111111000010" => data_out <= rom_array(12226);
		when "0010111111000011" => data_out <= rom_array(12227);
		when "0010111111000100" => data_out <= rom_array(12228);
		when "0010111111000101" => data_out <= rom_array(12229);
		when "0010111111000110" => data_out <= rom_array(12230);
		when "0010111111000111" => data_out <= rom_array(12231);
		when "0010111111001000" => data_out <= rom_array(12232);
		when "0010111111001001" => data_out <= rom_array(12233);
		when "0010111111001010" => data_out <= rom_array(12234);
		when "0010111111001011" => data_out <= rom_array(12235);
		when "0010111111001100" => data_out <= rom_array(12236);
		when "0010111111001101" => data_out <= rom_array(12237);
		when "0010111111001110" => data_out <= rom_array(12238);
		when "0010111111001111" => data_out <= rom_array(12239);
		when "0010111111010000" => data_out <= rom_array(12240);
		when "0010111111010001" => data_out <= rom_array(12241);
		when "0010111111010010" => data_out <= rom_array(12242);
		when "0010111111010011" => data_out <= rom_array(12243);
		when "0010111111010100" => data_out <= rom_array(12244);
		when "0010111111010101" => data_out <= rom_array(12245);
		when "0010111111010110" => data_out <= rom_array(12246);
		when "0010111111010111" => data_out <= rom_array(12247);
		when "0010111111011000" => data_out <= rom_array(12248);
		when "0010111111011001" => data_out <= rom_array(12249);
		when "0010111111011010" => data_out <= rom_array(12250);
		when "0010111111011011" => data_out <= rom_array(12251);
		when "0010111111011100" => data_out <= rom_array(12252);
		when "0010111111011101" => data_out <= rom_array(12253);
		when "0010111111011110" => data_out <= rom_array(12254);
		when "0010111111011111" => data_out <= rom_array(12255);
		when "0010111111100000" => data_out <= rom_array(12256);
		when "0010111111100001" => data_out <= rom_array(12257);
		when "0010111111100010" => data_out <= rom_array(12258);
		when "0010111111100011" => data_out <= rom_array(12259);
		when "0010111111100100" => data_out <= rom_array(12260);
		when "0010111111100101" => data_out <= rom_array(12261);
		when "0010111111100110" => data_out <= rom_array(12262);
		when "0010111111100111" => data_out <= rom_array(12263);
		when "0010111111101000" => data_out <= rom_array(12264);
		when "0010111111101001" => data_out <= rom_array(12265);
		when "0010111111101010" => data_out <= rom_array(12266);
		when "0010111111101011" => data_out <= rom_array(12267);
		when "0010111111101100" => data_out <= rom_array(12268);
		when "0010111111101101" => data_out <= rom_array(12269);
		when "0010111111101110" => data_out <= rom_array(12270);
		when "0010111111101111" => data_out <= rom_array(12271);
		when "0010111111110000" => data_out <= rom_array(12272);
		when "0010111111110001" => data_out <= rom_array(12273);
		when "0010111111110010" => data_out <= rom_array(12274);
		when "0010111111110011" => data_out <= rom_array(12275);
		when "0010111111110100" => data_out <= rom_array(12276);
		when "0010111111110101" => data_out <= rom_array(12277);
		when "0010111111110110" => data_out <= rom_array(12278);
		when "0010111111110111" => data_out <= rom_array(12279);
		when "0010111111111000" => data_out <= rom_array(12280);
		when "0010111111111001" => data_out <= rom_array(12281);
		when "0010111111111010" => data_out <= rom_array(12282);
		when "0010111111111011" => data_out <= rom_array(12283);
		when "0010111111111100" => data_out <= rom_array(12284);
		when "0010111111111101" => data_out <= rom_array(12285);
		when "0010111111111110" => data_out <= rom_array(12286);
		when "0010111111111111" => data_out <= rom_array(12287);
		when "0011000000000000" => data_out <= rom_array(12288);
		when "0011000000000001" => data_out <= rom_array(12289);
		when "0011000000000010" => data_out <= rom_array(12290);
		when "0011000000000011" => data_out <= rom_array(12291);
		when "0011000000000100" => data_out <= rom_array(12292);
		when "0011000000000101" => data_out <= rom_array(12293);
		when "0011000000000110" => data_out <= rom_array(12294);
		when "0011000000000111" => data_out <= rom_array(12295);
		when "0011000000001000" => data_out <= rom_array(12296);
		when "0011000000001001" => data_out <= rom_array(12297);
		when "0011000000001010" => data_out <= rom_array(12298);
		when "0011000000001011" => data_out <= rom_array(12299);
		when "0011000000001100" => data_out <= rom_array(12300);
		when "0011000000001101" => data_out <= rom_array(12301);
		when "0011000000001110" => data_out <= rom_array(12302);
		when "0011000000001111" => data_out <= rom_array(12303);
		when "0011000000010000" => data_out <= rom_array(12304);
		when "0011000000010001" => data_out <= rom_array(12305);
		when "0011000000010010" => data_out <= rom_array(12306);
		when "0011000000010011" => data_out <= rom_array(12307);
		when "0011000000010100" => data_out <= rom_array(12308);
		when "0011000000010101" => data_out <= rom_array(12309);
		when "0011000000010110" => data_out <= rom_array(12310);
		when "0011000000010111" => data_out <= rom_array(12311);
		when "0011000000011000" => data_out <= rom_array(12312);
		when "0011000000011001" => data_out <= rom_array(12313);
		when "0011000000011010" => data_out <= rom_array(12314);
		when "0011000000011011" => data_out <= rom_array(12315);
		when "0011000000011100" => data_out <= rom_array(12316);
		when "0011000000011101" => data_out <= rom_array(12317);
		when "0011000000011110" => data_out <= rom_array(12318);
		when "0011000000011111" => data_out <= rom_array(12319);
		when "0011000000100000" => data_out <= rom_array(12320);
		when "0011000000100001" => data_out <= rom_array(12321);
		when "0011000000100010" => data_out <= rom_array(12322);
		when "0011000000100011" => data_out <= rom_array(12323);
		when "0011000000100100" => data_out <= rom_array(12324);
		when "0011000000100101" => data_out <= rom_array(12325);
		when "0011000000100110" => data_out <= rom_array(12326);
		when "0011000000100111" => data_out <= rom_array(12327);
		when "0011000000101000" => data_out <= rom_array(12328);
		when "0011000000101001" => data_out <= rom_array(12329);
		when "0011000000101010" => data_out <= rom_array(12330);
		when "0011000000101011" => data_out <= rom_array(12331);
		when "0011000000101100" => data_out <= rom_array(12332);
		when "0011000000101101" => data_out <= rom_array(12333);
		when "0011000000101110" => data_out <= rom_array(12334);
		when "0011000000101111" => data_out <= rom_array(12335);
		when "0011000000110000" => data_out <= rom_array(12336);
		when "0011000000110001" => data_out <= rom_array(12337);
		when "0011000000110010" => data_out <= rom_array(12338);
		when "0011000000110011" => data_out <= rom_array(12339);
		when "0011000000110100" => data_out <= rom_array(12340);
		when "0011000000110101" => data_out <= rom_array(12341);
		when "0011000000110110" => data_out <= rom_array(12342);
		when "0011000000110111" => data_out <= rom_array(12343);
		when "0011000000111000" => data_out <= rom_array(12344);
		when "0011000000111001" => data_out <= rom_array(12345);
		when "0011000000111010" => data_out <= rom_array(12346);
		when "0011000000111011" => data_out <= rom_array(12347);
		when "0011000000111100" => data_out <= rom_array(12348);
		when "0011000000111101" => data_out <= rom_array(12349);
		when "0011000000111110" => data_out <= rom_array(12350);
		when "0011000000111111" => data_out <= rom_array(12351);
		when "0011000001000000" => data_out <= rom_array(12352);
		when "0011000001000001" => data_out <= rom_array(12353);
		when "0011000001000010" => data_out <= rom_array(12354);
		when "0011000001000011" => data_out <= rom_array(12355);
		when "0011000001000100" => data_out <= rom_array(12356);
		when "0011000001000101" => data_out <= rom_array(12357);
		when "0011000001000110" => data_out <= rom_array(12358);
		when "0011000001000111" => data_out <= rom_array(12359);
		when "0011000001001000" => data_out <= rom_array(12360);
		when "0011000001001001" => data_out <= rom_array(12361);
		when "0011000001001010" => data_out <= rom_array(12362);
		when "0011000001001011" => data_out <= rom_array(12363);
		when "0011000001001100" => data_out <= rom_array(12364);
		when "0011000001001101" => data_out <= rom_array(12365);
		when "0011000001001110" => data_out <= rom_array(12366);
		when "0011000001001111" => data_out <= rom_array(12367);
		when "0011000001010000" => data_out <= rom_array(12368);
		when "0011000001010001" => data_out <= rom_array(12369);
		when "0011000001010010" => data_out <= rom_array(12370);
		when "0011000001010011" => data_out <= rom_array(12371);
		when "0011000001010100" => data_out <= rom_array(12372);
		when "0011000001010101" => data_out <= rom_array(12373);
		when "0011000001010110" => data_out <= rom_array(12374);
		when "0011000001010111" => data_out <= rom_array(12375);
		when "0011000001011000" => data_out <= rom_array(12376);
		when "0011000001011001" => data_out <= rom_array(12377);
		when "0011000001011010" => data_out <= rom_array(12378);
		when "0011000001011011" => data_out <= rom_array(12379);
		when "0011000001011100" => data_out <= rom_array(12380);
		when "0011000001011101" => data_out <= rom_array(12381);
		when "0011000001011110" => data_out <= rom_array(12382);
		when "0011000001011111" => data_out <= rom_array(12383);
		when "0011000001100000" => data_out <= rom_array(12384);
		when "0011000001100001" => data_out <= rom_array(12385);
		when "0011000001100010" => data_out <= rom_array(12386);
		when "0011000001100011" => data_out <= rom_array(12387);
		when "0011000001100100" => data_out <= rom_array(12388);
		when "0011000001100101" => data_out <= rom_array(12389);
		when "0011000001100110" => data_out <= rom_array(12390);
		when "0011000001100111" => data_out <= rom_array(12391);
		when "0011000001101000" => data_out <= rom_array(12392);
		when "0011000001101001" => data_out <= rom_array(12393);
		when "0011000001101010" => data_out <= rom_array(12394);
		when "0011000001101011" => data_out <= rom_array(12395);
		when "0011000001101100" => data_out <= rom_array(12396);
		when "0011000001101101" => data_out <= rom_array(12397);
		when "0011000001101110" => data_out <= rom_array(12398);
		when "0011000001101111" => data_out <= rom_array(12399);
		when "0011000001110000" => data_out <= rom_array(12400);
		when "0011000001110001" => data_out <= rom_array(12401);
		when "0011000001110010" => data_out <= rom_array(12402);
		when "0011000001110011" => data_out <= rom_array(12403);
		when "0011000001110100" => data_out <= rom_array(12404);
		when "0011000001110101" => data_out <= rom_array(12405);
		when "0011000001110110" => data_out <= rom_array(12406);
		when "0011000001110111" => data_out <= rom_array(12407);
		when "0011000001111000" => data_out <= rom_array(12408);
		when "0011000001111001" => data_out <= rom_array(12409);
		when "0011000001111010" => data_out <= rom_array(12410);
		when "0011000001111011" => data_out <= rom_array(12411);
		when "0011000001111100" => data_out <= rom_array(12412);
		when "0011000001111101" => data_out <= rom_array(12413);
		when "0011000001111110" => data_out <= rom_array(12414);
		when "0011000001111111" => data_out <= rom_array(12415);
		when "0011000010000000" => data_out <= rom_array(12416);
		when "0011000010000001" => data_out <= rom_array(12417);
		when "0011000010000010" => data_out <= rom_array(12418);
		when "0011000010000011" => data_out <= rom_array(12419);
		when "0011000010000100" => data_out <= rom_array(12420);
		when "0011000010000101" => data_out <= rom_array(12421);
		when "0011000010000110" => data_out <= rom_array(12422);
		when "0011000010000111" => data_out <= rom_array(12423);
		when "0011000010001000" => data_out <= rom_array(12424);
		when "0011000010001001" => data_out <= rom_array(12425);
		when "0011000010001010" => data_out <= rom_array(12426);
		when "0011000010001011" => data_out <= rom_array(12427);
		when "0011000010001100" => data_out <= rom_array(12428);
		when "0011000010001101" => data_out <= rom_array(12429);
		when "0011000010001110" => data_out <= rom_array(12430);
		when "0011000010001111" => data_out <= rom_array(12431);
		when "0011000010010000" => data_out <= rom_array(12432);
		when "0011000010010001" => data_out <= rom_array(12433);
		when "0011000010010010" => data_out <= rom_array(12434);
		when "0011000010010011" => data_out <= rom_array(12435);
		when "0011000010010100" => data_out <= rom_array(12436);
		when "0011000010010101" => data_out <= rom_array(12437);
		when "0011000010010110" => data_out <= rom_array(12438);
		when "0011000010010111" => data_out <= rom_array(12439);
		when "0011000010011000" => data_out <= rom_array(12440);
		when "0011000010011001" => data_out <= rom_array(12441);
		when "0011000010011010" => data_out <= rom_array(12442);
		when "0011000010011011" => data_out <= rom_array(12443);
		when "0011000010011100" => data_out <= rom_array(12444);
		when "0011000010011101" => data_out <= rom_array(12445);
		when "0011000010011110" => data_out <= rom_array(12446);
		when "0011000010011111" => data_out <= rom_array(12447);
		when "0011000010100000" => data_out <= rom_array(12448);
		when "0011000010100001" => data_out <= rom_array(12449);
		when "0011000010100010" => data_out <= rom_array(12450);
		when "0011000010100011" => data_out <= rom_array(12451);
		when "0011000010100100" => data_out <= rom_array(12452);
		when "0011000010100101" => data_out <= rom_array(12453);
		when "0011000010100110" => data_out <= rom_array(12454);
		when "0011000010100111" => data_out <= rom_array(12455);
		when "0011000010101000" => data_out <= rom_array(12456);
		when "0011000010101001" => data_out <= rom_array(12457);
		when "0011000010101010" => data_out <= rom_array(12458);
		when "0011000010101011" => data_out <= rom_array(12459);
		when "0011000010101100" => data_out <= rom_array(12460);
		when "0011000010101101" => data_out <= rom_array(12461);
		when "0011000010101110" => data_out <= rom_array(12462);
		when "0011000010101111" => data_out <= rom_array(12463);
		when "0011000010110000" => data_out <= rom_array(12464);
		when "0011000010110001" => data_out <= rom_array(12465);
		when "0011000010110010" => data_out <= rom_array(12466);
		when "0011000010110011" => data_out <= rom_array(12467);
		when "0011000010110100" => data_out <= rom_array(12468);
		when "0011000010110101" => data_out <= rom_array(12469);
		when "0011000010110110" => data_out <= rom_array(12470);
		when "0011000010110111" => data_out <= rom_array(12471);
		when "0011000010111000" => data_out <= rom_array(12472);
		when "0011000010111001" => data_out <= rom_array(12473);
		when "0011000010111010" => data_out <= rom_array(12474);
		when "0011000010111011" => data_out <= rom_array(12475);
		when "0011000010111100" => data_out <= rom_array(12476);
		when "0011000010111101" => data_out <= rom_array(12477);
		when "0011000010111110" => data_out <= rom_array(12478);
		when "0011000010111111" => data_out <= rom_array(12479);
		when "0011000011000000" => data_out <= rom_array(12480);
		when "0011000011000001" => data_out <= rom_array(12481);
		when "0011000011000010" => data_out <= rom_array(12482);
		when "0011000011000011" => data_out <= rom_array(12483);
		when "0011000011000100" => data_out <= rom_array(12484);
		when "0011000011000101" => data_out <= rom_array(12485);
		when "0011000011000110" => data_out <= rom_array(12486);
		when "0011000011000111" => data_out <= rom_array(12487);
		when "0011000011001000" => data_out <= rom_array(12488);
		when "0011000011001001" => data_out <= rom_array(12489);
		when "0011000011001010" => data_out <= rom_array(12490);
		when "0011000011001011" => data_out <= rom_array(12491);
		when "0011000011001100" => data_out <= rom_array(12492);
		when "0011000011001101" => data_out <= rom_array(12493);
		when "0011000011001110" => data_out <= rom_array(12494);
		when "0011000011001111" => data_out <= rom_array(12495);
		when "0011000011010000" => data_out <= rom_array(12496);
		when "0011000011010001" => data_out <= rom_array(12497);
		when "0011000011010010" => data_out <= rom_array(12498);
		when "0011000011010011" => data_out <= rom_array(12499);
		when "0011000011010100" => data_out <= rom_array(12500);
		when "0011000011010101" => data_out <= rom_array(12501);
		when "0011000011010110" => data_out <= rom_array(12502);
		when "0011000011010111" => data_out <= rom_array(12503);
		when "0011000011011000" => data_out <= rom_array(12504);
		when "0011000011011001" => data_out <= rom_array(12505);
		when "0011000011011010" => data_out <= rom_array(12506);
		when "0011000011011011" => data_out <= rom_array(12507);
		when "0011000011011100" => data_out <= rom_array(12508);
		when "0011000011011101" => data_out <= rom_array(12509);
		when "0011000011011110" => data_out <= rom_array(12510);
		when "0011000011011111" => data_out <= rom_array(12511);
		when "0011000011100000" => data_out <= rom_array(12512);
		when "0011000011100001" => data_out <= rom_array(12513);
		when "0011000011100010" => data_out <= rom_array(12514);
		when "0011000011100011" => data_out <= rom_array(12515);
		when "0011000011100100" => data_out <= rom_array(12516);
		when "0011000011100101" => data_out <= rom_array(12517);
		when "0011000011100110" => data_out <= rom_array(12518);
		when "0011000011100111" => data_out <= rom_array(12519);
		when "0011000011101000" => data_out <= rom_array(12520);
		when "0011000011101001" => data_out <= rom_array(12521);
		when "0011000011101010" => data_out <= rom_array(12522);
		when "0011000011101011" => data_out <= rom_array(12523);
		when "0011000011101100" => data_out <= rom_array(12524);
		when "0011000011101101" => data_out <= rom_array(12525);
		when "0011000011101110" => data_out <= rom_array(12526);
		when "0011000011101111" => data_out <= rom_array(12527);
		when "0011000011110000" => data_out <= rom_array(12528);
		when "0011000011110001" => data_out <= rom_array(12529);
		when "0011000011110010" => data_out <= rom_array(12530);
		when "0011000011110011" => data_out <= rom_array(12531);
		when "0011000011110100" => data_out <= rom_array(12532);
		when "0011000011110101" => data_out <= rom_array(12533);
		when "0011000011110110" => data_out <= rom_array(12534);
		when "0011000011110111" => data_out <= rom_array(12535);
		when "0011000011111000" => data_out <= rom_array(12536);
		when "0011000011111001" => data_out <= rom_array(12537);
		when "0011000011111010" => data_out <= rom_array(12538);
		when "0011000011111011" => data_out <= rom_array(12539);
		when "0011000011111100" => data_out <= rom_array(12540);
		when "0011000011111101" => data_out <= rom_array(12541);
		when "0011000011111110" => data_out <= rom_array(12542);
		when "0011000011111111" => data_out <= rom_array(12543);
		when "0011000100000000" => data_out <= rom_array(12544);
		when "0011000100000001" => data_out <= rom_array(12545);
		when "0011000100000010" => data_out <= rom_array(12546);
		when "0011000100000011" => data_out <= rom_array(12547);
		when "0011000100000100" => data_out <= rom_array(12548);
		when "0011000100000101" => data_out <= rom_array(12549);
		when "0011000100000110" => data_out <= rom_array(12550);
		when "0011000100000111" => data_out <= rom_array(12551);
		when "0011000100001000" => data_out <= rom_array(12552);
		when "0011000100001001" => data_out <= rom_array(12553);
		when "0011000100001010" => data_out <= rom_array(12554);
		when "0011000100001011" => data_out <= rom_array(12555);
		when "0011000100001100" => data_out <= rom_array(12556);
		when "0011000100001101" => data_out <= rom_array(12557);
		when "0011000100001110" => data_out <= rom_array(12558);
		when "0011000100001111" => data_out <= rom_array(12559);
		when "0011000100010000" => data_out <= rom_array(12560);
		when "0011000100010001" => data_out <= rom_array(12561);
		when "0011000100010010" => data_out <= rom_array(12562);
		when "0011000100010011" => data_out <= rom_array(12563);
		when "0011000100010100" => data_out <= rom_array(12564);
		when "0011000100010101" => data_out <= rom_array(12565);
		when "0011000100010110" => data_out <= rom_array(12566);
		when "0011000100010111" => data_out <= rom_array(12567);
		when "0011000100011000" => data_out <= rom_array(12568);
		when "0011000100011001" => data_out <= rom_array(12569);
		when "0011000100011010" => data_out <= rom_array(12570);
		when "0011000100011011" => data_out <= rom_array(12571);
		when "0011000100011100" => data_out <= rom_array(12572);
		when "0011000100011101" => data_out <= rom_array(12573);
		when "0011000100011110" => data_out <= rom_array(12574);
		when "0011000100011111" => data_out <= rom_array(12575);
		when "0011000100100000" => data_out <= rom_array(12576);
		when "0011000100100001" => data_out <= rom_array(12577);
		when "0011000100100010" => data_out <= rom_array(12578);
		when "0011000100100011" => data_out <= rom_array(12579);
		when "0011000100100100" => data_out <= rom_array(12580);
		when "0011000100100101" => data_out <= rom_array(12581);
		when "0011000100100110" => data_out <= rom_array(12582);
		when "0011000100100111" => data_out <= rom_array(12583);
		when "0011000100101000" => data_out <= rom_array(12584);
		when "0011000100101001" => data_out <= rom_array(12585);
		when "0011000100101010" => data_out <= rom_array(12586);
		when "0011000100101011" => data_out <= rom_array(12587);
		when "0011000100101100" => data_out <= rom_array(12588);
		when "0011000100101101" => data_out <= rom_array(12589);
		when "0011000100101110" => data_out <= rom_array(12590);
		when "0011000100101111" => data_out <= rom_array(12591);
		when "0011000100110000" => data_out <= rom_array(12592);
		when "0011000100110001" => data_out <= rom_array(12593);
		when "0011000100110010" => data_out <= rom_array(12594);
		when "0011000100110011" => data_out <= rom_array(12595);
		when "0011000100110100" => data_out <= rom_array(12596);
		when "0011000100110101" => data_out <= rom_array(12597);
		when "0011000100110110" => data_out <= rom_array(12598);
		when "0011000100110111" => data_out <= rom_array(12599);
		when "0011000100111000" => data_out <= rom_array(12600);
		when "0011000100111001" => data_out <= rom_array(12601);
		when "0011000100111010" => data_out <= rom_array(12602);
		when "0011000100111011" => data_out <= rom_array(12603);
		when "0011000100111100" => data_out <= rom_array(12604);
		when "0011000100111101" => data_out <= rom_array(12605);
		when "0011000100111110" => data_out <= rom_array(12606);
		when "0011000100111111" => data_out <= rom_array(12607);
		when "0011000101000000" => data_out <= rom_array(12608);
		when "0011000101000001" => data_out <= rom_array(12609);
		when "0011000101000010" => data_out <= rom_array(12610);
		when "0011000101000011" => data_out <= rom_array(12611);
		when "0011000101000100" => data_out <= rom_array(12612);
		when "0011000101000101" => data_out <= rom_array(12613);
		when "0011000101000110" => data_out <= rom_array(12614);
		when "0011000101000111" => data_out <= rom_array(12615);
		when "0011000101001000" => data_out <= rom_array(12616);
		when "0011000101001001" => data_out <= rom_array(12617);
		when "0011000101001010" => data_out <= rom_array(12618);
		when "0011000101001011" => data_out <= rom_array(12619);
		when "0011000101001100" => data_out <= rom_array(12620);
		when "0011000101001101" => data_out <= rom_array(12621);
		when "0011000101001110" => data_out <= rom_array(12622);
		when "0011000101001111" => data_out <= rom_array(12623);
		when "0011000101010000" => data_out <= rom_array(12624);
		when "0011000101010001" => data_out <= rom_array(12625);
		when "0011000101010010" => data_out <= rom_array(12626);
		when "0011000101010011" => data_out <= rom_array(12627);
		when "0011000101010100" => data_out <= rom_array(12628);
		when "0011000101010101" => data_out <= rom_array(12629);
		when "0011000101010110" => data_out <= rom_array(12630);
		when "0011000101010111" => data_out <= rom_array(12631);
		when "0011000101011000" => data_out <= rom_array(12632);
		when "0011000101011001" => data_out <= rom_array(12633);
		when "0011000101011010" => data_out <= rom_array(12634);
		when "0011000101011011" => data_out <= rom_array(12635);
		when "0011000101011100" => data_out <= rom_array(12636);
		when "0011000101011101" => data_out <= rom_array(12637);
		when "0011000101011110" => data_out <= rom_array(12638);
		when "0011000101011111" => data_out <= rom_array(12639);
		when "0011000101100000" => data_out <= rom_array(12640);
		when "0011000101100001" => data_out <= rom_array(12641);
		when "0011000101100010" => data_out <= rom_array(12642);
		when "0011000101100011" => data_out <= rom_array(12643);
		when "0011000101100100" => data_out <= rom_array(12644);
		when "0011000101100101" => data_out <= rom_array(12645);
		when "0011000101100110" => data_out <= rom_array(12646);
		when "0011000101100111" => data_out <= rom_array(12647);
		when "0011000101101000" => data_out <= rom_array(12648);
		when "0011000101101001" => data_out <= rom_array(12649);
		when "0011000101101010" => data_out <= rom_array(12650);
		when "0011000101101011" => data_out <= rom_array(12651);
		when "0011000101101100" => data_out <= rom_array(12652);
		when "0011000101101101" => data_out <= rom_array(12653);
		when "0011000101101110" => data_out <= rom_array(12654);
		when "0011000101101111" => data_out <= rom_array(12655);
		when "0011000101110000" => data_out <= rom_array(12656);
		when "0011000101110001" => data_out <= rom_array(12657);
		when "0011000101110010" => data_out <= rom_array(12658);
		when "0011000101110011" => data_out <= rom_array(12659);
		when "0011000101110100" => data_out <= rom_array(12660);
		when "0011000101110101" => data_out <= rom_array(12661);
		when "0011000101110110" => data_out <= rom_array(12662);
		when "0011000101110111" => data_out <= rom_array(12663);
		when "0011000101111000" => data_out <= rom_array(12664);
		when "0011000101111001" => data_out <= rom_array(12665);
		when "0011000101111010" => data_out <= rom_array(12666);
		when "0011000101111011" => data_out <= rom_array(12667);
		when "0011000101111100" => data_out <= rom_array(12668);
		when "0011000101111101" => data_out <= rom_array(12669);
		when "0011000101111110" => data_out <= rom_array(12670);
		when "0011000101111111" => data_out <= rom_array(12671);
		when "0011000110000000" => data_out <= rom_array(12672);
		when "0011000110000001" => data_out <= rom_array(12673);
		when "0011000110000010" => data_out <= rom_array(12674);
		when "0011000110000011" => data_out <= rom_array(12675);
		when "0011000110000100" => data_out <= rom_array(12676);
		when "0011000110000101" => data_out <= rom_array(12677);
		when "0011000110000110" => data_out <= rom_array(12678);
		when "0011000110000111" => data_out <= rom_array(12679);
		when "0011000110001000" => data_out <= rom_array(12680);
		when "0011000110001001" => data_out <= rom_array(12681);
		when "0011000110001010" => data_out <= rom_array(12682);
		when "0011000110001011" => data_out <= rom_array(12683);
		when "0011000110001100" => data_out <= rom_array(12684);
		when "0011000110001101" => data_out <= rom_array(12685);
		when "0011000110001110" => data_out <= rom_array(12686);
		when "0011000110001111" => data_out <= rom_array(12687);
		when "0011000110010000" => data_out <= rom_array(12688);
		when "0011000110010001" => data_out <= rom_array(12689);
		when "0011000110010010" => data_out <= rom_array(12690);
		when "0011000110010011" => data_out <= rom_array(12691);
		when "0011000110010100" => data_out <= rom_array(12692);
		when "0011000110010101" => data_out <= rom_array(12693);
		when "0011000110010110" => data_out <= rom_array(12694);
		when "0011000110010111" => data_out <= rom_array(12695);
		when "0011000110011000" => data_out <= rom_array(12696);
		when "0011000110011001" => data_out <= rom_array(12697);
		when "0011000110011010" => data_out <= rom_array(12698);
		when "0011000110011011" => data_out <= rom_array(12699);
		when "0011000110011100" => data_out <= rom_array(12700);
		when "0011000110011101" => data_out <= rom_array(12701);
		when "0011000110011110" => data_out <= rom_array(12702);
		when "0011000110011111" => data_out <= rom_array(12703);
		when "0011000110100000" => data_out <= rom_array(12704);
		when "0011000110100001" => data_out <= rom_array(12705);
		when "0011000110100010" => data_out <= rom_array(12706);
		when "0011000110100011" => data_out <= rom_array(12707);
		when "0011000110100100" => data_out <= rom_array(12708);
		when "0011000110100101" => data_out <= rom_array(12709);
		when "0011000110100110" => data_out <= rom_array(12710);
		when "0011000110100111" => data_out <= rom_array(12711);
		when "0011000110101000" => data_out <= rom_array(12712);
		when "0011000110101001" => data_out <= rom_array(12713);
		when "0011000110101010" => data_out <= rom_array(12714);
		when "0011000110101011" => data_out <= rom_array(12715);
		when "0011000110101100" => data_out <= rom_array(12716);
		when "0011000110101101" => data_out <= rom_array(12717);
		when "0011000110101110" => data_out <= rom_array(12718);
		when "0011000110101111" => data_out <= rom_array(12719);
		when "0011000110110000" => data_out <= rom_array(12720);
		when "0011000110110001" => data_out <= rom_array(12721);
		when "0011000110110010" => data_out <= rom_array(12722);
		when "0011000110110011" => data_out <= rom_array(12723);
		when "0011000110110100" => data_out <= rom_array(12724);
		when "0011000110110101" => data_out <= rom_array(12725);
		when "0011000110110110" => data_out <= rom_array(12726);
		when "0011000110110111" => data_out <= rom_array(12727);
		when "0011000110111000" => data_out <= rom_array(12728);
		when "0011000110111001" => data_out <= rom_array(12729);
		when "0011000110111010" => data_out <= rom_array(12730);
		when "0011000110111011" => data_out <= rom_array(12731);
		when "0011000110111100" => data_out <= rom_array(12732);
		when "0011000110111101" => data_out <= rom_array(12733);
		when "0011000110111110" => data_out <= rom_array(12734);
		when "0011000110111111" => data_out <= rom_array(12735);
		when "0011000111000000" => data_out <= rom_array(12736);
		when "0011000111000001" => data_out <= rom_array(12737);
		when "0011000111000010" => data_out <= rom_array(12738);
		when "0011000111000011" => data_out <= rom_array(12739);
		when "0011000111000100" => data_out <= rom_array(12740);
		when "0011000111000101" => data_out <= rom_array(12741);
		when "0011000111000110" => data_out <= rom_array(12742);
		when "0011000111000111" => data_out <= rom_array(12743);
		when "0011000111001000" => data_out <= rom_array(12744);
		when "0011000111001001" => data_out <= rom_array(12745);
		when "0011000111001010" => data_out <= rom_array(12746);
		when "0011000111001011" => data_out <= rom_array(12747);
		when "0011000111001100" => data_out <= rom_array(12748);
		when "0011000111001101" => data_out <= rom_array(12749);
		when "0011000111001110" => data_out <= rom_array(12750);
		when "0011000111001111" => data_out <= rom_array(12751);
		when "0011000111010000" => data_out <= rom_array(12752);
		when "0011000111010001" => data_out <= rom_array(12753);
		when "0011000111010010" => data_out <= rom_array(12754);
		when "0011000111010011" => data_out <= rom_array(12755);
		when "0011000111010100" => data_out <= rom_array(12756);
		when "0011000111010101" => data_out <= rom_array(12757);
		when "0011000111010110" => data_out <= rom_array(12758);
		when "0011000111010111" => data_out <= rom_array(12759);
		when "0011000111011000" => data_out <= rom_array(12760);
		when "0011000111011001" => data_out <= rom_array(12761);
		when "0011000111011010" => data_out <= rom_array(12762);
		when "0011000111011011" => data_out <= rom_array(12763);
		when "0011000111011100" => data_out <= rom_array(12764);
		when "0011000111011101" => data_out <= rom_array(12765);
		when "0011000111011110" => data_out <= rom_array(12766);
		when "0011000111011111" => data_out <= rom_array(12767);
		when "0011000111100000" => data_out <= rom_array(12768);
		when "0011000111100001" => data_out <= rom_array(12769);
		when "0011000111100010" => data_out <= rom_array(12770);
		when "0011000111100011" => data_out <= rom_array(12771);
		when "0011000111100100" => data_out <= rom_array(12772);
		when "0011000111100101" => data_out <= rom_array(12773);
		when "0011000111100110" => data_out <= rom_array(12774);
		when "0011000111100111" => data_out <= rom_array(12775);
		when "0011000111101000" => data_out <= rom_array(12776);
		when "0011000111101001" => data_out <= rom_array(12777);
		when "0011000111101010" => data_out <= rom_array(12778);
		when "0011000111101011" => data_out <= rom_array(12779);
		when "0011000111101100" => data_out <= rom_array(12780);
		when "0011000111101101" => data_out <= rom_array(12781);
		when "0011000111101110" => data_out <= rom_array(12782);
		when "0011000111101111" => data_out <= rom_array(12783);
		when "0011000111110000" => data_out <= rom_array(12784);
		when "0011000111110001" => data_out <= rom_array(12785);
		when "0011000111110010" => data_out <= rom_array(12786);
		when "0011000111110011" => data_out <= rom_array(12787);
		when "0011000111110100" => data_out <= rom_array(12788);
		when "0011000111110101" => data_out <= rom_array(12789);
		when "0011000111110110" => data_out <= rom_array(12790);
		when "0011000111110111" => data_out <= rom_array(12791);
		when "0011000111111000" => data_out <= rom_array(12792);
		when "0011000111111001" => data_out <= rom_array(12793);
		when "0011000111111010" => data_out <= rom_array(12794);
		when "0011000111111011" => data_out <= rom_array(12795);
		when "0011000111111100" => data_out <= rom_array(12796);
		when "0011000111111101" => data_out <= rom_array(12797);
		when "0011000111111110" => data_out <= rom_array(12798);
		when "0011000111111111" => data_out <= rom_array(12799);
		when "0011001000000000" => data_out <= rom_array(12800);
		when "0011001000000001" => data_out <= rom_array(12801);
		when "0011001000000010" => data_out <= rom_array(12802);
		when "0011001000000011" => data_out <= rom_array(12803);
		when "0011001000000100" => data_out <= rom_array(12804);
		when "0011001000000101" => data_out <= rom_array(12805);
		when "0011001000000110" => data_out <= rom_array(12806);
		when "0011001000000111" => data_out <= rom_array(12807);
		when "0011001000001000" => data_out <= rom_array(12808);
		when "0011001000001001" => data_out <= rom_array(12809);
		when "0011001000001010" => data_out <= rom_array(12810);
		when "0011001000001011" => data_out <= rom_array(12811);
		when "0011001000001100" => data_out <= rom_array(12812);
		when "0011001000001101" => data_out <= rom_array(12813);
		when "0011001000001110" => data_out <= rom_array(12814);
		when "0011001000001111" => data_out <= rom_array(12815);
		when "0011001000010000" => data_out <= rom_array(12816);
		when "0011001000010001" => data_out <= rom_array(12817);
		when "0011001000010010" => data_out <= rom_array(12818);
		when "0011001000010011" => data_out <= rom_array(12819);
		when "0011001000010100" => data_out <= rom_array(12820);
		when "0011001000010101" => data_out <= rom_array(12821);
		when "0011001000010110" => data_out <= rom_array(12822);
		when "0011001000010111" => data_out <= rom_array(12823);
		when "0011001000011000" => data_out <= rom_array(12824);
		when "0011001000011001" => data_out <= rom_array(12825);
		when "0011001000011010" => data_out <= rom_array(12826);
		when "0011001000011011" => data_out <= rom_array(12827);
		when "0011001000011100" => data_out <= rom_array(12828);
		when "0011001000011101" => data_out <= rom_array(12829);
		when "0011001000011110" => data_out <= rom_array(12830);
		when "0011001000011111" => data_out <= rom_array(12831);
		when "0011001000100000" => data_out <= rom_array(12832);
		when "0011001000100001" => data_out <= rom_array(12833);
		when "0011001000100010" => data_out <= rom_array(12834);
		when "0011001000100011" => data_out <= rom_array(12835);
		when "0011001000100100" => data_out <= rom_array(12836);
		when "0011001000100101" => data_out <= rom_array(12837);
		when "0011001000100110" => data_out <= rom_array(12838);
		when "0011001000100111" => data_out <= rom_array(12839);
		when "0011001000101000" => data_out <= rom_array(12840);
		when "0011001000101001" => data_out <= rom_array(12841);
		when "0011001000101010" => data_out <= rom_array(12842);
		when "0011001000101011" => data_out <= rom_array(12843);
		when "0011001000101100" => data_out <= rom_array(12844);
		when "0011001000101101" => data_out <= rom_array(12845);
		when "0011001000101110" => data_out <= rom_array(12846);
		when "0011001000101111" => data_out <= rom_array(12847);
		when "0011001000110000" => data_out <= rom_array(12848);
		when "0011001000110001" => data_out <= rom_array(12849);
		when "0011001000110010" => data_out <= rom_array(12850);
		when "0011001000110011" => data_out <= rom_array(12851);
		when "0011001000110100" => data_out <= rom_array(12852);
		when "0011001000110101" => data_out <= rom_array(12853);
		when "0011001000110110" => data_out <= rom_array(12854);
		when "0011001000110111" => data_out <= rom_array(12855);
		when "0011001000111000" => data_out <= rom_array(12856);
		when "0011001000111001" => data_out <= rom_array(12857);
		when "0011001000111010" => data_out <= rom_array(12858);
		when "0011001000111011" => data_out <= rom_array(12859);
		when "0011001000111100" => data_out <= rom_array(12860);
		when "0011001000111101" => data_out <= rom_array(12861);
		when "0011001000111110" => data_out <= rom_array(12862);
		when "0011001000111111" => data_out <= rom_array(12863);
		when "0011001001000000" => data_out <= rom_array(12864);
		when "0011001001000001" => data_out <= rom_array(12865);
		when "0011001001000010" => data_out <= rom_array(12866);
		when "0011001001000011" => data_out <= rom_array(12867);
		when "0011001001000100" => data_out <= rom_array(12868);
		when "0011001001000101" => data_out <= rom_array(12869);
		when "0011001001000110" => data_out <= rom_array(12870);
		when "0011001001000111" => data_out <= rom_array(12871);
		when "0011001001001000" => data_out <= rom_array(12872);
		when "0011001001001001" => data_out <= rom_array(12873);
		when "0011001001001010" => data_out <= rom_array(12874);
		when "0011001001001011" => data_out <= rom_array(12875);
		when "0011001001001100" => data_out <= rom_array(12876);
		when "0011001001001101" => data_out <= rom_array(12877);
		when "0011001001001110" => data_out <= rom_array(12878);
		when "0011001001001111" => data_out <= rom_array(12879);
		when "0011001001010000" => data_out <= rom_array(12880);
		when "0011001001010001" => data_out <= rom_array(12881);
		when "0011001001010010" => data_out <= rom_array(12882);
		when "0011001001010011" => data_out <= rom_array(12883);
		when "0011001001010100" => data_out <= rom_array(12884);
		when "0011001001010101" => data_out <= rom_array(12885);
		when "0011001001010110" => data_out <= rom_array(12886);
		when "0011001001010111" => data_out <= rom_array(12887);
		when "0011001001011000" => data_out <= rom_array(12888);
		when "0011001001011001" => data_out <= rom_array(12889);
		when "0011001001011010" => data_out <= rom_array(12890);
		when "0011001001011011" => data_out <= rom_array(12891);
		when "0011001001011100" => data_out <= rom_array(12892);
		when "0011001001011101" => data_out <= rom_array(12893);
		when "0011001001011110" => data_out <= rom_array(12894);
		when "0011001001011111" => data_out <= rom_array(12895);
		when "0011001001100000" => data_out <= rom_array(12896);
		when "0011001001100001" => data_out <= rom_array(12897);
		when "0011001001100010" => data_out <= rom_array(12898);
		when "0011001001100011" => data_out <= rom_array(12899);
		when "0011001001100100" => data_out <= rom_array(12900);
		when "0011001001100101" => data_out <= rom_array(12901);
		when "0011001001100110" => data_out <= rom_array(12902);
		when "0011001001100111" => data_out <= rom_array(12903);
		when "0011001001101000" => data_out <= rom_array(12904);
		when "0011001001101001" => data_out <= rom_array(12905);
		when "0011001001101010" => data_out <= rom_array(12906);
		when "0011001001101011" => data_out <= rom_array(12907);
		when "0011001001101100" => data_out <= rom_array(12908);
		when "0011001001101101" => data_out <= rom_array(12909);
		when "0011001001101110" => data_out <= rom_array(12910);
		when "0011001001101111" => data_out <= rom_array(12911);
		when "0011001001110000" => data_out <= rom_array(12912);
		when "0011001001110001" => data_out <= rom_array(12913);
		when "0011001001110010" => data_out <= rom_array(12914);
		when "0011001001110011" => data_out <= rom_array(12915);
		when "0011001001110100" => data_out <= rom_array(12916);
		when "0011001001110101" => data_out <= rom_array(12917);
		when "0011001001110110" => data_out <= rom_array(12918);
		when "0011001001110111" => data_out <= rom_array(12919);
		when "0011001001111000" => data_out <= rom_array(12920);
		when "0011001001111001" => data_out <= rom_array(12921);
		when "0011001001111010" => data_out <= rom_array(12922);
		when "0011001001111011" => data_out <= rom_array(12923);
		when "0011001001111100" => data_out <= rom_array(12924);
		when "0011001001111101" => data_out <= rom_array(12925);
		when "0011001001111110" => data_out <= rom_array(12926);
		when "0011001001111111" => data_out <= rom_array(12927);
		when "0011001010000000" => data_out <= rom_array(12928);
		when "0011001010000001" => data_out <= rom_array(12929);
		when "0011001010000010" => data_out <= rom_array(12930);
		when "0011001010000011" => data_out <= rom_array(12931);
		when "0011001010000100" => data_out <= rom_array(12932);
		when "0011001010000101" => data_out <= rom_array(12933);
		when "0011001010000110" => data_out <= rom_array(12934);
		when "0011001010000111" => data_out <= rom_array(12935);
		when "0011001010001000" => data_out <= rom_array(12936);
		when "0011001010001001" => data_out <= rom_array(12937);
		when "0011001010001010" => data_out <= rom_array(12938);
		when "0011001010001011" => data_out <= rom_array(12939);
		when "0011001010001100" => data_out <= rom_array(12940);
		when "0011001010001101" => data_out <= rom_array(12941);
		when "0011001010001110" => data_out <= rom_array(12942);
		when "0011001010001111" => data_out <= rom_array(12943);
		when "0011001010010000" => data_out <= rom_array(12944);
		when "0011001010010001" => data_out <= rom_array(12945);
		when "0011001010010010" => data_out <= rom_array(12946);
		when "0011001010010011" => data_out <= rom_array(12947);
		when "0011001010010100" => data_out <= rom_array(12948);
		when "0011001010010101" => data_out <= rom_array(12949);
		when "0011001010010110" => data_out <= rom_array(12950);
		when "0011001010010111" => data_out <= rom_array(12951);
		when "0011001010011000" => data_out <= rom_array(12952);
		when "0011001010011001" => data_out <= rom_array(12953);
		when "0011001010011010" => data_out <= rom_array(12954);
		when "0011001010011011" => data_out <= rom_array(12955);
		when "0011001010011100" => data_out <= rom_array(12956);
		when "0011001010011101" => data_out <= rom_array(12957);
		when "0011001010011110" => data_out <= rom_array(12958);
		when "0011001010011111" => data_out <= rom_array(12959);
		when "0011001010100000" => data_out <= rom_array(12960);
		when "0011001010100001" => data_out <= rom_array(12961);
		when "0011001010100010" => data_out <= rom_array(12962);
		when "0011001010100011" => data_out <= rom_array(12963);
		when "0011001010100100" => data_out <= rom_array(12964);
		when "0011001010100101" => data_out <= rom_array(12965);
		when "0011001010100110" => data_out <= rom_array(12966);
		when "0011001010100111" => data_out <= rom_array(12967);
		when "0011001010101000" => data_out <= rom_array(12968);
		when "0011001010101001" => data_out <= rom_array(12969);
		when "0011001010101010" => data_out <= rom_array(12970);
		when "0011001010101011" => data_out <= rom_array(12971);
		when "0011001010101100" => data_out <= rom_array(12972);
		when "0011001010101101" => data_out <= rom_array(12973);
		when "0011001010101110" => data_out <= rom_array(12974);
		when "0011001010101111" => data_out <= rom_array(12975);
		when "0011001010110000" => data_out <= rom_array(12976);
		when "0011001010110001" => data_out <= rom_array(12977);
		when "0011001010110010" => data_out <= rom_array(12978);
		when "0011001010110011" => data_out <= rom_array(12979);
		when "0011001010110100" => data_out <= rom_array(12980);
		when "0011001010110101" => data_out <= rom_array(12981);
		when "0011001010110110" => data_out <= rom_array(12982);
		when "0011001010110111" => data_out <= rom_array(12983);
		when "0011001010111000" => data_out <= rom_array(12984);
		when "0011001010111001" => data_out <= rom_array(12985);
		when "0011001010111010" => data_out <= rom_array(12986);
		when "0011001010111011" => data_out <= rom_array(12987);
		when "0011001010111100" => data_out <= rom_array(12988);
		when "0011001010111101" => data_out <= rom_array(12989);
		when "0011001010111110" => data_out <= rom_array(12990);
		when "0011001010111111" => data_out <= rom_array(12991);
		when "0011001011000000" => data_out <= rom_array(12992);
		when "0011001011000001" => data_out <= rom_array(12993);
		when "0011001011000010" => data_out <= rom_array(12994);
		when "0011001011000011" => data_out <= rom_array(12995);
		when "0011001011000100" => data_out <= rom_array(12996);
		when "0011001011000101" => data_out <= rom_array(12997);
		when "0011001011000110" => data_out <= rom_array(12998);
		when "0011001011000111" => data_out <= rom_array(12999);
		when "0011001011001000" => data_out <= rom_array(13000);
		when "0011001011001001" => data_out <= rom_array(13001);
		when "0011001011001010" => data_out <= rom_array(13002);
		when "0011001011001011" => data_out <= rom_array(13003);
		when "0011001011001100" => data_out <= rom_array(13004);
		when "0011001011001101" => data_out <= rom_array(13005);
		when "0011001011001110" => data_out <= rom_array(13006);
		when "0011001011001111" => data_out <= rom_array(13007);
		when "0011001011010000" => data_out <= rom_array(13008);
		when "0011001011010001" => data_out <= rom_array(13009);
		when "0011001011010010" => data_out <= rom_array(13010);
		when "0011001011010011" => data_out <= rom_array(13011);
		when "0011001011010100" => data_out <= rom_array(13012);
		when "0011001011010101" => data_out <= rom_array(13013);
		when "0011001011010110" => data_out <= rom_array(13014);
		when "0011001011010111" => data_out <= rom_array(13015);
		when "0011001011011000" => data_out <= rom_array(13016);
		when "0011001011011001" => data_out <= rom_array(13017);
		when "0011001011011010" => data_out <= rom_array(13018);
		when "0011001011011011" => data_out <= rom_array(13019);
		when "0011001011011100" => data_out <= rom_array(13020);
		when "0011001011011101" => data_out <= rom_array(13021);
		when "0011001011011110" => data_out <= rom_array(13022);
		when "0011001011011111" => data_out <= rom_array(13023);
		when "0011001011100000" => data_out <= rom_array(13024);
		when "0011001011100001" => data_out <= rom_array(13025);
		when "0011001011100010" => data_out <= rom_array(13026);
		when "0011001011100011" => data_out <= rom_array(13027);
		when "0011001011100100" => data_out <= rom_array(13028);
		when "0011001011100101" => data_out <= rom_array(13029);
		when "0011001011100110" => data_out <= rom_array(13030);
		when "0011001011100111" => data_out <= rom_array(13031);
		when "0011001011101000" => data_out <= rom_array(13032);
		when "0011001011101001" => data_out <= rom_array(13033);
		when "0011001011101010" => data_out <= rom_array(13034);
		when "0011001011101011" => data_out <= rom_array(13035);
		when "0011001011101100" => data_out <= rom_array(13036);
		when "0011001011101101" => data_out <= rom_array(13037);
		when "0011001011101110" => data_out <= rom_array(13038);
		when "0011001011101111" => data_out <= rom_array(13039);
		when "0011001011110000" => data_out <= rom_array(13040);
		when "0011001011110001" => data_out <= rom_array(13041);
		when "0011001011110010" => data_out <= rom_array(13042);
		when "0011001011110011" => data_out <= rom_array(13043);
		when "0011001011110100" => data_out <= rom_array(13044);
		when "0011001011110101" => data_out <= rom_array(13045);
		when "0011001011110110" => data_out <= rom_array(13046);
		when "0011001011110111" => data_out <= rom_array(13047);
		when "0011001011111000" => data_out <= rom_array(13048);
		when "0011001011111001" => data_out <= rom_array(13049);
		when "0011001011111010" => data_out <= rom_array(13050);
		when "0011001011111011" => data_out <= rom_array(13051);
		when "0011001011111100" => data_out <= rom_array(13052);
		when "0011001011111101" => data_out <= rom_array(13053);
		when "0011001011111110" => data_out <= rom_array(13054);
		when "0011001011111111" => data_out <= rom_array(13055);
		when "0011001100000000" => data_out <= rom_array(13056);
		when "0011001100000001" => data_out <= rom_array(13057);
		when "0011001100000010" => data_out <= rom_array(13058);
		when "0011001100000011" => data_out <= rom_array(13059);
		when "0011001100000100" => data_out <= rom_array(13060);
		when "0011001100000101" => data_out <= rom_array(13061);
		when "0011001100000110" => data_out <= rom_array(13062);
		when "0011001100000111" => data_out <= rom_array(13063);
		when "0011001100001000" => data_out <= rom_array(13064);
		when "0011001100001001" => data_out <= rom_array(13065);
		when "0011001100001010" => data_out <= rom_array(13066);
		when "0011001100001011" => data_out <= rom_array(13067);
		when "0011001100001100" => data_out <= rom_array(13068);
		when "0011001100001101" => data_out <= rom_array(13069);
		when "0011001100001110" => data_out <= rom_array(13070);
		when "0011001100001111" => data_out <= rom_array(13071);
		when "0011001100010000" => data_out <= rom_array(13072);
		when "0011001100010001" => data_out <= rom_array(13073);
		when "0011001100010010" => data_out <= rom_array(13074);
		when "0011001100010011" => data_out <= rom_array(13075);
		when "0011001100010100" => data_out <= rom_array(13076);
		when "0011001100010101" => data_out <= rom_array(13077);
		when "0011001100010110" => data_out <= rom_array(13078);
		when "0011001100010111" => data_out <= rom_array(13079);
		when "0011001100011000" => data_out <= rom_array(13080);
		when "0011001100011001" => data_out <= rom_array(13081);
		when "0011001100011010" => data_out <= rom_array(13082);
		when "0011001100011011" => data_out <= rom_array(13083);
		when "0011001100011100" => data_out <= rom_array(13084);
		when "0011001100011101" => data_out <= rom_array(13085);
		when "0011001100011110" => data_out <= rom_array(13086);
		when "0011001100011111" => data_out <= rom_array(13087);
		when "0011001100100000" => data_out <= rom_array(13088);
		when "0011001100100001" => data_out <= rom_array(13089);
		when "0011001100100010" => data_out <= rom_array(13090);
		when "0011001100100011" => data_out <= rom_array(13091);
		when "0011001100100100" => data_out <= rom_array(13092);
		when "0011001100100101" => data_out <= rom_array(13093);
		when "0011001100100110" => data_out <= rom_array(13094);
		when "0011001100100111" => data_out <= rom_array(13095);
		when "0011001100101000" => data_out <= rom_array(13096);
		when "0011001100101001" => data_out <= rom_array(13097);
		when "0011001100101010" => data_out <= rom_array(13098);
		when "0011001100101011" => data_out <= rom_array(13099);
		when "0011001100101100" => data_out <= rom_array(13100);
		when "0011001100101101" => data_out <= rom_array(13101);
		when "0011001100101110" => data_out <= rom_array(13102);
		when "0011001100101111" => data_out <= rom_array(13103);
		when "0011001100110000" => data_out <= rom_array(13104);
		when "0011001100110001" => data_out <= rom_array(13105);
		when "0011001100110010" => data_out <= rom_array(13106);
		when "0011001100110011" => data_out <= rom_array(13107);
		when "0011001100110100" => data_out <= rom_array(13108);
		when "0011001100110101" => data_out <= rom_array(13109);
		when "0011001100110110" => data_out <= rom_array(13110);
		when "0011001100110111" => data_out <= rom_array(13111);
		when "0011001100111000" => data_out <= rom_array(13112);
		when "0011001100111001" => data_out <= rom_array(13113);
		when "0011001100111010" => data_out <= rom_array(13114);
		when "0011001100111011" => data_out <= rom_array(13115);
		when "0011001100111100" => data_out <= rom_array(13116);
		when "0011001100111101" => data_out <= rom_array(13117);
		when "0011001100111110" => data_out <= rom_array(13118);
		when "0011001100111111" => data_out <= rom_array(13119);
		when "0011001101000000" => data_out <= rom_array(13120);
		when "0011001101000001" => data_out <= rom_array(13121);
		when "0011001101000010" => data_out <= rom_array(13122);
		when "0011001101000011" => data_out <= rom_array(13123);
		when "0011001101000100" => data_out <= rom_array(13124);
		when "0011001101000101" => data_out <= rom_array(13125);
		when "0011001101000110" => data_out <= rom_array(13126);
		when "0011001101000111" => data_out <= rom_array(13127);
		when "0011001101001000" => data_out <= rom_array(13128);
		when "0011001101001001" => data_out <= rom_array(13129);
		when "0011001101001010" => data_out <= rom_array(13130);
		when "0011001101001011" => data_out <= rom_array(13131);
		when "0011001101001100" => data_out <= rom_array(13132);
		when "0011001101001101" => data_out <= rom_array(13133);
		when "0011001101001110" => data_out <= rom_array(13134);
		when "0011001101001111" => data_out <= rom_array(13135);
		when "0011001101010000" => data_out <= rom_array(13136);
		when "0011001101010001" => data_out <= rom_array(13137);
		when "0011001101010010" => data_out <= rom_array(13138);
		when "0011001101010011" => data_out <= rom_array(13139);
		when "0011001101010100" => data_out <= rom_array(13140);
		when "0011001101010101" => data_out <= rom_array(13141);
		when "0011001101010110" => data_out <= rom_array(13142);
		when "0011001101010111" => data_out <= rom_array(13143);
		when "0011001101011000" => data_out <= rom_array(13144);
		when "0011001101011001" => data_out <= rom_array(13145);
		when "0011001101011010" => data_out <= rom_array(13146);
		when "0011001101011011" => data_out <= rom_array(13147);
		when "0011001101011100" => data_out <= rom_array(13148);
		when "0011001101011101" => data_out <= rom_array(13149);
		when "0011001101011110" => data_out <= rom_array(13150);
		when "0011001101011111" => data_out <= rom_array(13151);
		when "0011001101100000" => data_out <= rom_array(13152);
		when "0011001101100001" => data_out <= rom_array(13153);
		when "0011001101100010" => data_out <= rom_array(13154);
		when "0011001101100011" => data_out <= rom_array(13155);
		when "0011001101100100" => data_out <= rom_array(13156);
		when "0011001101100101" => data_out <= rom_array(13157);
		when "0011001101100110" => data_out <= rom_array(13158);
		when "0011001101100111" => data_out <= rom_array(13159);
		when "0011001101101000" => data_out <= rom_array(13160);
		when "0011001101101001" => data_out <= rom_array(13161);
		when "0011001101101010" => data_out <= rom_array(13162);
		when "0011001101101011" => data_out <= rom_array(13163);
		when "0011001101101100" => data_out <= rom_array(13164);
		when "0011001101101101" => data_out <= rom_array(13165);
		when "0011001101101110" => data_out <= rom_array(13166);
		when "0011001101101111" => data_out <= rom_array(13167);
		when "0011001101110000" => data_out <= rom_array(13168);
		when "0011001101110001" => data_out <= rom_array(13169);
		when "0011001101110010" => data_out <= rom_array(13170);
		when "0011001101110011" => data_out <= rom_array(13171);
		when "0011001101110100" => data_out <= rom_array(13172);
		when "0011001101110101" => data_out <= rom_array(13173);
		when "0011001101110110" => data_out <= rom_array(13174);
		when "0011001101110111" => data_out <= rom_array(13175);
		when "0011001101111000" => data_out <= rom_array(13176);
		when "0011001101111001" => data_out <= rom_array(13177);
		when "0011001101111010" => data_out <= rom_array(13178);
		when "0011001101111011" => data_out <= rom_array(13179);
		when "0011001101111100" => data_out <= rom_array(13180);
		when "0011001101111101" => data_out <= rom_array(13181);
		when "0011001101111110" => data_out <= rom_array(13182);
		when "0011001101111111" => data_out <= rom_array(13183);
		when "0011001110000000" => data_out <= rom_array(13184);
		when "0011001110000001" => data_out <= rom_array(13185);
		when "0011001110000010" => data_out <= rom_array(13186);
		when "0011001110000011" => data_out <= rom_array(13187);
		when "0011001110000100" => data_out <= rom_array(13188);
		when "0011001110000101" => data_out <= rom_array(13189);
		when "0011001110000110" => data_out <= rom_array(13190);
		when "0011001110000111" => data_out <= rom_array(13191);
		when "0011001110001000" => data_out <= rom_array(13192);
		when "0011001110001001" => data_out <= rom_array(13193);
		when "0011001110001010" => data_out <= rom_array(13194);
		when "0011001110001011" => data_out <= rom_array(13195);
		when "0011001110001100" => data_out <= rom_array(13196);
		when "0011001110001101" => data_out <= rom_array(13197);
		when "0011001110001110" => data_out <= rom_array(13198);
		when "0011001110001111" => data_out <= rom_array(13199);
		when "0011001110010000" => data_out <= rom_array(13200);
		when "0011001110010001" => data_out <= rom_array(13201);
		when "0011001110010010" => data_out <= rom_array(13202);
		when "0011001110010011" => data_out <= rom_array(13203);
		when "0011001110010100" => data_out <= rom_array(13204);
		when "0011001110010101" => data_out <= rom_array(13205);
		when "0011001110010110" => data_out <= rom_array(13206);
		when "0011001110010111" => data_out <= rom_array(13207);
		when "0011001110011000" => data_out <= rom_array(13208);
		when "0011001110011001" => data_out <= rom_array(13209);
		when "0011001110011010" => data_out <= rom_array(13210);
		when "0011001110011011" => data_out <= rom_array(13211);
		when "0011001110011100" => data_out <= rom_array(13212);
		when "0011001110011101" => data_out <= rom_array(13213);
		when "0011001110011110" => data_out <= rom_array(13214);
		when "0011001110011111" => data_out <= rom_array(13215);
		when "0011001110100000" => data_out <= rom_array(13216);
		when "0011001110100001" => data_out <= rom_array(13217);
		when "0011001110100010" => data_out <= rom_array(13218);
		when "0011001110100011" => data_out <= rom_array(13219);
		when "0011001110100100" => data_out <= rom_array(13220);
		when "0011001110100101" => data_out <= rom_array(13221);
		when "0011001110100110" => data_out <= rom_array(13222);
		when "0011001110100111" => data_out <= rom_array(13223);
		when "0011001110101000" => data_out <= rom_array(13224);
		when "0011001110101001" => data_out <= rom_array(13225);
		when "0011001110101010" => data_out <= rom_array(13226);
		when "0011001110101011" => data_out <= rom_array(13227);
		when "0011001110101100" => data_out <= rom_array(13228);
		when "0011001110101101" => data_out <= rom_array(13229);
		when "0011001110101110" => data_out <= rom_array(13230);
		when "0011001110101111" => data_out <= rom_array(13231);
		when "0011001110110000" => data_out <= rom_array(13232);
		when "0011001110110001" => data_out <= rom_array(13233);
		when "0011001110110010" => data_out <= rom_array(13234);
		when "0011001110110011" => data_out <= rom_array(13235);
		when "0011001110110100" => data_out <= rom_array(13236);
		when "0011001110110101" => data_out <= rom_array(13237);
		when "0011001110110110" => data_out <= rom_array(13238);
		when "0011001110110111" => data_out <= rom_array(13239);
		when "0011001110111000" => data_out <= rom_array(13240);
		when "0011001110111001" => data_out <= rom_array(13241);
		when "0011001110111010" => data_out <= rom_array(13242);
		when "0011001110111011" => data_out <= rom_array(13243);
		when "0011001110111100" => data_out <= rom_array(13244);
		when "0011001110111101" => data_out <= rom_array(13245);
		when "0011001110111110" => data_out <= rom_array(13246);
		when "0011001110111111" => data_out <= rom_array(13247);
		when "0011001111000000" => data_out <= rom_array(13248);
		when "0011001111000001" => data_out <= rom_array(13249);
		when "0011001111000010" => data_out <= rom_array(13250);
		when "0011001111000011" => data_out <= rom_array(13251);
		when "0011001111000100" => data_out <= rom_array(13252);
		when "0011001111000101" => data_out <= rom_array(13253);
		when "0011001111000110" => data_out <= rom_array(13254);
		when "0011001111000111" => data_out <= rom_array(13255);
		when "0011001111001000" => data_out <= rom_array(13256);
		when "0011001111001001" => data_out <= rom_array(13257);
		when "0011001111001010" => data_out <= rom_array(13258);
		when "0011001111001011" => data_out <= rom_array(13259);
		when "0011001111001100" => data_out <= rom_array(13260);
		when "0011001111001101" => data_out <= rom_array(13261);
		when "0011001111001110" => data_out <= rom_array(13262);
		when "0011001111001111" => data_out <= rom_array(13263);
		when "0011001111010000" => data_out <= rom_array(13264);
		when "0011001111010001" => data_out <= rom_array(13265);
		when "0011001111010010" => data_out <= rom_array(13266);
		when "0011001111010011" => data_out <= rom_array(13267);
		when "0011001111010100" => data_out <= rom_array(13268);
		when "0011001111010101" => data_out <= rom_array(13269);
		when "0011001111010110" => data_out <= rom_array(13270);
		when "0011001111010111" => data_out <= rom_array(13271);
		when "0011001111011000" => data_out <= rom_array(13272);
		when "0011001111011001" => data_out <= rom_array(13273);
		when "0011001111011010" => data_out <= rom_array(13274);
		when "0011001111011011" => data_out <= rom_array(13275);
		when "0011001111011100" => data_out <= rom_array(13276);
		when "0011001111011101" => data_out <= rom_array(13277);
		when "0011001111011110" => data_out <= rom_array(13278);
		when "0011001111011111" => data_out <= rom_array(13279);
		when "0011001111100000" => data_out <= rom_array(13280);
		when "0011001111100001" => data_out <= rom_array(13281);
		when "0011001111100010" => data_out <= rom_array(13282);
		when "0011001111100011" => data_out <= rom_array(13283);
		when "0011001111100100" => data_out <= rom_array(13284);
		when "0011001111100101" => data_out <= rom_array(13285);
		when "0011001111100110" => data_out <= rom_array(13286);
		when "0011001111100111" => data_out <= rom_array(13287);
		when "0011001111101000" => data_out <= rom_array(13288);
		when "0011001111101001" => data_out <= rom_array(13289);
		when "0011001111101010" => data_out <= rom_array(13290);
		when "0011001111101011" => data_out <= rom_array(13291);
		when "0011001111101100" => data_out <= rom_array(13292);
		when "0011001111101101" => data_out <= rom_array(13293);
		when "0011001111101110" => data_out <= rom_array(13294);
		when "0011001111101111" => data_out <= rom_array(13295);
		when "0011001111110000" => data_out <= rom_array(13296);
		when "0011001111110001" => data_out <= rom_array(13297);
		when "0011001111110010" => data_out <= rom_array(13298);
		when "0011001111110011" => data_out <= rom_array(13299);
		when "0011001111110100" => data_out <= rom_array(13300);
		when "0011001111110101" => data_out <= rom_array(13301);
		when "0011001111110110" => data_out <= rom_array(13302);
		when "0011001111110111" => data_out <= rom_array(13303);
		when "0011001111111000" => data_out <= rom_array(13304);
		when "0011001111111001" => data_out <= rom_array(13305);
		when "0011001111111010" => data_out <= rom_array(13306);
		when "0011001111111011" => data_out <= rom_array(13307);
		when "0011001111111100" => data_out <= rom_array(13308);
		when "0011001111111101" => data_out <= rom_array(13309);
		when "0011001111111110" => data_out <= rom_array(13310);
		when "0011001111111111" => data_out <= rom_array(13311);
		when "0011010000000000" => data_out <= rom_array(13312);
		when "0011010000000001" => data_out <= rom_array(13313);
		when "0011010000000010" => data_out <= rom_array(13314);
		when "0011010000000011" => data_out <= rom_array(13315);
		when "0011010000000100" => data_out <= rom_array(13316);
		when "0011010000000101" => data_out <= rom_array(13317);
		when "0011010000000110" => data_out <= rom_array(13318);
		when "0011010000000111" => data_out <= rom_array(13319);
		when "0011010000001000" => data_out <= rom_array(13320);
		when "0011010000001001" => data_out <= rom_array(13321);
		when "0011010000001010" => data_out <= rom_array(13322);
		when "0011010000001011" => data_out <= rom_array(13323);
		when "0011010000001100" => data_out <= rom_array(13324);
		when "0011010000001101" => data_out <= rom_array(13325);
		when "0011010000001110" => data_out <= rom_array(13326);
		when "0011010000001111" => data_out <= rom_array(13327);
		when "0011010000010000" => data_out <= rom_array(13328);
		when "0011010000010001" => data_out <= rom_array(13329);
		when "0011010000010010" => data_out <= rom_array(13330);
		when "0011010000010011" => data_out <= rom_array(13331);
		when "0011010000010100" => data_out <= rom_array(13332);
		when "0011010000010101" => data_out <= rom_array(13333);
		when "0011010000010110" => data_out <= rom_array(13334);
		when "0011010000010111" => data_out <= rom_array(13335);
		when "0011010000011000" => data_out <= rom_array(13336);
		when "0011010000011001" => data_out <= rom_array(13337);
		when "0011010000011010" => data_out <= rom_array(13338);
		when "0011010000011011" => data_out <= rom_array(13339);
		when "0011010000011100" => data_out <= rom_array(13340);
		when "0011010000011101" => data_out <= rom_array(13341);
		when "0011010000011110" => data_out <= rom_array(13342);
		when "0011010000011111" => data_out <= rom_array(13343);
		when "0011010000100000" => data_out <= rom_array(13344);
		when "0011010000100001" => data_out <= rom_array(13345);
		when "0011010000100010" => data_out <= rom_array(13346);
		when "0011010000100011" => data_out <= rom_array(13347);
		when "0011010000100100" => data_out <= rom_array(13348);
		when "0011010000100101" => data_out <= rom_array(13349);
		when "0011010000100110" => data_out <= rom_array(13350);
		when "0011010000100111" => data_out <= rom_array(13351);
		when "0011010000101000" => data_out <= rom_array(13352);
		when "0011010000101001" => data_out <= rom_array(13353);
		when "0011010000101010" => data_out <= rom_array(13354);
		when "0011010000101011" => data_out <= rom_array(13355);
		when "0011010000101100" => data_out <= rom_array(13356);
		when "0011010000101101" => data_out <= rom_array(13357);
		when "0011010000101110" => data_out <= rom_array(13358);
		when "0011010000101111" => data_out <= rom_array(13359);
		when "0011010000110000" => data_out <= rom_array(13360);
		when "0011010000110001" => data_out <= rom_array(13361);
		when "0011010000110010" => data_out <= rom_array(13362);
		when "0011010000110011" => data_out <= rom_array(13363);
		when "0011010000110100" => data_out <= rom_array(13364);
		when "0011010000110101" => data_out <= rom_array(13365);
		when "0011010000110110" => data_out <= rom_array(13366);
		when "0011010000110111" => data_out <= rom_array(13367);
		when "0011010000111000" => data_out <= rom_array(13368);
		when "0011010000111001" => data_out <= rom_array(13369);
		when "0011010000111010" => data_out <= rom_array(13370);
		when "0011010000111011" => data_out <= rom_array(13371);
		when "0011010000111100" => data_out <= rom_array(13372);
		when "0011010000111101" => data_out <= rom_array(13373);
		when "0011010000111110" => data_out <= rom_array(13374);
		when "0011010000111111" => data_out <= rom_array(13375);
		when "0011010001000000" => data_out <= rom_array(13376);
		when "0011010001000001" => data_out <= rom_array(13377);
		when "0011010001000010" => data_out <= rom_array(13378);
		when "0011010001000011" => data_out <= rom_array(13379);
		when "0011010001000100" => data_out <= rom_array(13380);
		when "0011010001000101" => data_out <= rom_array(13381);
		when "0011010001000110" => data_out <= rom_array(13382);
		when "0011010001000111" => data_out <= rom_array(13383);
		when "0011010001001000" => data_out <= rom_array(13384);
		when "0011010001001001" => data_out <= rom_array(13385);
		when "0011010001001010" => data_out <= rom_array(13386);
		when "0011010001001011" => data_out <= rom_array(13387);
		when "0011010001001100" => data_out <= rom_array(13388);
		when "0011010001001101" => data_out <= rom_array(13389);
		when "0011010001001110" => data_out <= rom_array(13390);
		when "0011010001001111" => data_out <= rom_array(13391);
		when "0011010001010000" => data_out <= rom_array(13392);
		when "0011010001010001" => data_out <= rom_array(13393);
		when "0011010001010010" => data_out <= rom_array(13394);
		when "0011010001010011" => data_out <= rom_array(13395);
		when "0011010001010100" => data_out <= rom_array(13396);
		when "0011010001010101" => data_out <= rom_array(13397);
		when "0011010001010110" => data_out <= rom_array(13398);
		when "0011010001010111" => data_out <= rom_array(13399);
		when "0011010001011000" => data_out <= rom_array(13400);
		when "0011010001011001" => data_out <= rom_array(13401);
		when "0011010001011010" => data_out <= rom_array(13402);
		when "0011010001011011" => data_out <= rom_array(13403);
		when "0011010001011100" => data_out <= rom_array(13404);
		when "0011010001011101" => data_out <= rom_array(13405);
		when "0011010001011110" => data_out <= rom_array(13406);
		when "0011010001011111" => data_out <= rom_array(13407);
		when "0011010001100000" => data_out <= rom_array(13408);
		when "0011010001100001" => data_out <= rom_array(13409);
		when "0011010001100010" => data_out <= rom_array(13410);
		when "0011010001100011" => data_out <= rom_array(13411);
		when "0011010001100100" => data_out <= rom_array(13412);
		when "0011010001100101" => data_out <= rom_array(13413);
		when "0011010001100110" => data_out <= rom_array(13414);
		when "0011010001100111" => data_out <= rom_array(13415);
		when "0011010001101000" => data_out <= rom_array(13416);
		when "0011010001101001" => data_out <= rom_array(13417);
		when "0011010001101010" => data_out <= rom_array(13418);
		when "0011010001101011" => data_out <= rom_array(13419);
		when "0011010001101100" => data_out <= rom_array(13420);
		when "0011010001101101" => data_out <= rom_array(13421);
		when "0011010001101110" => data_out <= rom_array(13422);
		when "0011010001101111" => data_out <= rom_array(13423);
		when "0011010001110000" => data_out <= rom_array(13424);
		when "0011010001110001" => data_out <= rom_array(13425);
		when "0011010001110010" => data_out <= rom_array(13426);
		when "0011010001110011" => data_out <= rom_array(13427);
		when "0011010001110100" => data_out <= rom_array(13428);
		when "0011010001110101" => data_out <= rom_array(13429);
		when "0011010001110110" => data_out <= rom_array(13430);
		when "0011010001110111" => data_out <= rom_array(13431);
		when "0011010001111000" => data_out <= rom_array(13432);
		when "0011010001111001" => data_out <= rom_array(13433);
		when "0011010001111010" => data_out <= rom_array(13434);
		when "0011010001111011" => data_out <= rom_array(13435);
		when "0011010001111100" => data_out <= rom_array(13436);
		when "0011010001111101" => data_out <= rom_array(13437);
		when "0011010001111110" => data_out <= rom_array(13438);
		when "0011010001111111" => data_out <= rom_array(13439);
		when "0011010010000000" => data_out <= rom_array(13440);
		when "0011010010000001" => data_out <= rom_array(13441);
		when "0011010010000010" => data_out <= rom_array(13442);
		when "0011010010000011" => data_out <= rom_array(13443);
		when "0011010010000100" => data_out <= rom_array(13444);
		when "0011010010000101" => data_out <= rom_array(13445);
		when "0011010010000110" => data_out <= rom_array(13446);
		when "0011010010000111" => data_out <= rom_array(13447);
		when "0011010010001000" => data_out <= rom_array(13448);
		when "0011010010001001" => data_out <= rom_array(13449);
		when "0011010010001010" => data_out <= rom_array(13450);
		when "0011010010001011" => data_out <= rom_array(13451);
		when "0011010010001100" => data_out <= rom_array(13452);
		when "0011010010001101" => data_out <= rom_array(13453);
		when "0011010010001110" => data_out <= rom_array(13454);
		when "0011010010001111" => data_out <= rom_array(13455);
		when "0011010010010000" => data_out <= rom_array(13456);
		when "0011010010010001" => data_out <= rom_array(13457);
		when "0011010010010010" => data_out <= rom_array(13458);
		when "0011010010010011" => data_out <= rom_array(13459);
		when "0011010010010100" => data_out <= rom_array(13460);
		when "0011010010010101" => data_out <= rom_array(13461);
		when "0011010010010110" => data_out <= rom_array(13462);
		when "0011010010010111" => data_out <= rom_array(13463);
		when "0011010010011000" => data_out <= rom_array(13464);
		when "0011010010011001" => data_out <= rom_array(13465);
		when "0011010010011010" => data_out <= rom_array(13466);
		when "0011010010011011" => data_out <= rom_array(13467);
		when "0011010010011100" => data_out <= rom_array(13468);
		when "0011010010011101" => data_out <= rom_array(13469);
		when "0011010010011110" => data_out <= rom_array(13470);
		when "0011010010011111" => data_out <= rom_array(13471);
		when "0011010010100000" => data_out <= rom_array(13472);
		when "0011010010100001" => data_out <= rom_array(13473);
		when "0011010010100010" => data_out <= rom_array(13474);
		when "0011010010100011" => data_out <= rom_array(13475);
		when "0011010010100100" => data_out <= rom_array(13476);
		when "0011010010100101" => data_out <= rom_array(13477);
		when "0011010010100110" => data_out <= rom_array(13478);
		when "0011010010100111" => data_out <= rom_array(13479);
		when "0011010010101000" => data_out <= rom_array(13480);
		when "0011010010101001" => data_out <= rom_array(13481);
		when "0011010010101010" => data_out <= rom_array(13482);
		when "0011010010101011" => data_out <= rom_array(13483);
		when "0011010010101100" => data_out <= rom_array(13484);
		when "0011010010101101" => data_out <= rom_array(13485);
		when "0011010010101110" => data_out <= rom_array(13486);
		when "0011010010101111" => data_out <= rom_array(13487);
		when "0011010010110000" => data_out <= rom_array(13488);
		when "0011010010110001" => data_out <= rom_array(13489);
		when "0011010010110010" => data_out <= rom_array(13490);
		when "0011010010110011" => data_out <= rom_array(13491);
		when "0011010010110100" => data_out <= rom_array(13492);
		when "0011010010110101" => data_out <= rom_array(13493);
		when "0011010010110110" => data_out <= rom_array(13494);
		when "0011010010110111" => data_out <= rom_array(13495);
		when "0011010010111000" => data_out <= rom_array(13496);
		when "0011010010111001" => data_out <= rom_array(13497);
		when "0011010010111010" => data_out <= rom_array(13498);
		when "0011010010111011" => data_out <= rom_array(13499);
		when "0011010010111100" => data_out <= rom_array(13500);
		when "0011010010111101" => data_out <= rom_array(13501);
		when "0011010010111110" => data_out <= rom_array(13502);
		when "0011010010111111" => data_out <= rom_array(13503);
		when "0011010011000000" => data_out <= rom_array(13504);
		when "0011010011000001" => data_out <= rom_array(13505);
		when "0011010011000010" => data_out <= rom_array(13506);
		when "0011010011000011" => data_out <= rom_array(13507);
		when "0011010011000100" => data_out <= rom_array(13508);
		when "0011010011000101" => data_out <= rom_array(13509);
		when "0011010011000110" => data_out <= rom_array(13510);
		when "0011010011000111" => data_out <= rom_array(13511);
		when "0011010011001000" => data_out <= rom_array(13512);
		when "0011010011001001" => data_out <= rom_array(13513);
		when "0011010011001010" => data_out <= rom_array(13514);
		when "0011010011001011" => data_out <= rom_array(13515);
		when "0011010011001100" => data_out <= rom_array(13516);
		when "0011010011001101" => data_out <= rom_array(13517);
		when "0011010011001110" => data_out <= rom_array(13518);
		when "0011010011001111" => data_out <= rom_array(13519);
		when "0011010011010000" => data_out <= rom_array(13520);
		when "0011010011010001" => data_out <= rom_array(13521);
		when "0011010011010010" => data_out <= rom_array(13522);
		when "0011010011010011" => data_out <= rom_array(13523);
		when "0011010011010100" => data_out <= rom_array(13524);
		when "0011010011010101" => data_out <= rom_array(13525);
		when "0011010011010110" => data_out <= rom_array(13526);
		when "0011010011010111" => data_out <= rom_array(13527);
		when "0011010011011000" => data_out <= rom_array(13528);
		when "0011010011011001" => data_out <= rom_array(13529);
		when "0011010011011010" => data_out <= rom_array(13530);
		when "0011010011011011" => data_out <= rom_array(13531);
		when "0011010011011100" => data_out <= rom_array(13532);
		when "0011010011011101" => data_out <= rom_array(13533);
		when "0011010011011110" => data_out <= rom_array(13534);
		when "0011010011011111" => data_out <= rom_array(13535);
		when "0011010011100000" => data_out <= rom_array(13536);
		when "0011010011100001" => data_out <= rom_array(13537);
		when "0011010011100010" => data_out <= rom_array(13538);
		when "0011010011100011" => data_out <= rom_array(13539);
		when "0011010011100100" => data_out <= rom_array(13540);
		when "0011010011100101" => data_out <= rom_array(13541);
		when "0011010011100110" => data_out <= rom_array(13542);
		when "0011010011100111" => data_out <= rom_array(13543);
		when "0011010011101000" => data_out <= rom_array(13544);
		when "0011010011101001" => data_out <= rom_array(13545);
		when "0011010011101010" => data_out <= rom_array(13546);
		when "0011010011101011" => data_out <= rom_array(13547);
		when "0011010011101100" => data_out <= rom_array(13548);
		when "0011010011101101" => data_out <= rom_array(13549);
		when "0011010011101110" => data_out <= rom_array(13550);
		when "0011010011101111" => data_out <= rom_array(13551);
		when "0011010011110000" => data_out <= rom_array(13552);
		when "0011010011110001" => data_out <= rom_array(13553);
		when "0011010011110010" => data_out <= rom_array(13554);
		when "0011010011110011" => data_out <= rom_array(13555);
		when "0011010011110100" => data_out <= rom_array(13556);
		when "0011010011110101" => data_out <= rom_array(13557);
		when "0011010011110110" => data_out <= rom_array(13558);
		when "0011010011110111" => data_out <= rom_array(13559);
		when "0011010011111000" => data_out <= rom_array(13560);
		when "0011010011111001" => data_out <= rom_array(13561);
		when "0011010011111010" => data_out <= rom_array(13562);
		when "0011010011111011" => data_out <= rom_array(13563);
		when "0011010011111100" => data_out <= rom_array(13564);
		when "0011010011111101" => data_out <= rom_array(13565);
		when "0011010011111110" => data_out <= rom_array(13566);
		when "0011010011111111" => data_out <= rom_array(13567);
		when "0011010100000000" => data_out <= rom_array(13568);
		when "0011010100000001" => data_out <= rom_array(13569);
		when "0011010100000010" => data_out <= rom_array(13570);
		when "0011010100000011" => data_out <= rom_array(13571);
		when "0011010100000100" => data_out <= rom_array(13572);
		when "0011010100000101" => data_out <= rom_array(13573);
		when "0011010100000110" => data_out <= rom_array(13574);
		when "0011010100000111" => data_out <= rom_array(13575);
		when "0011010100001000" => data_out <= rom_array(13576);
		when "0011010100001001" => data_out <= rom_array(13577);
		when "0011010100001010" => data_out <= rom_array(13578);
		when "0011010100001011" => data_out <= rom_array(13579);
		when "0011010100001100" => data_out <= rom_array(13580);
		when "0011010100001101" => data_out <= rom_array(13581);
		when "0011010100001110" => data_out <= rom_array(13582);
		when "0011010100001111" => data_out <= rom_array(13583);
		when "0011010100010000" => data_out <= rom_array(13584);
		when "0011010100010001" => data_out <= rom_array(13585);
		when "0011010100010010" => data_out <= rom_array(13586);
		when "0011010100010011" => data_out <= rom_array(13587);
		when "0011010100010100" => data_out <= rom_array(13588);
		when "0011010100010101" => data_out <= rom_array(13589);
		when "0011010100010110" => data_out <= rom_array(13590);
		when "0011010100010111" => data_out <= rom_array(13591);
		when "0011010100011000" => data_out <= rom_array(13592);
		when "0011010100011001" => data_out <= rom_array(13593);
		when "0011010100011010" => data_out <= rom_array(13594);
		when "0011010100011011" => data_out <= rom_array(13595);
		when "0011010100011100" => data_out <= rom_array(13596);
		when "0011010100011101" => data_out <= rom_array(13597);
		when "0011010100011110" => data_out <= rom_array(13598);
		when "0011010100011111" => data_out <= rom_array(13599);
		when "0011010100100000" => data_out <= rom_array(13600);
		when "0011010100100001" => data_out <= rom_array(13601);
		when "0011010100100010" => data_out <= rom_array(13602);
		when "0011010100100011" => data_out <= rom_array(13603);
		when "0011010100100100" => data_out <= rom_array(13604);
		when "0011010100100101" => data_out <= rom_array(13605);
		when "0011010100100110" => data_out <= rom_array(13606);
		when "0011010100100111" => data_out <= rom_array(13607);
		when "0011010100101000" => data_out <= rom_array(13608);
		when "0011010100101001" => data_out <= rom_array(13609);
		when "0011010100101010" => data_out <= rom_array(13610);
		when "0011010100101011" => data_out <= rom_array(13611);
		when "0011010100101100" => data_out <= rom_array(13612);
		when "0011010100101101" => data_out <= rom_array(13613);
		when "0011010100101110" => data_out <= rom_array(13614);
		when "0011010100101111" => data_out <= rom_array(13615);
		when "0011010100110000" => data_out <= rom_array(13616);
		when "0011010100110001" => data_out <= rom_array(13617);
		when "0011010100110010" => data_out <= rom_array(13618);
		when "0011010100110011" => data_out <= rom_array(13619);
		when "0011010100110100" => data_out <= rom_array(13620);
		when "0011010100110101" => data_out <= rom_array(13621);
		when "0011010100110110" => data_out <= rom_array(13622);
		when "0011010100110111" => data_out <= rom_array(13623);
		when "0011010100111000" => data_out <= rom_array(13624);
		when "0011010100111001" => data_out <= rom_array(13625);
		when "0011010100111010" => data_out <= rom_array(13626);
		when "0011010100111011" => data_out <= rom_array(13627);
		when "0011010100111100" => data_out <= rom_array(13628);
		when "0011010100111101" => data_out <= rom_array(13629);
		when "0011010100111110" => data_out <= rom_array(13630);
		when "0011010100111111" => data_out <= rom_array(13631);
		when "0011010101000000" => data_out <= rom_array(13632);
		when "0011010101000001" => data_out <= rom_array(13633);
		when "0011010101000010" => data_out <= rom_array(13634);
		when "0011010101000011" => data_out <= rom_array(13635);
		when "0011010101000100" => data_out <= rom_array(13636);
		when "0011010101000101" => data_out <= rom_array(13637);
		when "0011010101000110" => data_out <= rom_array(13638);
		when "0011010101000111" => data_out <= rom_array(13639);
		when "0011010101001000" => data_out <= rom_array(13640);
		when "0011010101001001" => data_out <= rom_array(13641);
		when "0011010101001010" => data_out <= rom_array(13642);
		when "0011010101001011" => data_out <= rom_array(13643);
		when "0011010101001100" => data_out <= rom_array(13644);
		when "0011010101001101" => data_out <= rom_array(13645);
		when "0011010101001110" => data_out <= rom_array(13646);
		when "0011010101001111" => data_out <= rom_array(13647);
		when "0011010101010000" => data_out <= rom_array(13648);
		when "0011010101010001" => data_out <= rom_array(13649);
		when "0011010101010010" => data_out <= rom_array(13650);
		when "0011010101010011" => data_out <= rom_array(13651);
		when "0011010101010100" => data_out <= rom_array(13652);
		when "0011010101010101" => data_out <= rom_array(13653);
		when "0011010101010110" => data_out <= rom_array(13654);
		when "0011010101010111" => data_out <= rom_array(13655);
		when "0011010101011000" => data_out <= rom_array(13656);
		when "0011010101011001" => data_out <= rom_array(13657);
		when "0011010101011010" => data_out <= rom_array(13658);
		when "0011010101011011" => data_out <= rom_array(13659);
		when "0011010101011100" => data_out <= rom_array(13660);
		when "0011010101011101" => data_out <= rom_array(13661);
		when "0011010101011110" => data_out <= rom_array(13662);
		when "0011010101011111" => data_out <= rom_array(13663);
		when "0011010101100000" => data_out <= rom_array(13664);
		when "0011010101100001" => data_out <= rom_array(13665);
		when "0011010101100010" => data_out <= rom_array(13666);
		when "0011010101100011" => data_out <= rom_array(13667);
		when "0011010101100100" => data_out <= rom_array(13668);
		when "0011010101100101" => data_out <= rom_array(13669);
		when "0011010101100110" => data_out <= rom_array(13670);
		when "0011010101100111" => data_out <= rom_array(13671);
		when "0011010101101000" => data_out <= rom_array(13672);
		when "0011010101101001" => data_out <= rom_array(13673);
		when "0011010101101010" => data_out <= rom_array(13674);
		when "0011010101101011" => data_out <= rom_array(13675);
		when "0011010101101100" => data_out <= rom_array(13676);
		when "0011010101101101" => data_out <= rom_array(13677);
		when "0011010101101110" => data_out <= rom_array(13678);
		when "0011010101101111" => data_out <= rom_array(13679);
		when "0011010101110000" => data_out <= rom_array(13680);
		when "0011010101110001" => data_out <= rom_array(13681);
		when "0011010101110010" => data_out <= rom_array(13682);
		when "0011010101110011" => data_out <= rom_array(13683);
		when "0011010101110100" => data_out <= rom_array(13684);
		when "0011010101110101" => data_out <= rom_array(13685);
		when "0011010101110110" => data_out <= rom_array(13686);
		when "0011010101110111" => data_out <= rom_array(13687);
		when "0011010101111000" => data_out <= rom_array(13688);
		when "0011010101111001" => data_out <= rom_array(13689);
		when "0011010101111010" => data_out <= rom_array(13690);
		when "0011010101111011" => data_out <= rom_array(13691);
		when "0011010101111100" => data_out <= rom_array(13692);
		when "0011010101111101" => data_out <= rom_array(13693);
		when "0011010101111110" => data_out <= rom_array(13694);
		when "0011010101111111" => data_out <= rom_array(13695);
		when "0011010110000000" => data_out <= rom_array(13696);
		when "0011010110000001" => data_out <= rom_array(13697);
		when "0011010110000010" => data_out <= rom_array(13698);
		when "0011010110000011" => data_out <= rom_array(13699);
		when "0011010110000100" => data_out <= rom_array(13700);
		when "0011010110000101" => data_out <= rom_array(13701);
		when "0011010110000110" => data_out <= rom_array(13702);
		when "0011010110000111" => data_out <= rom_array(13703);
		when "0011010110001000" => data_out <= rom_array(13704);
		when "0011010110001001" => data_out <= rom_array(13705);
		when "0011010110001010" => data_out <= rom_array(13706);
		when "0011010110001011" => data_out <= rom_array(13707);
		when "0011010110001100" => data_out <= rom_array(13708);
		when "0011010110001101" => data_out <= rom_array(13709);
		when "0011010110001110" => data_out <= rom_array(13710);
		when "0011010110001111" => data_out <= rom_array(13711);
		when "0011010110010000" => data_out <= rom_array(13712);
		when "0011010110010001" => data_out <= rom_array(13713);
		when "0011010110010010" => data_out <= rom_array(13714);
		when "0011010110010011" => data_out <= rom_array(13715);
		when "0011010110010100" => data_out <= rom_array(13716);
		when "0011010110010101" => data_out <= rom_array(13717);
		when "0011010110010110" => data_out <= rom_array(13718);
		when "0011010110010111" => data_out <= rom_array(13719);
		when "0011010110011000" => data_out <= rom_array(13720);
		when "0011010110011001" => data_out <= rom_array(13721);
		when "0011010110011010" => data_out <= rom_array(13722);
		when "0011010110011011" => data_out <= rom_array(13723);
		when "0011010110011100" => data_out <= rom_array(13724);
		when "0011010110011101" => data_out <= rom_array(13725);
		when "0011010110011110" => data_out <= rom_array(13726);
		when "0011010110011111" => data_out <= rom_array(13727);
		when "0011010110100000" => data_out <= rom_array(13728);
		when "0011010110100001" => data_out <= rom_array(13729);
		when "0011010110100010" => data_out <= rom_array(13730);
		when "0011010110100011" => data_out <= rom_array(13731);
		when "0011010110100100" => data_out <= rom_array(13732);
		when "0011010110100101" => data_out <= rom_array(13733);
		when "0011010110100110" => data_out <= rom_array(13734);
		when "0011010110100111" => data_out <= rom_array(13735);
		when "0011010110101000" => data_out <= rom_array(13736);
		when "0011010110101001" => data_out <= rom_array(13737);
		when "0011010110101010" => data_out <= rom_array(13738);
		when "0011010110101011" => data_out <= rom_array(13739);
		when "0011010110101100" => data_out <= rom_array(13740);
		when "0011010110101101" => data_out <= rom_array(13741);
		when "0011010110101110" => data_out <= rom_array(13742);
		when "0011010110101111" => data_out <= rom_array(13743);
		when "0011010110110000" => data_out <= rom_array(13744);
		when "0011010110110001" => data_out <= rom_array(13745);
		when "0011010110110010" => data_out <= rom_array(13746);
		when "0011010110110011" => data_out <= rom_array(13747);
		when "0011010110110100" => data_out <= rom_array(13748);
		when "0011010110110101" => data_out <= rom_array(13749);
		when "0011010110110110" => data_out <= rom_array(13750);
		when "0011010110110111" => data_out <= rom_array(13751);
		when "0011010110111000" => data_out <= rom_array(13752);
		when "0011010110111001" => data_out <= rom_array(13753);
		when "0011010110111010" => data_out <= rom_array(13754);
		when "0011010110111011" => data_out <= rom_array(13755);
		when "0011010110111100" => data_out <= rom_array(13756);
		when "0011010110111101" => data_out <= rom_array(13757);
		when "0011010110111110" => data_out <= rom_array(13758);
		when "0011010110111111" => data_out <= rom_array(13759);
		when "0011010111000000" => data_out <= rom_array(13760);
		when "0011010111000001" => data_out <= rom_array(13761);
		when "0011010111000010" => data_out <= rom_array(13762);
		when "0011010111000011" => data_out <= rom_array(13763);
		when "0011010111000100" => data_out <= rom_array(13764);
		when "0011010111000101" => data_out <= rom_array(13765);
		when "0011010111000110" => data_out <= rom_array(13766);
		when "0011010111000111" => data_out <= rom_array(13767);
		when "0011010111001000" => data_out <= rom_array(13768);
		when "0011010111001001" => data_out <= rom_array(13769);
		when "0011010111001010" => data_out <= rom_array(13770);
		when "0011010111001011" => data_out <= rom_array(13771);
		when "0011010111001100" => data_out <= rom_array(13772);
		when "0011010111001101" => data_out <= rom_array(13773);
		when "0011010111001110" => data_out <= rom_array(13774);
		when "0011010111001111" => data_out <= rom_array(13775);
		when "0011010111010000" => data_out <= rom_array(13776);
		when "0011010111010001" => data_out <= rom_array(13777);
		when "0011010111010010" => data_out <= rom_array(13778);
		when "0011010111010011" => data_out <= rom_array(13779);
		when "0011010111010100" => data_out <= rom_array(13780);
		when "0011010111010101" => data_out <= rom_array(13781);
		when "0011010111010110" => data_out <= rom_array(13782);
		when "0011010111010111" => data_out <= rom_array(13783);
		when "0011010111011000" => data_out <= rom_array(13784);
		when "0011010111011001" => data_out <= rom_array(13785);
		when "0011010111011010" => data_out <= rom_array(13786);
		when "0011010111011011" => data_out <= rom_array(13787);
		when "0011010111011100" => data_out <= rom_array(13788);
		when "0011010111011101" => data_out <= rom_array(13789);
		when "0011010111011110" => data_out <= rom_array(13790);
		when "0011010111011111" => data_out <= rom_array(13791);
		when "0011010111100000" => data_out <= rom_array(13792);
		when "0011010111100001" => data_out <= rom_array(13793);
		when "0011010111100010" => data_out <= rom_array(13794);
		when "0011010111100011" => data_out <= rom_array(13795);
		when "0011010111100100" => data_out <= rom_array(13796);
		when "0011010111100101" => data_out <= rom_array(13797);
		when "0011010111100110" => data_out <= rom_array(13798);
		when "0011010111100111" => data_out <= rom_array(13799);
		when "0011010111101000" => data_out <= rom_array(13800);
		when "0011010111101001" => data_out <= rom_array(13801);
		when "0011010111101010" => data_out <= rom_array(13802);
		when "0011010111101011" => data_out <= rom_array(13803);
		when "0011010111101100" => data_out <= rom_array(13804);
		when "0011010111101101" => data_out <= rom_array(13805);
		when "0011010111101110" => data_out <= rom_array(13806);
		when "0011010111101111" => data_out <= rom_array(13807);
		when "0011010111110000" => data_out <= rom_array(13808);
		when "0011010111110001" => data_out <= rom_array(13809);
		when "0011010111110010" => data_out <= rom_array(13810);
		when "0011010111110011" => data_out <= rom_array(13811);
		when "0011010111110100" => data_out <= rom_array(13812);
		when "0011010111110101" => data_out <= rom_array(13813);
		when "0011010111110110" => data_out <= rom_array(13814);
		when "0011010111110111" => data_out <= rom_array(13815);
		when "0011010111111000" => data_out <= rom_array(13816);
		when "0011010111111001" => data_out <= rom_array(13817);
		when "0011010111111010" => data_out <= rom_array(13818);
		when "0011010111111011" => data_out <= rom_array(13819);
		when "0011010111111100" => data_out <= rom_array(13820);
		when "0011010111111101" => data_out <= rom_array(13821);
		when "0011010111111110" => data_out <= rom_array(13822);
		when "0011010111111111" => data_out <= rom_array(13823);
		when "0011011000000000" => data_out <= rom_array(13824);
		when "0011011000000001" => data_out <= rom_array(13825);
		when "0011011000000010" => data_out <= rom_array(13826);
		when "0011011000000011" => data_out <= rom_array(13827);
		when "0011011000000100" => data_out <= rom_array(13828);
		when "0011011000000101" => data_out <= rom_array(13829);
		when "0011011000000110" => data_out <= rom_array(13830);
		when "0011011000000111" => data_out <= rom_array(13831);
		when "0011011000001000" => data_out <= rom_array(13832);
		when "0011011000001001" => data_out <= rom_array(13833);
		when "0011011000001010" => data_out <= rom_array(13834);
		when "0011011000001011" => data_out <= rom_array(13835);
		when "0011011000001100" => data_out <= rom_array(13836);
		when "0011011000001101" => data_out <= rom_array(13837);
		when "0011011000001110" => data_out <= rom_array(13838);
		when "0011011000001111" => data_out <= rom_array(13839);
		when "0011011000010000" => data_out <= rom_array(13840);
		when "0011011000010001" => data_out <= rom_array(13841);
		when "0011011000010010" => data_out <= rom_array(13842);
		when "0011011000010011" => data_out <= rom_array(13843);
		when "0011011000010100" => data_out <= rom_array(13844);
		when "0011011000010101" => data_out <= rom_array(13845);
		when "0011011000010110" => data_out <= rom_array(13846);
		when "0011011000010111" => data_out <= rom_array(13847);
		when "0011011000011000" => data_out <= rom_array(13848);
		when "0011011000011001" => data_out <= rom_array(13849);
		when "0011011000011010" => data_out <= rom_array(13850);
		when "0011011000011011" => data_out <= rom_array(13851);
		when "0011011000011100" => data_out <= rom_array(13852);
		when "0011011000011101" => data_out <= rom_array(13853);
		when "0011011000011110" => data_out <= rom_array(13854);
		when "0011011000011111" => data_out <= rom_array(13855);
		when "0011011000100000" => data_out <= rom_array(13856);
		when "0011011000100001" => data_out <= rom_array(13857);
		when "0011011000100010" => data_out <= rom_array(13858);
		when "0011011000100011" => data_out <= rom_array(13859);
		when "0011011000100100" => data_out <= rom_array(13860);
		when "0011011000100101" => data_out <= rom_array(13861);
		when "0011011000100110" => data_out <= rom_array(13862);
		when "0011011000100111" => data_out <= rom_array(13863);
		when "0011011000101000" => data_out <= rom_array(13864);
		when "0011011000101001" => data_out <= rom_array(13865);
		when "0011011000101010" => data_out <= rom_array(13866);
		when "0011011000101011" => data_out <= rom_array(13867);
		when "0011011000101100" => data_out <= rom_array(13868);
		when "0011011000101101" => data_out <= rom_array(13869);
		when "0011011000101110" => data_out <= rom_array(13870);
		when "0011011000101111" => data_out <= rom_array(13871);
		when "0011011000110000" => data_out <= rom_array(13872);
		when "0011011000110001" => data_out <= rom_array(13873);
		when "0011011000110010" => data_out <= rom_array(13874);
		when "0011011000110011" => data_out <= rom_array(13875);
		when "0011011000110100" => data_out <= rom_array(13876);
		when "0011011000110101" => data_out <= rom_array(13877);
		when "0011011000110110" => data_out <= rom_array(13878);
		when "0011011000110111" => data_out <= rom_array(13879);
		when "0011011000111000" => data_out <= rom_array(13880);
		when "0011011000111001" => data_out <= rom_array(13881);
		when "0011011000111010" => data_out <= rom_array(13882);
		when "0011011000111011" => data_out <= rom_array(13883);
		when "0011011000111100" => data_out <= rom_array(13884);
		when "0011011000111101" => data_out <= rom_array(13885);
		when "0011011000111110" => data_out <= rom_array(13886);
		when "0011011000111111" => data_out <= rom_array(13887);
		when "0011011001000000" => data_out <= rom_array(13888);
		when "0011011001000001" => data_out <= rom_array(13889);
		when "0011011001000010" => data_out <= rom_array(13890);
		when "0011011001000011" => data_out <= rom_array(13891);
		when "0011011001000100" => data_out <= rom_array(13892);
		when "0011011001000101" => data_out <= rom_array(13893);
		when "0011011001000110" => data_out <= rom_array(13894);
		when "0011011001000111" => data_out <= rom_array(13895);
		when "0011011001001000" => data_out <= rom_array(13896);
		when "0011011001001001" => data_out <= rom_array(13897);
		when "0011011001001010" => data_out <= rom_array(13898);
		when "0011011001001011" => data_out <= rom_array(13899);
		when "0011011001001100" => data_out <= rom_array(13900);
		when "0011011001001101" => data_out <= rom_array(13901);
		when "0011011001001110" => data_out <= rom_array(13902);
		when "0011011001001111" => data_out <= rom_array(13903);
		when "0011011001010000" => data_out <= rom_array(13904);
		when "0011011001010001" => data_out <= rom_array(13905);
		when "0011011001010010" => data_out <= rom_array(13906);
		when "0011011001010011" => data_out <= rom_array(13907);
		when "0011011001010100" => data_out <= rom_array(13908);
		when "0011011001010101" => data_out <= rom_array(13909);
		when "0011011001010110" => data_out <= rom_array(13910);
		when "0011011001010111" => data_out <= rom_array(13911);
		when "0011011001011000" => data_out <= rom_array(13912);
		when "0011011001011001" => data_out <= rom_array(13913);
		when "0011011001011010" => data_out <= rom_array(13914);
		when "0011011001011011" => data_out <= rom_array(13915);
		when "0011011001011100" => data_out <= rom_array(13916);
		when "0011011001011101" => data_out <= rom_array(13917);
		when "0011011001011110" => data_out <= rom_array(13918);
		when "0011011001011111" => data_out <= rom_array(13919);
		when "0011011001100000" => data_out <= rom_array(13920);
		when "0011011001100001" => data_out <= rom_array(13921);
		when "0011011001100010" => data_out <= rom_array(13922);
		when "0011011001100011" => data_out <= rom_array(13923);
		when "0011011001100100" => data_out <= rom_array(13924);
		when "0011011001100101" => data_out <= rom_array(13925);
		when "0011011001100110" => data_out <= rom_array(13926);
		when "0011011001100111" => data_out <= rom_array(13927);
		when "0011011001101000" => data_out <= rom_array(13928);
		when "0011011001101001" => data_out <= rom_array(13929);
		when "0011011001101010" => data_out <= rom_array(13930);
		when "0011011001101011" => data_out <= rom_array(13931);
		when "0011011001101100" => data_out <= rom_array(13932);
		when "0011011001101101" => data_out <= rom_array(13933);
		when "0011011001101110" => data_out <= rom_array(13934);
		when "0011011001101111" => data_out <= rom_array(13935);
		when "0011011001110000" => data_out <= rom_array(13936);
		when "0011011001110001" => data_out <= rom_array(13937);
		when "0011011001110010" => data_out <= rom_array(13938);
		when "0011011001110011" => data_out <= rom_array(13939);
		when "0011011001110100" => data_out <= rom_array(13940);
		when "0011011001110101" => data_out <= rom_array(13941);
		when "0011011001110110" => data_out <= rom_array(13942);
		when "0011011001110111" => data_out <= rom_array(13943);
		when "0011011001111000" => data_out <= rom_array(13944);
		when "0011011001111001" => data_out <= rom_array(13945);
		when "0011011001111010" => data_out <= rom_array(13946);
		when "0011011001111011" => data_out <= rom_array(13947);
		when "0011011001111100" => data_out <= rom_array(13948);
		when "0011011001111101" => data_out <= rom_array(13949);
		when "0011011001111110" => data_out <= rom_array(13950);
		when "0011011001111111" => data_out <= rom_array(13951);
		when "0011011010000000" => data_out <= rom_array(13952);
		when "0011011010000001" => data_out <= rom_array(13953);
		when "0011011010000010" => data_out <= rom_array(13954);
		when "0011011010000011" => data_out <= rom_array(13955);
		when "0011011010000100" => data_out <= rom_array(13956);
		when "0011011010000101" => data_out <= rom_array(13957);
		when "0011011010000110" => data_out <= rom_array(13958);
		when "0011011010000111" => data_out <= rom_array(13959);
		when "0011011010001000" => data_out <= rom_array(13960);
		when "0011011010001001" => data_out <= rom_array(13961);
		when "0011011010001010" => data_out <= rom_array(13962);
		when "0011011010001011" => data_out <= rom_array(13963);
		when "0011011010001100" => data_out <= rom_array(13964);
		when "0011011010001101" => data_out <= rom_array(13965);
		when "0011011010001110" => data_out <= rom_array(13966);
		when "0011011010001111" => data_out <= rom_array(13967);
		when "0011011010010000" => data_out <= rom_array(13968);
		when "0011011010010001" => data_out <= rom_array(13969);
		when "0011011010010010" => data_out <= rom_array(13970);
		when "0011011010010011" => data_out <= rom_array(13971);
		when "0011011010010100" => data_out <= rom_array(13972);
		when "0011011010010101" => data_out <= rom_array(13973);
		when "0011011010010110" => data_out <= rom_array(13974);
		when "0011011010010111" => data_out <= rom_array(13975);
		when "0011011010011000" => data_out <= rom_array(13976);
		when "0011011010011001" => data_out <= rom_array(13977);
		when "0011011010011010" => data_out <= rom_array(13978);
		when "0011011010011011" => data_out <= rom_array(13979);
		when "0011011010011100" => data_out <= rom_array(13980);
		when "0011011010011101" => data_out <= rom_array(13981);
		when "0011011010011110" => data_out <= rom_array(13982);
		when "0011011010011111" => data_out <= rom_array(13983);
		when "0011011010100000" => data_out <= rom_array(13984);
		when "0011011010100001" => data_out <= rom_array(13985);
		when "0011011010100010" => data_out <= rom_array(13986);
		when "0011011010100011" => data_out <= rom_array(13987);
		when "0011011010100100" => data_out <= rom_array(13988);
		when "0011011010100101" => data_out <= rom_array(13989);
		when "0011011010100110" => data_out <= rom_array(13990);
		when "0011011010100111" => data_out <= rom_array(13991);
		when "0011011010101000" => data_out <= rom_array(13992);
		when "0011011010101001" => data_out <= rom_array(13993);
		when "0011011010101010" => data_out <= rom_array(13994);
		when "0011011010101011" => data_out <= rom_array(13995);
		when "0011011010101100" => data_out <= rom_array(13996);
		when "0011011010101101" => data_out <= rom_array(13997);
		when "0011011010101110" => data_out <= rom_array(13998);
		when "0011011010101111" => data_out <= rom_array(13999);
		when "0011011010110000" => data_out <= rom_array(14000);
		when "0011011010110001" => data_out <= rom_array(14001);
		when "0011011010110010" => data_out <= rom_array(14002);
		when "0011011010110011" => data_out <= rom_array(14003);
		when "0011011010110100" => data_out <= rom_array(14004);
		when "0011011010110101" => data_out <= rom_array(14005);
		when "0011011010110110" => data_out <= rom_array(14006);
		when "0011011010110111" => data_out <= rom_array(14007);
		when "0011011010111000" => data_out <= rom_array(14008);
		when "0011011010111001" => data_out <= rom_array(14009);
		when "0011011010111010" => data_out <= rom_array(14010);
		when "0011011010111011" => data_out <= rom_array(14011);
		when "0011011010111100" => data_out <= rom_array(14012);
		when "0011011010111101" => data_out <= rom_array(14013);
		when "0011011010111110" => data_out <= rom_array(14014);
		when "0011011010111111" => data_out <= rom_array(14015);
		when "0011011011000000" => data_out <= rom_array(14016);
		when "0011011011000001" => data_out <= rom_array(14017);
		when "0011011011000010" => data_out <= rom_array(14018);
		when "0011011011000011" => data_out <= rom_array(14019);
		when "0011011011000100" => data_out <= rom_array(14020);
		when "0011011011000101" => data_out <= rom_array(14021);
		when "0011011011000110" => data_out <= rom_array(14022);
		when "0011011011000111" => data_out <= rom_array(14023);
		when "0011011011001000" => data_out <= rom_array(14024);
		when "0011011011001001" => data_out <= rom_array(14025);
		when "0011011011001010" => data_out <= rom_array(14026);
		when "0011011011001011" => data_out <= rom_array(14027);
		when "0011011011001100" => data_out <= rom_array(14028);
		when "0011011011001101" => data_out <= rom_array(14029);
		when "0011011011001110" => data_out <= rom_array(14030);
		when "0011011011001111" => data_out <= rom_array(14031);
		when "0011011011010000" => data_out <= rom_array(14032);
		when "0011011011010001" => data_out <= rom_array(14033);
		when "0011011011010010" => data_out <= rom_array(14034);
		when "0011011011010011" => data_out <= rom_array(14035);
		when "0011011011010100" => data_out <= rom_array(14036);
		when "0011011011010101" => data_out <= rom_array(14037);
		when "0011011011010110" => data_out <= rom_array(14038);
		when "0011011011010111" => data_out <= rom_array(14039);
		when "0011011011011000" => data_out <= rom_array(14040);
		when "0011011011011001" => data_out <= rom_array(14041);
		when "0011011011011010" => data_out <= rom_array(14042);
		when "0011011011011011" => data_out <= rom_array(14043);
		when "0011011011011100" => data_out <= rom_array(14044);
		when "0011011011011101" => data_out <= rom_array(14045);
		when "0011011011011110" => data_out <= rom_array(14046);
		when "0011011011011111" => data_out <= rom_array(14047);
		when "0011011011100000" => data_out <= rom_array(14048);
		when "0011011011100001" => data_out <= rom_array(14049);
		when "0011011011100010" => data_out <= rom_array(14050);
		when "0011011011100011" => data_out <= rom_array(14051);
		when "0011011011100100" => data_out <= rom_array(14052);
		when "0011011011100101" => data_out <= rom_array(14053);
		when "0011011011100110" => data_out <= rom_array(14054);
		when "0011011011100111" => data_out <= rom_array(14055);
		when "0011011011101000" => data_out <= rom_array(14056);
		when "0011011011101001" => data_out <= rom_array(14057);
		when "0011011011101010" => data_out <= rom_array(14058);
		when "0011011011101011" => data_out <= rom_array(14059);
		when "0011011011101100" => data_out <= rom_array(14060);
		when "0011011011101101" => data_out <= rom_array(14061);
		when "0011011011101110" => data_out <= rom_array(14062);
		when "0011011011101111" => data_out <= rom_array(14063);
		when "0011011011110000" => data_out <= rom_array(14064);
		when "0011011011110001" => data_out <= rom_array(14065);
		when "0011011011110010" => data_out <= rom_array(14066);
		when "0011011011110011" => data_out <= rom_array(14067);
		when "0011011011110100" => data_out <= rom_array(14068);
		when "0011011011110101" => data_out <= rom_array(14069);
		when "0011011011110110" => data_out <= rom_array(14070);
		when "0011011011110111" => data_out <= rom_array(14071);
		when "0011011011111000" => data_out <= rom_array(14072);
		when "0011011011111001" => data_out <= rom_array(14073);
		when "0011011011111010" => data_out <= rom_array(14074);
		when "0011011011111011" => data_out <= rom_array(14075);
		when "0011011011111100" => data_out <= rom_array(14076);
		when "0011011011111101" => data_out <= rom_array(14077);
		when "0011011011111110" => data_out <= rom_array(14078);
		when "0011011011111111" => data_out <= rom_array(14079);
		when "0011011100000000" => data_out <= rom_array(14080);
		when "0011011100000001" => data_out <= rom_array(14081);
		when "0011011100000010" => data_out <= rom_array(14082);
		when "0011011100000011" => data_out <= rom_array(14083);
		when "0011011100000100" => data_out <= rom_array(14084);
		when "0011011100000101" => data_out <= rom_array(14085);
		when "0011011100000110" => data_out <= rom_array(14086);
		when "0011011100000111" => data_out <= rom_array(14087);
		when "0011011100001000" => data_out <= rom_array(14088);
		when "0011011100001001" => data_out <= rom_array(14089);
		when "0011011100001010" => data_out <= rom_array(14090);
		when "0011011100001011" => data_out <= rom_array(14091);
		when "0011011100001100" => data_out <= rom_array(14092);
		when "0011011100001101" => data_out <= rom_array(14093);
		when "0011011100001110" => data_out <= rom_array(14094);
		when "0011011100001111" => data_out <= rom_array(14095);
		when "0011011100010000" => data_out <= rom_array(14096);
		when "0011011100010001" => data_out <= rom_array(14097);
		when "0011011100010010" => data_out <= rom_array(14098);
		when "0011011100010011" => data_out <= rom_array(14099);
		when "0011011100010100" => data_out <= rom_array(14100);
		when "0011011100010101" => data_out <= rom_array(14101);
		when "0011011100010110" => data_out <= rom_array(14102);
		when "0011011100010111" => data_out <= rom_array(14103);
		when "0011011100011000" => data_out <= rom_array(14104);
		when "0011011100011001" => data_out <= rom_array(14105);
		when "0011011100011010" => data_out <= rom_array(14106);
		when "0011011100011011" => data_out <= rom_array(14107);
		when "0011011100011100" => data_out <= rom_array(14108);
		when "0011011100011101" => data_out <= rom_array(14109);
		when "0011011100011110" => data_out <= rom_array(14110);
		when "0011011100011111" => data_out <= rom_array(14111);
		when "0011011100100000" => data_out <= rom_array(14112);
		when "0011011100100001" => data_out <= rom_array(14113);
		when "0011011100100010" => data_out <= rom_array(14114);
		when "0011011100100011" => data_out <= rom_array(14115);
		when "0011011100100100" => data_out <= rom_array(14116);
		when "0011011100100101" => data_out <= rom_array(14117);
		when "0011011100100110" => data_out <= rom_array(14118);
		when "0011011100100111" => data_out <= rom_array(14119);
		when "0011011100101000" => data_out <= rom_array(14120);
		when "0011011100101001" => data_out <= rom_array(14121);
		when "0011011100101010" => data_out <= rom_array(14122);
		when "0011011100101011" => data_out <= rom_array(14123);
		when "0011011100101100" => data_out <= rom_array(14124);
		when "0011011100101101" => data_out <= rom_array(14125);
		when "0011011100101110" => data_out <= rom_array(14126);
		when "0011011100101111" => data_out <= rom_array(14127);
		when "0011011100110000" => data_out <= rom_array(14128);
		when "0011011100110001" => data_out <= rom_array(14129);
		when "0011011100110010" => data_out <= rom_array(14130);
		when "0011011100110011" => data_out <= rom_array(14131);
		when "0011011100110100" => data_out <= rom_array(14132);
		when "0011011100110101" => data_out <= rom_array(14133);
		when "0011011100110110" => data_out <= rom_array(14134);
		when "0011011100110111" => data_out <= rom_array(14135);
		when "0011011100111000" => data_out <= rom_array(14136);
		when "0011011100111001" => data_out <= rom_array(14137);
		when "0011011100111010" => data_out <= rom_array(14138);
		when "0011011100111011" => data_out <= rom_array(14139);
		when "0011011100111100" => data_out <= rom_array(14140);
		when "0011011100111101" => data_out <= rom_array(14141);
		when "0011011100111110" => data_out <= rom_array(14142);
		when "0011011100111111" => data_out <= rom_array(14143);
		when "0011011101000000" => data_out <= rom_array(14144);
		when "0011011101000001" => data_out <= rom_array(14145);
		when "0011011101000010" => data_out <= rom_array(14146);
		when "0011011101000011" => data_out <= rom_array(14147);
		when "0011011101000100" => data_out <= rom_array(14148);
		when "0011011101000101" => data_out <= rom_array(14149);
		when "0011011101000110" => data_out <= rom_array(14150);
		when "0011011101000111" => data_out <= rom_array(14151);
		when "0011011101001000" => data_out <= rom_array(14152);
		when "0011011101001001" => data_out <= rom_array(14153);
		when "0011011101001010" => data_out <= rom_array(14154);
		when "0011011101001011" => data_out <= rom_array(14155);
		when "0011011101001100" => data_out <= rom_array(14156);
		when "0011011101001101" => data_out <= rom_array(14157);
		when "0011011101001110" => data_out <= rom_array(14158);
		when "0011011101001111" => data_out <= rom_array(14159);
		when "0011011101010000" => data_out <= rom_array(14160);
		when "0011011101010001" => data_out <= rom_array(14161);
		when "0011011101010010" => data_out <= rom_array(14162);
		when "0011011101010011" => data_out <= rom_array(14163);
		when "0011011101010100" => data_out <= rom_array(14164);
		when "0011011101010101" => data_out <= rom_array(14165);
		when "0011011101010110" => data_out <= rom_array(14166);
		when "0011011101010111" => data_out <= rom_array(14167);
		when "0011011101011000" => data_out <= rom_array(14168);
		when "0011011101011001" => data_out <= rom_array(14169);
		when "0011011101011010" => data_out <= rom_array(14170);
		when "0011011101011011" => data_out <= rom_array(14171);
		when "0011011101011100" => data_out <= rom_array(14172);
		when "0011011101011101" => data_out <= rom_array(14173);
		when "0011011101011110" => data_out <= rom_array(14174);
		when "0011011101011111" => data_out <= rom_array(14175);
		when "0011011101100000" => data_out <= rom_array(14176);
		when "0011011101100001" => data_out <= rom_array(14177);
		when "0011011101100010" => data_out <= rom_array(14178);
		when "0011011101100011" => data_out <= rom_array(14179);
		when "0011011101100100" => data_out <= rom_array(14180);
		when "0011011101100101" => data_out <= rom_array(14181);
		when "0011011101100110" => data_out <= rom_array(14182);
		when "0011011101100111" => data_out <= rom_array(14183);
		when "0011011101101000" => data_out <= rom_array(14184);
		when "0011011101101001" => data_out <= rom_array(14185);
		when "0011011101101010" => data_out <= rom_array(14186);
		when "0011011101101011" => data_out <= rom_array(14187);
		when "0011011101101100" => data_out <= rom_array(14188);
		when "0011011101101101" => data_out <= rom_array(14189);
		when "0011011101101110" => data_out <= rom_array(14190);
		when "0011011101101111" => data_out <= rom_array(14191);
		when "0011011101110000" => data_out <= rom_array(14192);
		when "0011011101110001" => data_out <= rom_array(14193);
		when "0011011101110010" => data_out <= rom_array(14194);
		when "0011011101110011" => data_out <= rom_array(14195);
		when "0011011101110100" => data_out <= rom_array(14196);
		when "0011011101110101" => data_out <= rom_array(14197);
		when "0011011101110110" => data_out <= rom_array(14198);
		when "0011011101110111" => data_out <= rom_array(14199);
		when "0011011101111000" => data_out <= rom_array(14200);
		when "0011011101111001" => data_out <= rom_array(14201);
		when "0011011101111010" => data_out <= rom_array(14202);
		when "0011011101111011" => data_out <= rom_array(14203);
		when "0011011101111100" => data_out <= rom_array(14204);
		when "0011011101111101" => data_out <= rom_array(14205);
		when "0011011101111110" => data_out <= rom_array(14206);
		when "0011011101111111" => data_out <= rom_array(14207);
		when "0011011110000000" => data_out <= rom_array(14208);
		when "0011011110000001" => data_out <= rom_array(14209);
		when "0011011110000010" => data_out <= rom_array(14210);
		when "0011011110000011" => data_out <= rom_array(14211);
		when "0011011110000100" => data_out <= rom_array(14212);
		when "0011011110000101" => data_out <= rom_array(14213);
		when "0011011110000110" => data_out <= rom_array(14214);
		when "0011011110000111" => data_out <= rom_array(14215);
		when "0011011110001000" => data_out <= rom_array(14216);
		when "0011011110001001" => data_out <= rom_array(14217);
		when "0011011110001010" => data_out <= rom_array(14218);
		when "0011011110001011" => data_out <= rom_array(14219);
		when "0011011110001100" => data_out <= rom_array(14220);
		when "0011011110001101" => data_out <= rom_array(14221);
		when "0011011110001110" => data_out <= rom_array(14222);
		when "0011011110001111" => data_out <= rom_array(14223);
		when "0011011110010000" => data_out <= rom_array(14224);
		when "0011011110010001" => data_out <= rom_array(14225);
		when "0011011110010010" => data_out <= rom_array(14226);
		when "0011011110010011" => data_out <= rom_array(14227);
		when "0011011110010100" => data_out <= rom_array(14228);
		when "0011011110010101" => data_out <= rom_array(14229);
		when "0011011110010110" => data_out <= rom_array(14230);
		when "0011011110010111" => data_out <= rom_array(14231);
		when "0011011110011000" => data_out <= rom_array(14232);
		when "0011011110011001" => data_out <= rom_array(14233);
		when "0011011110011010" => data_out <= rom_array(14234);
		when "0011011110011011" => data_out <= rom_array(14235);
		when "0011011110011100" => data_out <= rom_array(14236);
		when "0011011110011101" => data_out <= rom_array(14237);
		when "0011011110011110" => data_out <= rom_array(14238);
		when "0011011110011111" => data_out <= rom_array(14239);
		when "0011011110100000" => data_out <= rom_array(14240);
		when "0011011110100001" => data_out <= rom_array(14241);
		when "0011011110100010" => data_out <= rom_array(14242);
		when "0011011110100011" => data_out <= rom_array(14243);
		when "0011011110100100" => data_out <= rom_array(14244);
		when "0011011110100101" => data_out <= rom_array(14245);
		when "0011011110100110" => data_out <= rom_array(14246);
		when "0011011110100111" => data_out <= rom_array(14247);
		when "0011011110101000" => data_out <= rom_array(14248);
		when "0011011110101001" => data_out <= rom_array(14249);
		when "0011011110101010" => data_out <= rom_array(14250);
		when "0011011110101011" => data_out <= rom_array(14251);
		when "0011011110101100" => data_out <= rom_array(14252);
		when "0011011110101101" => data_out <= rom_array(14253);
		when "0011011110101110" => data_out <= rom_array(14254);
		when "0011011110101111" => data_out <= rom_array(14255);
		when "0011011110110000" => data_out <= rom_array(14256);
		when "0011011110110001" => data_out <= rom_array(14257);
		when "0011011110110010" => data_out <= rom_array(14258);
		when "0011011110110011" => data_out <= rom_array(14259);
		when "0011011110110100" => data_out <= rom_array(14260);
		when "0011011110110101" => data_out <= rom_array(14261);
		when "0011011110110110" => data_out <= rom_array(14262);
		when "0011011110110111" => data_out <= rom_array(14263);
		when "0011011110111000" => data_out <= rom_array(14264);
		when "0011011110111001" => data_out <= rom_array(14265);
		when "0011011110111010" => data_out <= rom_array(14266);
		when "0011011110111011" => data_out <= rom_array(14267);
		when "0011011110111100" => data_out <= rom_array(14268);
		when "0011011110111101" => data_out <= rom_array(14269);
		when "0011011110111110" => data_out <= rom_array(14270);
		when "0011011110111111" => data_out <= rom_array(14271);
		when "0011011111000000" => data_out <= rom_array(14272);
		when "0011011111000001" => data_out <= rom_array(14273);
		when "0011011111000010" => data_out <= rom_array(14274);
		when "0011011111000011" => data_out <= rom_array(14275);
		when "0011011111000100" => data_out <= rom_array(14276);
		when "0011011111000101" => data_out <= rom_array(14277);
		when "0011011111000110" => data_out <= rom_array(14278);
		when "0011011111000111" => data_out <= rom_array(14279);
		when "0011011111001000" => data_out <= rom_array(14280);
		when "0011011111001001" => data_out <= rom_array(14281);
		when "0011011111001010" => data_out <= rom_array(14282);
		when "0011011111001011" => data_out <= rom_array(14283);
		when "0011011111001100" => data_out <= rom_array(14284);
		when "0011011111001101" => data_out <= rom_array(14285);
		when "0011011111001110" => data_out <= rom_array(14286);
		when "0011011111001111" => data_out <= rom_array(14287);
		when "0011011111010000" => data_out <= rom_array(14288);
		when "0011011111010001" => data_out <= rom_array(14289);
		when "0011011111010010" => data_out <= rom_array(14290);
		when "0011011111010011" => data_out <= rom_array(14291);
		when "0011011111010100" => data_out <= rom_array(14292);
		when "0011011111010101" => data_out <= rom_array(14293);
		when "0011011111010110" => data_out <= rom_array(14294);
		when "0011011111010111" => data_out <= rom_array(14295);
		when "0011011111011000" => data_out <= rom_array(14296);
		when "0011011111011001" => data_out <= rom_array(14297);
		when "0011011111011010" => data_out <= rom_array(14298);
		when "0011011111011011" => data_out <= rom_array(14299);
		when "0011011111011100" => data_out <= rom_array(14300);
		when "0011011111011101" => data_out <= rom_array(14301);
		when "0011011111011110" => data_out <= rom_array(14302);
		when "0011011111011111" => data_out <= rom_array(14303);
		when "0011011111100000" => data_out <= rom_array(14304);
		when "0011011111100001" => data_out <= rom_array(14305);
		when "0011011111100010" => data_out <= rom_array(14306);
		when "0011011111100011" => data_out <= rom_array(14307);
		when "0011011111100100" => data_out <= rom_array(14308);
		when "0011011111100101" => data_out <= rom_array(14309);
		when "0011011111100110" => data_out <= rom_array(14310);
		when "0011011111100111" => data_out <= rom_array(14311);
		when "0011011111101000" => data_out <= rom_array(14312);
		when "0011011111101001" => data_out <= rom_array(14313);
		when "0011011111101010" => data_out <= rom_array(14314);
		when "0011011111101011" => data_out <= rom_array(14315);
		when "0011011111101100" => data_out <= rom_array(14316);
		when "0011011111101101" => data_out <= rom_array(14317);
		when "0011011111101110" => data_out <= rom_array(14318);
		when "0011011111101111" => data_out <= rom_array(14319);
		when "0011011111110000" => data_out <= rom_array(14320);
		when "0011011111110001" => data_out <= rom_array(14321);
		when "0011011111110010" => data_out <= rom_array(14322);
		when "0011011111110011" => data_out <= rom_array(14323);
		when "0011011111110100" => data_out <= rom_array(14324);
		when "0011011111110101" => data_out <= rom_array(14325);
		when "0011011111110110" => data_out <= rom_array(14326);
		when "0011011111110111" => data_out <= rom_array(14327);
		when "0011011111111000" => data_out <= rom_array(14328);
		when "0011011111111001" => data_out <= rom_array(14329);
		when "0011011111111010" => data_out <= rom_array(14330);
		when "0011011111111011" => data_out <= rom_array(14331);
		when "0011011111111100" => data_out <= rom_array(14332);
		when "0011011111111101" => data_out <= rom_array(14333);
		when "0011011111111110" => data_out <= rom_array(14334);
		when "0011011111111111" => data_out <= rom_array(14335);
		when "0011100000000000" => data_out <= rom_array(14336);
		when "0011100000000001" => data_out <= rom_array(14337);
		when "0011100000000010" => data_out <= rom_array(14338);
		when "0011100000000011" => data_out <= rom_array(14339);
		when "0011100000000100" => data_out <= rom_array(14340);
		when "0011100000000101" => data_out <= rom_array(14341);
		when "0011100000000110" => data_out <= rom_array(14342);
		when "0011100000000111" => data_out <= rom_array(14343);
		when "0011100000001000" => data_out <= rom_array(14344);
		when "0011100000001001" => data_out <= rom_array(14345);
		when "0011100000001010" => data_out <= rom_array(14346);
		when "0011100000001011" => data_out <= rom_array(14347);
		when "0011100000001100" => data_out <= rom_array(14348);
		when "0011100000001101" => data_out <= rom_array(14349);
		when "0011100000001110" => data_out <= rom_array(14350);
		when "0011100000001111" => data_out <= rom_array(14351);
		when "0011100000010000" => data_out <= rom_array(14352);
		when "0011100000010001" => data_out <= rom_array(14353);
		when "0011100000010010" => data_out <= rom_array(14354);
		when "0011100000010011" => data_out <= rom_array(14355);
		when "0011100000010100" => data_out <= rom_array(14356);
		when "0011100000010101" => data_out <= rom_array(14357);
		when "0011100000010110" => data_out <= rom_array(14358);
		when "0011100000010111" => data_out <= rom_array(14359);
		when "0011100000011000" => data_out <= rom_array(14360);
		when "0011100000011001" => data_out <= rom_array(14361);
		when "0011100000011010" => data_out <= rom_array(14362);
		when "0011100000011011" => data_out <= rom_array(14363);
		when "0011100000011100" => data_out <= rom_array(14364);
		when "0011100000011101" => data_out <= rom_array(14365);
		when "0011100000011110" => data_out <= rom_array(14366);
		when "0011100000011111" => data_out <= rom_array(14367);
		when "0011100000100000" => data_out <= rom_array(14368);
		when "0011100000100001" => data_out <= rom_array(14369);
		when "0011100000100010" => data_out <= rom_array(14370);
		when "0011100000100011" => data_out <= rom_array(14371);
		when "0011100000100100" => data_out <= rom_array(14372);
		when "0011100000100101" => data_out <= rom_array(14373);
		when "0011100000100110" => data_out <= rom_array(14374);
		when "0011100000100111" => data_out <= rom_array(14375);
		when "0011100000101000" => data_out <= rom_array(14376);
		when "0011100000101001" => data_out <= rom_array(14377);
		when "0011100000101010" => data_out <= rom_array(14378);
		when "0011100000101011" => data_out <= rom_array(14379);
		when "0011100000101100" => data_out <= rom_array(14380);
		when "0011100000101101" => data_out <= rom_array(14381);
		when "0011100000101110" => data_out <= rom_array(14382);
		when "0011100000101111" => data_out <= rom_array(14383);
		when "0011100000110000" => data_out <= rom_array(14384);
		when "0011100000110001" => data_out <= rom_array(14385);
		when "0011100000110010" => data_out <= rom_array(14386);
		when "0011100000110011" => data_out <= rom_array(14387);
		when "0011100000110100" => data_out <= rom_array(14388);
		when "0011100000110101" => data_out <= rom_array(14389);
		when "0011100000110110" => data_out <= rom_array(14390);
		when "0011100000110111" => data_out <= rom_array(14391);
		when "0011100000111000" => data_out <= rom_array(14392);
		when "0011100000111001" => data_out <= rom_array(14393);
		when "0011100000111010" => data_out <= rom_array(14394);
		when "0011100000111011" => data_out <= rom_array(14395);
		when "0011100000111100" => data_out <= rom_array(14396);
		when "0011100000111101" => data_out <= rom_array(14397);
		when "0011100000111110" => data_out <= rom_array(14398);
		when "0011100000111111" => data_out <= rom_array(14399);
		when "0011100001000000" => data_out <= rom_array(14400);
		when "0011100001000001" => data_out <= rom_array(14401);
		when "0011100001000010" => data_out <= rom_array(14402);
		when "0011100001000011" => data_out <= rom_array(14403);
		when "0011100001000100" => data_out <= rom_array(14404);
		when "0011100001000101" => data_out <= rom_array(14405);
		when "0011100001000110" => data_out <= rom_array(14406);
		when "0011100001000111" => data_out <= rom_array(14407);
		when "0011100001001000" => data_out <= rom_array(14408);
		when "0011100001001001" => data_out <= rom_array(14409);
		when "0011100001001010" => data_out <= rom_array(14410);
		when "0011100001001011" => data_out <= rom_array(14411);
		when "0011100001001100" => data_out <= rom_array(14412);
		when "0011100001001101" => data_out <= rom_array(14413);
		when "0011100001001110" => data_out <= rom_array(14414);
		when "0011100001001111" => data_out <= rom_array(14415);
		when "0011100001010000" => data_out <= rom_array(14416);
		when "0011100001010001" => data_out <= rom_array(14417);
		when "0011100001010010" => data_out <= rom_array(14418);
		when "0011100001010011" => data_out <= rom_array(14419);
		when "0011100001010100" => data_out <= rom_array(14420);
		when "0011100001010101" => data_out <= rom_array(14421);
		when "0011100001010110" => data_out <= rom_array(14422);
		when "0011100001010111" => data_out <= rom_array(14423);
		when "0011100001011000" => data_out <= rom_array(14424);
		when "0011100001011001" => data_out <= rom_array(14425);
		when "0011100001011010" => data_out <= rom_array(14426);
		when "0011100001011011" => data_out <= rom_array(14427);
		when "0011100001011100" => data_out <= rom_array(14428);
		when "0011100001011101" => data_out <= rom_array(14429);
		when "0011100001011110" => data_out <= rom_array(14430);
		when "0011100001011111" => data_out <= rom_array(14431);
		when "0011100001100000" => data_out <= rom_array(14432);
		when "0011100001100001" => data_out <= rom_array(14433);
		when "0011100001100010" => data_out <= rom_array(14434);
		when "0011100001100011" => data_out <= rom_array(14435);
		when "0011100001100100" => data_out <= rom_array(14436);
		when "0011100001100101" => data_out <= rom_array(14437);
		when "0011100001100110" => data_out <= rom_array(14438);
		when "0011100001100111" => data_out <= rom_array(14439);
		when "0011100001101000" => data_out <= rom_array(14440);
		when "0011100001101001" => data_out <= rom_array(14441);
		when "0011100001101010" => data_out <= rom_array(14442);
		when "0011100001101011" => data_out <= rom_array(14443);
		when "0011100001101100" => data_out <= rom_array(14444);
		when "0011100001101101" => data_out <= rom_array(14445);
		when "0011100001101110" => data_out <= rom_array(14446);
		when "0011100001101111" => data_out <= rom_array(14447);
		when "0011100001110000" => data_out <= rom_array(14448);
		when "0011100001110001" => data_out <= rom_array(14449);
		when "0011100001110010" => data_out <= rom_array(14450);
		when "0011100001110011" => data_out <= rom_array(14451);
		when "0011100001110100" => data_out <= rom_array(14452);
		when "0011100001110101" => data_out <= rom_array(14453);
		when "0011100001110110" => data_out <= rom_array(14454);
		when "0011100001110111" => data_out <= rom_array(14455);
		when "0011100001111000" => data_out <= rom_array(14456);
		when "0011100001111001" => data_out <= rom_array(14457);
		when "0011100001111010" => data_out <= rom_array(14458);
		when "0011100001111011" => data_out <= rom_array(14459);
		when "0011100001111100" => data_out <= rom_array(14460);
		when "0011100001111101" => data_out <= rom_array(14461);
		when "0011100001111110" => data_out <= rom_array(14462);
		when "0011100001111111" => data_out <= rom_array(14463);
		when "0011100010000000" => data_out <= rom_array(14464);
		when "0011100010000001" => data_out <= rom_array(14465);
		when "0011100010000010" => data_out <= rom_array(14466);
		when "0011100010000011" => data_out <= rom_array(14467);
		when "0011100010000100" => data_out <= rom_array(14468);
		when "0011100010000101" => data_out <= rom_array(14469);
		when "0011100010000110" => data_out <= rom_array(14470);
		when "0011100010000111" => data_out <= rom_array(14471);
		when "0011100010001000" => data_out <= rom_array(14472);
		when "0011100010001001" => data_out <= rom_array(14473);
		when "0011100010001010" => data_out <= rom_array(14474);
		when "0011100010001011" => data_out <= rom_array(14475);
		when "0011100010001100" => data_out <= rom_array(14476);
		when "0011100010001101" => data_out <= rom_array(14477);
		when "0011100010001110" => data_out <= rom_array(14478);
		when "0011100010001111" => data_out <= rom_array(14479);
		when "0011100010010000" => data_out <= rom_array(14480);
		when "0011100010010001" => data_out <= rom_array(14481);
		when "0011100010010010" => data_out <= rom_array(14482);
		when "0011100010010011" => data_out <= rom_array(14483);
		when "0011100010010100" => data_out <= rom_array(14484);
		when "0011100010010101" => data_out <= rom_array(14485);
		when "0011100010010110" => data_out <= rom_array(14486);
		when "0011100010010111" => data_out <= rom_array(14487);
		when "0011100010011000" => data_out <= rom_array(14488);
		when "0011100010011001" => data_out <= rom_array(14489);
		when "0011100010011010" => data_out <= rom_array(14490);
		when "0011100010011011" => data_out <= rom_array(14491);
		when "0011100010011100" => data_out <= rom_array(14492);
		when "0011100010011101" => data_out <= rom_array(14493);
		when "0011100010011110" => data_out <= rom_array(14494);
		when "0011100010011111" => data_out <= rom_array(14495);
		when "0011100010100000" => data_out <= rom_array(14496);
		when "0011100010100001" => data_out <= rom_array(14497);
		when "0011100010100010" => data_out <= rom_array(14498);
		when "0011100010100011" => data_out <= rom_array(14499);
		when "0011100010100100" => data_out <= rom_array(14500);
		when "0011100010100101" => data_out <= rom_array(14501);
		when "0011100010100110" => data_out <= rom_array(14502);
		when "0011100010100111" => data_out <= rom_array(14503);
		when "0011100010101000" => data_out <= rom_array(14504);
		when "0011100010101001" => data_out <= rom_array(14505);
		when "0011100010101010" => data_out <= rom_array(14506);
		when "0011100010101011" => data_out <= rom_array(14507);
		when "0011100010101100" => data_out <= rom_array(14508);
		when "0011100010101101" => data_out <= rom_array(14509);
		when "0011100010101110" => data_out <= rom_array(14510);
		when "0011100010101111" => data_out <= rom_array(14511);
		when "0011100010110000" => data_out <= rom_array(14512);
		when "0011100010110001" => data_out <= rom_array(14513);
		when "0011100010110010" => data_out <= rom_array(14514);
		when "0011100010110011" => data_out <= rom_array(14515);
		when "0011100010110100" => data_out <= rom_array(14516);
		when "0011100010110101" => data_out <= rom_array(14517);
		when "0011100010110110" => data_out <= rom_array(14518);
		when "0011100010110111" => data_out <= rom_array(14519);
		when "0011100010111000" => data_out <= rom_array(14520);
		when "0011100010111001" => data_out <= rom_array(14521);
		when "0011100010111010" => data_out <= rom_array(14522);
		when "0011100010111011" => data_out <= rom_array(14523);
		when "0011100010111100" => data_out <= rom_array(14524);
		when "0011100010111101" => data_out <= rom_array(14525);
		when "0011100010111110" => data_out <= rom_array(14526);
		when "0011100010111111" => data_out <= rom_array(14527);
		when "0011100011000000" => data_out <= rom_array(14528);
		when "0011100011000001" => data_out <= rom_array(14529);
		when "0011100011000010" => data_out <= rom_array(14530);
		when "0011100011000011" => data_out <= rom_array(14531);
		when "0011100011000100" => data_out <= rom_array(14532);
		when "0011100011000101" => data_out <= rom_array(14533);
		when "0011100011000110" => data_out <= rom_array(14534);
		when "0011100011000111" => data_out <= rom_array(14535);
		when "0011100011001000" => data_out <= rom_array(14536);
		when "0011100011001001" => data_out <= rom_array(14537);
		when "0011100011001010" => data_out <= rom_array(14538);
		when "0011100011001011" => data_out <= rom_array(14539);
		when "0011100011001100" => data_out <= rom_array(14540);
		when "0011100011001101" => data_out <= rom_array(14541);
		when "0011100011001110" => data_out <= rom_array(14542);
		when "0011100011001111" => data_out <= rom_array(14543);
		when "0011100011010000" => data_out <= rom_array(14544);
		when "0011100011010001" => data_out <= rom_array(14545);
		when "0011100011010010" => data_out <= rom_array(14546);
		when "0011100011010011" => data_out <= rom_array(14547);
		when "0011100011010100" => data_out <= rom_array(14548);
		when "0011100011010101" => data_out <= rom_array(14549);
		when "0011100011010110" => data_out <= rom_array(14550);
		when "0011100011010111" => data_out <= rom_array(14551);
		when "0011100011011000" => data_out <= rom_array(14552);
		when "0011100011011001" => data_out <= rom_array(14553);
		when "0011100011011010" => data_out <= rom_array(14554);
		when "0011100011011011" => data_out <= rom_array(14555);
		when "0011100011011100" => data_out <= rom_array(14556);
		when "0011100011011101" => data_out <= rom_array(14557);
		when "0011100011011110" => data_out <= rom_array(14558);
		when "0011100011011111" => data_out <= rom_array(14559);
		when "0011100011100000" => data_out <= rom_array(14560);
		when "0011100011100001" => data_out <= rom_array(14561);
		when "0011100011100010" => data_out <= rom_array(14562);
		when "0011100011100011" => data_out <= rom_array(14563);
		when "0011100011100100" => data_out <= rom_array(14564);
		when "0011100011100101" => data_out <= rom_array(14565);
		when "0011100011100110" => data_out <= rom_array(14566);
		when "0011100011100111" => data_out <= rom_array(14567);
		when "0011100011101000" => data_out <= rom_array(14568);
		when "0011100011101001" => data_out <= rom_array(14569);
		when "0011100011101010" => data_out <= rom_array(14570);
		when "0011100011101011" => data_out <= rom_array(14571);
		when "0011100011101100" => data_out <= rom_array(14572);
		when "0011100011101101" => data_out <= rom_array(14573);
		when "0011100011101110" => data_out <= rom_array(14574);
		when "0011100011101111" => data_out <= rom_array(14575);
		when "0011100011110000" => data_out <= rom_array(14576);
		when "0011100011110001" => data_out <= rom_array(14577);
		when "0011100011110010" => data_out <= rom_array(14578);
		when "0011100011110011" => data_out <= rom_array(14579);
		when "0011100011110100" => data_out <= rom_array(14580);
		when "0011100011110101" => data_out <= rom_array(14581);
		when "0011100011110110" => data_out <= rom_array(14582);
		when "0011100011110111" => data_out <= rom_array(14583);
		when "0011100011111000" => data_out <= rom_array(14584);
		when "0011100011111001" => data_out <= rom_array(14585);
		when "0011100011111010" => data_out <= rom_array(14586);
		when "0011100011111011" => data_out <= rom_array(14587);
		when "0011100011111100" => data_out <= rom_array(14588);
		when "0011100011111101" => data_out <= rom_array(14589);
		when "0011100011111110" => data_out <= rom_array(14590);
		when "0011100011111111" => data_out <= rom_array(14591);
		when "0011100100000000" => data_out <= rom_array(14592);
		when "0011100100000001" => data_out <= rom_array(14593);
		when "0011100100000010" => data_out <= rom_array(14594);
		when "0011100100000011" => data_out <= rom_array(14595);
		when "0011100100000100" => data_out <= rom_array(14596);
		when "0011100100000101" => data_out <= rom_array(14597);
		when "0011100100000110" => data_out <= rom_array(14598);
		when "0011100100000111" => data_out <= rom_array(14599);
		when "0011100100001000" => data_out <= rom_array(14600);
		when "0011100100001001" => data_out <= rom_array(14601);
		when "0011100100001010" => data_out <= rom_array(14602);
		when "0011100100001011" => data_out <= rom_array(14603);
		when "0011100100001100" => data_out <= rom_array(14604);
		when "0011100100001101" => data_out <= rom_array(14605);
		when "0011100100001110" => data_out <= rom_array(14606);
		when "0011100100001111" => data_out <= rom_array(14607);
		when "0011100100010000" => data_out <= rom_array(14608);
		when "0011100100010001" => data_out <= rom_array(14609);
		when "0011100100010010" => data_out <= rom_array(14610);
		when "0011100100010011" => data_out <= rom_array(14611);
		when "0011100100010100" => data_out <= rom_array(14612);
		when "0011100100010101" => data_out <= rom_array(14613);
		when "0011100100010110" => data_out <= rom_array(14614);
		when "0011100100010111" => data_out <= rom_array(14615);
		when "0011100100011000" => data_out <= rom_array(14616);
		when "0011100100011001" => data_out <= rom_array(14617);
		when "0011100100011010" => data_out <= rom_array(14618);
		when "0011100100011011" => data_out <= rom_array(14619);
		when "0011100100011100" => data_out <= rom_array(14620);
		when "0011100100011101" => data_out <= rom_array(14621);
		when "0011100100011110" => data_out <= rom_array(14622);
		when "0011100100011111" => data_out <= rom_array(14623);
		when "0011100100100000" => data_out <= rom_array(14624);
		when "0011100100100001" => data_out <= rom_array(14625);
		when "0011100100100010" => data_out <= rom_array(14626);
		when "0011100100100011" => data_out <= rom_array(14627);
		when "0011100100100100" => data_out <= rom_array(14628);
		when "0011100100100101" => data_out <= rom_array(14629);
		when "0011100100100110" => data_out <= rom_array(14630);
		when "0011100100100111" => data_out <= rom_array(14631);
		when "0011100100101000" => data_out <= rom_array(14632);
		when "0011100100101001" => data_out <= rom_array(14633);
		when "0011100100101010" => data_out <= rom_array(14634);
		when "0011100100101011" => data_out <= rom_array(14635);
		when "0011100100101100" => data_out <= rom_array(14636);
		when "0011100100101101" => data_out <= rom_array(14637);
		when "0011100100101110" => data_out <= rom_array(14638);
		when "0011100100101111" => data_out <= rom_array(14639);
		when "0011100100110000" => data_out <= rom_array(14640);
		when "0011100100110001" => data_out <= rom_array(14641);
		when "0011100100110010" => data_out <= rom_array(14642);
		when "0011100100110011" => data_out <= rom_array(14643);
		when "0011100100110100" => data_out <= rom_array(14644);
		when "0011100100110101" => data_out <= rom_array(14645);
		when "0011100100110110" => data_out <= rom_array(14646);
		when "0011100100110111" => data_out <= rom_array(14647);
		when "0011100100111000" => data_out <= rom_array(14648);
		when "0011100100111001" => data_out <= rom_array(14649);
		when "0011100100111010" => data_out <= rom_array(14650);
		when "0011100100111011" => data_out <= rom_array(14651);
		when "0011100100111100" => data_out <= rom_array(14652);
		when "0011100100111101" => data_out <= rom_array(14653);
		when "0011100100111110" => data_out <= rom_array(14654);
		when "0011100100111111" => data_out <= rom_array(14655);
		when "0011100101000000" => data_out <= rom_array(14656);
		when "0011100101000001" => data_out <= rom_array(14657);
		when "0011100101000010" => data_out <= rom_array(14658);
		when "0011100101000011" => data_out <= rom_array(14659);
		when "0011100101000100" => data_out <= rom_array(14660);
		when "0011100101000101" => data_out <= rom_array(14661);
		when "0011100101000110" => data_out <= rom_array(14662);
		when "0011100101000111" => data_out <= rom_array(14663);
		when "0011100101001000" => data_out <= rom_array(14664);
		when "0011100101001001" => data_out <= rom_array(14665);
		when "0011100101001010" => data_out <= rom_array(14666);
		when "0011100101001011" => data_out <= rom_array(14667);
		when "0011100101001100" => data_out <= rom_array(14668);
		when "0011100101001101" => data_out <= rom_array(14669);
		when "0011100101001110" => data_out <= rom_array(14670);
		when "0011100101001111" => data_out <= rom_array(14671);
		when "0011100101010000" => data_out <= rom_array(14672);
		when "0011100101010001" => data_out <= rom_array(14673);
		when "0011100101010010" => data_out <= rom_array(14674);
		when "0011100101010011" => data_out <= rom_array(14675);
		when "0011100101010100" => data_out <= rom_array(14676);
		when "0011100101010101" => data_out <= rom_array(14677);
		when "0011100101010110" => data_out <= rom_array(14678);
		when "0011100101010111" => data_out <= rom_array(14679);
		when "0011100101011000" => data_out <= rom_array(14680);
		when "0011100101011001" => data_out <= rom_array(14681);
		when "0011100101011010" => data_out <= rom_array(14682);
		when "0011100101011011" => data_out <= rom_array(14683);
		when "0011100101011100" => data_out <= rom_array(14684);
		when "0011100101011101" => data_out <= rom_array(14685);
		when "0011100101011110" => data_out <= rom_array(14686);
		when "0011100101011111" => data_out <= rom_array(14687);
		when "0011100101100000" => data_out <= rom_array(14688);
		when "0011100101100001" => data_out <= rom_array(14689);
		when "0011100101100010" => data_out <= rom_array(14690);
		when "0011100101100011" => data_out <= rom_array(14691);
		when "0011100101100100" => data_out <= rom_array(14692);
		when "0011100101100101" => data_out <= rom_array(14693);
		when "0011100101100110" => data_out <= rom_array(14694);
		when "0011100101100111" => data_out <= rom_array(14695);
		when "0011100101101000" => data_out <= rom_array(14696);
		when "0011100101101001" => data_out <= rom_array(14697);
		when "0011100101101010" => data_out <= rom_array(14698);
		when "0011100101101011" => data_out <= rom_array(14699);
		when "0011100101101100" => data_out <= rom_array(14700);
		when "0011100101101101" => data_out <= rom_array(14701);
		when "0011100101101110" => data_out <= rom_array(14702);
		when "0011100101101111" => data_out <= rom_array(14703);
		when "0011100101110000" => data_out <= rom_array(14704);
		when "0011100101110001" => data_out <= rom_array(14705);
		when "0011100101110010" => data_out <= rom_array(14706);
		when "0011100101110011" => data_out <= rom_array(14707);
		when "0011100101110100" => data_out <= rom_array(14708);
		when "0011100101110101" => data_out <= rom_array(14709);
		when "0011100101110110" => data_out <= rom_array(14710);
		when "0011100101110111" => data_out <= rom_array(14711);
		when "0011100101111000" => data_out <= rom_array(14712);
		when "0011100101111001" => data_out <= rom_array(14713);
		when "0011100101111010" => data_out <= rom_array(14714);
		when "0011100101111011" => data_out <= rom_array(14715);
		when "0011100101111100" => data_out <= rom_array(14716);
		when "0011100101111101" => data_out <= rom_array(14717);
		when "0011100101111110" => data_out <= rom_array(14718);
		when "0011100101111111" => data_out <= rom_array(14719);
		when "0011100110000000" => data_out <= rom_array(14720);
		when "0011100110000001" => data_out <= rom_array(14721);
		when "0011100110000010" => data_out <= rom_array(14722);
		when "0011100110000011" => data_out <= rom_array(14723);
		when "0011100110000100" => data_out <= rom_array(14724);
		when "0011100110000101" => data_out <= rom_array(14725);
		when "0011100110000110" => data_out <= rom_array(14726);
		when "0011100110000111" => data_out <= rom_array(14727);
		when "0011100110001000" => data_out <= rom_array(14728);
		when "0011100110001001" => data_out <= rom_array(14729);
		when "0011100110001010" => data_out <= rom_array(14730);
		when "0011100110001011" => data_out <= rom_array(14731);
		when "0011100110001100" => data_out <= rom_array(14732);
		when "0011100110001101" => data_out <= rom_array(14733);
		when "0011100110001110" => data_out <= rom_array(14734);
		when "0011100110001111" => data_out <= rom_array(14735);
		when "0011100110010000" => data_out <= rom_array(14736);
		when "0011100110010001" => data_out <= rom_array(14737);
		when "0011100110010010" => data_out <= rom_array(14738);
		when "0011100110010011" => data_out <= rom_array(14739);
		when "0011100110010100" => data_out <= rom_array(14740);
		when "0011100110010101" => data_out <= rom_array(14741);
		when "0011100110010110" => data_out <= rom_array(14742);
		when "0011100110010111" => data_out <= rom_array(14743);
		when "0011100110011000" => data_out <= rom_array(14744);
		when "0011100110011001" => data_out <= rom_array(14745);
		when "0011100110011010" => data_out <= rom_array(14746);
		when "0011100110011011" => data_out <= rom_array(14747);
		when "0011100110011100" => data_out <= rom_array(14748);
		when "0011100110011101" => data_out <= rom_array(14749);
		when "0011100110011110" => data_out <= rom_array(14750);
		when "0011100110011111" => data_out <= rom_array(14751);
		when "0011100110100000" => data_out <= rom_array(14752);
		when "0011100110100001" => data_out <= rom_array(14753);
		when "0011100110100010" => data_out <= rom_array(14754);
		when "0011100110100011" => data_out <= rom_array(14755);
		when "0011100110100100" => data_out <= rom_array(14756);
		when "0011100110100101" => data_out <= rom_array(14757);
		when "0011100110100110" => data_out <= rom_array(14758);
		when "0011100110100111" => data_out <= rom_array(14759);
		when "0011100110101000" => data_out <= rom_array(14760);
		when "0011100110101001" => data_out <= rom_array(14761);
		when "0011100110101010" => data_out <= rom_array(14762);
		when "0011100110101011" => data_out <= rom_array(14763);
		when "0011100110101100" => data_out <= rom_array(14764);
		when "0011100110101101" => data_out <= rom_array(14765);
		when "0011100110101110" => data_out <= rom_array(14766);
		when "0011100110101111" => data_out <= rom_array(14767);
		when "0011100110110000" => data_out <= rom_array(14768);
		when "0011100110110001" => data_out <= rom_array(14769);
		when "0011100110110010" => data_out <= rom_array(14770);
		when "0011100110110011" => data_out <= rom_array(14771);
		when "0011100110110100" => data_out <= rom_array(14772);
		when "0011100110110101" => data_out <= rom_array(14773);
		when "0011100110110110" => data_out <= rom_array(14774);
		when "0011100110110111" => data_out <= rom_array(14775);
		when "0011100110111000" => data_out <= rom_array(14776);
		when "0011100110111001" => data_out <= rom_array(14777);
		when "0011100110111010" => data_out <= rom_array(14778);
		when "0011100110111011" => data_out <= rom_array(14779);
		when "0011100110111100" => data_out <= rom_array(14780);
		when "0011100110111101" => data_out <= rom_array(14781);
		when "0011100110111110" => data_out <= rom_array(14782);
		when "0011100110111111" => data_out <= rom_array(14783);
		when "0011100111000000" => data_out <= rom_array(14784);
		when "0011100111000001" => data_out <= rom_array(14785);
		when "0011100111000010" => data_out <= rom_array(14786);
		when "0011100111000011" => data_out <= rom_array(14787);
		when "0011100111000100" => data_out <= rom_array(14788);
		when "0011100111000101" => data_out <= rom_array(14789);
		when "0011100111000110" => data_out <= rom_array(14790);
		when "0011100111000111" => data_out <= rom_array(14791);
		when "0011100111001000" => data_out <= rom_array(14792);
		when "0011100111001001" => data_out <= rom_array(14793);
		when "0011100111001010" => data_out <= rom_array(14794);
		when "0011100111001011" => data_out <= rom_array(14795);
		when "0011100111001100" => data_out <= rom_array(14796);
		when "0011100111001101" => data_out <= rom_array(14797);
		when "0011100111001110" => data_out <= rom_array(14798);
		when "0011100111001111" => data_out <= rom_array(14799);
		when "0011100111010000" => data_out <= rom_array(14800);
		when "0011100111010001" => data_out <= rom_array(14801);
		when "0011100111010010" => data_out <= rom_array(14802);
		when "0011100111010011" => data_out <= rom_array(14803);
		when "0011100111010100" => data_out <= rom_array(14804);
		when "0011100111010101" => data_out <= rom_array(14805);
		when "0011100111010110" => data_out <= rom_array(14806);
		when "0011100111010111" => data_out <= rom_array(14807);
		when "0011100111011000" => data_out <= rom_array(14808);
		when "0011100111011001" => data_out <= rom_array(14809);
		when "0011100111011010" => data_out <= rom_array(14810);
		when "0011100111011011" => data_out <= rom_array(14811);
		when "0011100111011100" => data_out <= rom_array(14812);
		when "0011100111011101" => data_out <= rom_array(14813);
		when "0011100111011110" => data_out <= rom_array(14814);
		when "0011100111011111" => data_out <= rom_array(14815);
		when "0011100111100000" => data_out <= rom_array(14816);
		when "0011100111100001" => data_out <= rom_array(14817);
		when "0011100111100010" => data_out <= rom_array(14818);
		when "0011100111100011" => data_out <= rom_array(14819);
		when "0011100111100100" => data_out <= rom_array(14820);
		when "0011100111100101" => data_out <= rom_array(14821);
		when "0011100111100110" => data_out <= rom_array(14822);
		when "0011100111100111" => data_out <= rom_array(14823);
		when "0011100111101000" => data_out <= rom_array(14824);
		when "0011100111101001" => data_out <= rom_array(14825);
		when "0011100111101010" => data_out <= rom_array(14826);
		when "0011100111101011" => data_out <= rom_array(14827);
		when "0011100111101100" => data_out <= rom_array(14828);
		when "0011100111101101" => data_out <= rom_array(14829);
		when "0011100111101110" => data_out <= rom_array(14830);
		when "0011100111101111" => data_out <= rom_array(14831);
		when "0011100111110000" => data_out <= rom_array(14832);
		when "0011100111110001" => data_out <= rom_array(14833);
		when "0011100111110010" => data_out <= rom_array(14834);
		when "0011100111110011" => data_out <= rom_array(14835);
		when "0011100111110100" => data_out <= rom_array(14836);
		when "0011100111110101" => data_out <= rom_array(14837);
		when "0011100111110110" => data_out <= rom_array(14838);
		when "0011100111110111" => data_out <= rom_array(14839);
		when "0011100111111000" => data_out <= rom_array(14840);
		when "0011100111111001" => data_out <= rom_array(14841);
		when "0011100111111010" => data_out <= rom_array(14842);
		when "0011100111111011" => data_out <= rom_array(14843);
		when "0011100111111100" => data_out <= rom_array(14844);
		when "0011100111111101" => data_out <= rom_array(14845);
		when "0011100111111110" => data_out <= rom_array(14846);
		when "0011100111111111" => data_out <= rom_array(14847);
		when "0011101000000000" => data_out <= rom_array(14848);
		when "0011101000000001" => data_out <= rom_array(14849);
		when "0011101000000010" => data_out <= rom_array(14850);
		when "0011101000000011" => data_out <= rom_array(14851);
		when "0011101000000100" => data_out <= rom_array(14852);
		when "0011101000000101" => data_out <= rom_array(14853);
		when "0011101000000110" => data_out <= rom_array(14854);
		when "0011101000000111" => data_out <= rom_array(14855);
		when "0011101000001000" => data_out <= rom_array(14856);
		when "0011101000001001" => data_out <= rom_array(14857);
		when "0011101000001010" => data_out <= rom_array(14858);
		when "0011101000001011" => data_out <= rom_array(14859);
		when "0011101000001100" => data_out <= rom_array(14860);
		when "0011101000001101" => data_out <= rom_array(14861);
		when "0011101000001110" => data_out <= rom_array(14862);
		when "0011101000001111" => data_out <= rom_array(14863);
		when "0011101000010000" => data_out <= rom_array(14864);
		when "0011101000010001" => data_out <= rom_array(14865);
		when "0011101000010010" => data_out <= rom_array(14866);
		when "0011101000010011" => data_out <= rom_array(14867);
		when "0011101000010100" => data_out <= rom_array(14868);
		when "0011101000010101" => data_out <= rom_array(14869);
		when "0011101000010110" => data_out <= rom_array(14870);
		when "0011101000010111" => data_out <= rom_array(14871);
		when "0011101000011000" => data_out <= rom_array(14872);
		when "0011101000011001" => data_out <= rom_array(14873);
		when "0011101000011010" => data_out <= rom_array(14874);
		when "0011101000011011" => data_out <= rom_array(14875);
		when "0011101000011100" => data_out <= rom_array(14876);
		when "0011101000011101" => data_out <= rom_array(14877);
		when "0011101000011110" => data_out <= rom_array(14878);
		when "0011101000011111" => data_out <= rom_array(14879);
		when "0011101000100000" => data_out <= rom_array(14880);
		when "0011101000100001" => data_out <= rom_array(14881);
		when "0011101000100010" => data_out <= rom_array(14882);
		when "0011101000100011" => data_out <= rom_array(14883);
		when "0011101000100100" => data_out <= rom_array(14884);
		when "0011101000100101" => data_out <= rom_array(14885);
		when "0011101000100110" => data_out <= rom_array(14886);
		when "0011101000100111" => data_out <= rom_array(14887);
		when "0011101000101000" => data_out <= rom_array(14888);
		when "0011101000101001" => data_out <= rom_array(14889);
		when "0011101000101010" => data_out <= rom_array(14890);
		when "0011101000101011" => data_out <= rom_array(14891);
		when "0011101000101100" => data_out <= rom_array(14892);
		when "0011101000101101" => data_out <= rom_array(14893);
		when "0011101000101110" => data_out <= rom_array(14894);
		when "0011101000101111" => data_out <= rom_array(14895);
		when "0011101000110000" => data_out <= rom_array(14896);
		when "0011101000110001" => data_out <= rom_array(14897);
		when "0011101000110010" => data_out <= rom_array(14898);
		when "0011101000110011" => data_out <= rom_array(14899);
		when "0011101000110100" => data_out <= rom_array(14900);
		when "0011101000110101" => data_out <= rom_array(14901);
		when "0011101000110110" => data_out <= rom_array(14902);
		when "0011101000110111" => data_out <= rom_array(14903);
		when "0011101000111000" => data_out <= rom_array(14904);
		when "0011101000111001" => data_out <= rom_array(14905);
		when "0011101000111010" => data_out <= rom_array(14906);
		when "0011101000111011" => data_out <= rom_array(14907);
		when "0011101000111100" => data_out <= rom_array(14908);
		when "0011101000111101" => data_out <= rom_array(14909);
		when "0011101000111110" => data_out <= rom_array(14910);
		when "0011101000111111" => data_out <= rom_array(14911);
		when "0011101001000000" => data_out <= rom_array(14912);
		when "0011101001000001" => data_out <= rom_array(14913);
		when "0011101001000010" => data_out <= rom_array(14914);
		when "0011101001000011" => data_out <= rom_array(14915);
		when "0011101001000100" => data_out <= rom_array(14916);
		when "0011101001000101" => data_out <= rom_array(14917);
		when "0011101001000110" => data_out <= rom_array(14918);
		when "0011101001000111" => data_out <= rom_array(14919);
		when "0011101001001000" => data_out <= rom_array(14920);
		when "0011101001001001" => data_out <= rom_array(14921);
		when "0011101001001010" => data_out <= rom_array(14922);
		when "0011101001001011" => data_out <= rom_array(14923);
		when "0011101001001100" => data_out <= rom_array(14924);
		when "0011101001001101" => data_out <= rom_array(14925);
		when "0011101001001110" => data_out <= rom_array(14926);
		when "0011101001001111" => data_out <= rom_array(14927);
		when "0011101001010000" => data_out <= rom_array(14928);
		when "0011101001010001" => data_out <= rom_array(14929);
		when "0011101001010010" => data_out <= rom_array(14930);
		when "0011101001010011" => data_out <= rom_array(14931);
		when "0011101001010100" => data_out <= rom_array(14932);
		when "0011101001010101" => data_out <= rom_array(14933);
		when "0011101001010110" => data_out <= rom_array(14934);
		when "0011101001010111" => data_out <= rom_array(14935);
		when "0011101001011000" => data_out <= rom_array(14936);
		when "0011101001011001" => data_out <= rom_array(14937);
		when "0011101001011010" => data_out <= rom_array(14938);
		when "0011101001011011" => data_out <= rom_array(14939);
		when "0011101001011100" => data_out <= rom_array(14940);
		when "0011101001011101" => data_out <= rom_array(14941);
		when "0011101001011110" => data_out <= rom_array(14942);
		when "0011101001011111" => data_out <= rom_array(14943);
		when "0011101001100000" => data_out <= rom_array(14944);
		when "0011101001100001" => data_out <= rom_array(14945);
		when "0011101001100010" => data_out <= rom_array(14946);
		when "0011101001100011" => data_out <= rom_array(14947);
		when "0011101001100100" => data_out <= rom_array(14948);
		when "0011101001100101" => data_out <= rom_array(14949);
		when "0011101001100110" => data_out <= rom_array(14950);
		when "0011101001100111" => data_out <= rom_array(14951);
		when "0011101001101000" => data_out <= rom_array(14952);
		when "0011101001101001" => data_out <= rom_array(14953);
		when "0011101001101010" => data_out <= rom_array(14954);
		when "0011101001101011" => data_out <= rom_array(14955);
		when "0011101001101100" => data_out <= rom_array(14956);
		when "0011101001101101" => data_out <= rom_array(14957);
		when "0011101001101110" => data_out <= rom_array(14958);
		when "0011101001101111" => data_out <= rom_array(14959);
		when "0011101001110000" => data_out <= rom_array(14960);
		when "0011101001110001" => data_out <= rom_array(14961);
		when "0011101001110010" => data_out <= rom_array(14962);
		when "0011101001110011" => data_out <= rom_array(14963);
		when "0011101001110100" => data_out <= rom_array(14964);
		when "0011101001110101" => data_out <= rom_array(14965);
		when "0011101001110110" => data_out <= rom_array(14966);
		when "0011101001110111" => data_out <= rom_array(14967);
		when "0011101001111000" => data_out <= rom_array(14968);
		when "0011101001111001" => data_out <= rom_array(14969);
		when "0011101001111010" => data_out <= rom_array(14970);
		when "0011101001111011" => data_out <= rom_array(14971);
		when "0011101001111100" => data_out <= rom_array(14972);
		when "0011101001111101" => data_out <= rom_array(14973);
		when "0011101001111110" => data_out <= rom_array(14974);
		when "0011101001111111" => data_out <= rom_array(14975);
		when "0011101010000000" => data_out <= rom_array(14976);
		when "0011101010000001" => data_out <= rom_array(14977);
		when "0011101010000010" => data_out <= rom_array(14978);
		when "0011101010000011" => data_out <= rom_array(14979);
		when "0011101010000100" => data_out <= rom_array(14980);
		when "0011101010000101" => data_out <= rom_array(14981);
		when "0011101010000110" => data_out <= rom_array(14982);
		when "0011101010000111" => data_out <= rom_array(14983);
		when "0011101010001000" => data_out <= rom_array(14984);
		when "0011101010001001" => data_out <= rom_array(14985);
		when "0011101010001010" => data_out <= rom_array(14986);
		when "0011101010001011" => data_out <= rom_array(14987);
		when "0011101010001100" => data_out <= rom_array(14988);
		when "0011101010001101" => data_out <= rom_array(14989);
		when "0011101010001110" => data_out <= rom_array(14990);
		when "0011101010001111" => data_out <= rom_array(14991);
		when "0011101010010000" => data_out <= rom_array(14992);
		when "0011101010010001" => data_out <= rom_array(14993);
		when "0011101010010010" => data_out <= rom_array(14994);
		when "0011101010010011" => data_out <= rom_array(14995);
		when "0011101010010100" => data_out <= rom_array(14996);
		when "0011101010010101" => data_out <= rom_array(14997);
		when "0011101010010110" => data_out <= rom_array(14998);
		when "0011101010010111" => data_out <= rom_array(14999);
		when "0011101010011000" => data_out <= rom_array(15000);
		when "0011101010011001" => data_out <= rom_array(15001);
		when "0011101010011010" => data_out <= rom_array(15002);
		when "0011101010011011" => data_out <= rom_array(15003);
		when "0011101010011100" => data_out <= rom_array(15004);
		when "0011101010011101" => data_out <= rom_array(15005);
		when "0011101010011110" => data_out <= rom_array(15006);
		when "0011101010011111" => data_out <= rom_array(15007);
		when "0011101010100000" => data_out <= rom_array(15008);
		when "0011101010100001" => data_out <= rom_array(15009);
		when "0011101010100010" => data_out <= rom_array(15010);
		when "0011101010100011" => data_out <= rom_array(15011);
		when "0011101010100100" => data_out <= rom_array(15012);
		when "0011101010100101" => data_out <= rom_array(15013);
		when "0011101010100110" => data_out <= rom_array(15014);
		when "0011101010100111" => data_out <= rom_array(15015);
		when "0011101010101000" => data_out <= rom_array(15016);
		when "0011101010101001" => data_out <= rom_array(15017);
		when "0011101010101010" => data_out <= rom_array(15018);
		when "0011101010101011" => data_out <= rom_array(15019);
		when "0011101010101100" => data_out <= rom_array(15020);
		when "0011101010101101" => data_out <= rom_array(15021);
		when "0011101010101110" => data_out <= rom_array(15022);
		when "0011101010101111" => data_out <= rom_array(15023);
		when "0011101010110000" => data_out <= rom_array(15024);
		when "0011101010110001" => data_out <= rom_array(15025);
		when "0011101010110010" => data_out <= rom_array(15026);
		when "0011101010110011" => data_out <= rom_array(15027);
		when "0011101010110100" => data_out <= rom_array(15028);
		when "0011101010110101" => data_out <= rom_array(15029);
		when "0011101010110110" => data_out <= rom_array(15030);
		when "0011101010110111" => data_out <= rom_array(15031);
		when "0011101010111000" => data_out <= rom_array(15032);
		when "0011101010111001" => data_out <= rom_array(15033);
		when "0011101010111010" => data_out <= rom_array(15034);
		when "0011101010111011" => data_out <= rom_array(15035);
		when "0011101010111100" => data_out <= rom_array(15036);
		when "0011101010111101" => data_out <= rom_array(15037);
		when "0011101010111110" => data_out <= rom_array(15038);
		when "0011101010111111" => data_out <= rom_array(15039);
		when "0011101011000000" => data_out <= rom_array(15040);
		when "0011101011000001" => data_out <= rom_array(15041);
		when "0011101011000010" => data_out <= rom_array(15042);
		when "0011101011000011" => data_out <= rom_array(15043);
		when "0011101011000100" => data_out <= rom_array(15044);
		when "0011101011000101" => data_out <= rom_array(15045);
		when "0011101011000110" => data_out <= rom_array(15046);
		when "0011101011000111" => data_out <= rom_array(15047);
		when "0011101011001000" => data_out <= rom_array(15048);
		when "0011101011001001" => data_out <= rom_array(15049);
		when "0011101011001010" => data_out <= rom_array(15050);
		when "0011101011001011" => data_out <= rom_array(15051);
		when "0011101011001100" => data_out <= rom_array(15052);
		when "0011101011001101" => data_out <= rom_array(15053);
		when "0011101011001110" => data_out <= rom_array(15054);
		when "0011101011001111" => data_out <= rom_array(15055);
		when "0011101011010000" => data_out <= rom_array(15056);
		when "0011101011010001" => data_out <= rom_array(15057);
		when "0011101011010010" => data_out <= rom_array(15058);
		when "0011101011010011" => data_out <= rom_array(15059);
		when "0011101011010100" => data_out <= rom_array(15060);
		when "0011101011010101" => data_out <= rom_array(15061);
		when "0011101011010110" => data_out <= rom_array(15062);
		when "0011101011010111" => data_out <= rom_array(15063);
		when "0011101011011000" => data_out <= rom_array(15064);
		when "0011101011011001" => data_out <= rom_array(15065);
		when "0011101011011010" => data_out <= rom_array(15066);
		when "0011101011011011" => data_out <= rom_array(15067);
		when "0011101011011100" => data_out <= rom_array(15068);
		when "0011101011011101" => data_out <= rom_array(15069);
		when "0011101011011110" => data_out <= rom_array(15070);
		when "0011101011011111" => data_out <= rom_array(15071);
		when "0011101011100000" => data_out <= rom_array(15072);
		when "0011101011100001" => data_out <= rom_array(15073);
		when "0011101011100010" => data_out <= rom_array(15074);
		when "0011101011100011" => data_out <= rom_array(15075);
		when "0011101011100100" => data_out <= rom_array(15076);
		when "0011101011100101" => data_out <= rom_array(15077);
		when "0011101011100110" => data_out <= rom_array(15078);
		when "0011101011100111" => data_out <= rom_array(15079);
		when "0011101011101000" => data_out <= rom_array(15080);
		when "0011101011101001" => data_out <= rom_array(15081);
		when "0011101011101010" => data_out <= rom_array(15082);
		when "0011101011101011" => data_out <= rom_array(15083);
		when "0011101011101100" => data_out <= rom_array(15084);
		when "0011101011101101" => data_out <= rom_array(15085);
		when "0011101011101110" => data_out <= rom_array(15086);
		when "0011101011101111" => data_out <= rom_array(15087);
		when "0011101011110000" => data_out <= rom_array(15088);
		when "0011101011110001" => data_out <= rom_array(15089);
		when "0011101011110010" => data_out <= rom_array(15090);
		when "0011101011110011" => data_out <= rom_array(15091);
		when "0011101011110100" => data_out <= rom_array(15092);
		when "0011101011110101" => data_out <= rom_array(15093);
		when "0011101011110110" => data_out <= rom_array(15094);
		when "0011101011110111" => data_out <= rom_array(15095);
		when "0011101011111000" => data_out <= rom_array(15096);
		when "0011101011111001" => data_out <= rom_array(15097);
		when "0011101011111010" => data_out <= rom_array(15098);
		when "0011101011111011" => data_out <= rom_array(15099);
		when "0011101011111100" => data_out <= rom_array(15100);
		when "0011101011111101" => data_out <= rom_array(15101);
		when "0011101011111110" => data_out <= rom_array(15102);
		when "0011101011111111" => data_out <= rom_array(15103);
		when "0011101100000000" => data_out <= rom_array(15104);
		when "0011101100000001" => data_out <= rom_array(15105);
		when "0011101100000010" => data_out <= rom_array(15106);
		when "0011101100000011" => data_out <= rom_array(15107);
		when "0011101100000100" => data_out <= rom_array(15108);
		when "0011101100000101" => data_out <= rom_array(15109);
		when "0011101100000110" => data_out <= rom_array(15110);
		when "0011101100000111" => data_out <= rom_array(15111);
		when "0011101100001000" => data_out <= rom_array(15112);
		when "0011101100001001" => data_out <= rom_array(15113);
		when "0011101100001010" => data_out <= rom_array(15114);
		when "0011101100001011" => data_out <= rom_array(15115);
		when "0011101100001100" => data_out <= rom_array(15116);
		when "0011101100001101" => data_out <= rom_array(15117);
		when "0011101100001110" => data_out <= rom_array(15118);
		when "0011101100001111" => data_out <= rom_array(15119);
		when "0011101100010000" => data_out <= rom_array(15120);
		when "0011101100010001" => data_out <= rom_array(15121);
		when "0011101100010010" => data_out <= rom_array(15122);
		when "0011101100010011" => data_out <= rom_array(15123);
		when "0011101100010100" => data_out <= rom_array(15124);
		when "0011101100010101" => data_out <= rom_array(15125);
		when "0011101100010110" => data_out <= rom_array(15126);
		when "0011101100010111" => data_out <= rom_array(15127);
		when "0011101100011000" => data_out <= rom_array(15128);
		when "0011101100011001" => data_out <= rom_array(15129);
		when "0011101100011010" => data_out <= rom_array(15130);
		when "0011101100011011" => data_out <= rom_array(15131);
		when "0011101100011100" => data_out <= rom_array(15132);
		when "0011101100011101" => data_out <= rom_array(15133);
		when "0011101100011110" => data_out <= rom_array(15134);
		when "0011101100011111" => data_out <= rom_array(15135);
		when "0011101100100000" => data_out <= rom_array(15136);
		when "0011101100100001" => data_out <= rom_array(15137);
		when "0011101100100010" => data_out <= rom_array(15138);
		when "0011101100100011" => data_out <= rom_array(15139);
		when "0011101100100100" => data_out <= rom_array(15140);
		when "0011101100100101" => data_out <= rom_array(15141);
		when "0011101100100110" => data_out <= rom_array(15142);
		when "0011101100100111" => data_out <= rom_array(15143);
		when "0011101100101000" => data_out <= rom_array(15144);
		when "0011101100101001" => data_out <= rom_array(15145);
		when "0011101100101010" => data_out <= rom_array(15146);
		when "0011101100101011" => data_out <= rom_array(15147);
		when "0011101100101100" => data_out <= rom_array(15148);
		when "0011101100101101" => data_out <= rom_array(15149);
		when "0011101100101110" => data_out <= rom_array(15150);
		when "0011101100101111" => data_out <= rom_array(15151);
		when "0011101100110000" => data_out <= rom_array(15152);
		when "0011101100110001" => data_out <= rom_array(15153);
		when "0011101100110010" => data_out <= rom_array(15154);
		when "0011101100110011" => data_out <= rom_array(15155);
		when "0011101100110100" => data_out <= rom_array(15156);
		when "0011101100110101" => data_out <= rom_array(15157);
		when "0011101100110110" => data_out <= rom_array(15158);
		when "0011101100110111" => data_out <= rom_array(15159);
		when "0011101100111000" => data_out <= rom_array(15160);
		when "0011101100111001" => data_out <= rom_array(15161);
		when "0011101100111010" => data_out <= rom_array(15162);
		when "0011101100111011" => data_out <= rom_array(15163);
		when "0011101100111100" => data_out <= rom_array(15164);
		when "0011101100111101" => data_out <= rom_array(15165);
		when "0011101100111110" => data_out <= rom_array(15166);
		when "0011101100111111" => data_out <= rom_array(15167);
		when "0011101101000000" => data_out <= rom_array(15168);
		when "0011101101000001" => data_out <= rom_array(15169);
		when "0011101101000010" => data_out <= rom_array(15170);
		when "0011101101000011" => data_out <= rom_array(15171);
		when "0011101101000100" => data_out <= rom_array(15172);
		when "0011101101000101" => data_out <= rom_array(15173);
		when "0011101101000110" => data_out <= rom_array(15174);
		when "0011101101000111" => data_out <= rom_array(15175);
		when "0011101101001000" => data_out <= rom_array(15176);
		when "0011101101001001" => data_out <= rom_array(15177);
		when "0011101101001010" => data_out <= rom_array(15178);
		when "0011101101001011" => data_out <= rom_array(15179);
		when "0011101101001100" => data_out <= rom_array(15180);
		when "0011101101001101" => data_out <= rom_array(15181);
		when "0011101101001110" => data_out <= rom_array(15182);
		when "0011101101001111" => data_out <= rom_array(15183);
		when "0011101101010000" => data_out <= rom_array(15184);
		when "0011101101010001" => data_out <= rom_array(15185);
		when "0011101101010010" => data_out <= rom_array(15186);
		when "0011101101010011" => data_out <= rom_array(15187);
		when "0011101101010100" => data_out <= rom_array(15188);
		when "0011101101010101" => data_out <= rom_array(15189);
		when "0011101101010110" => data_out <= rom_array(15190);
		when "0011101101010111" => data_out <= rom_array(15191);
		when "0011101101011000" => data_out <= rom_array(15192);
		when "0011101101011001" => data_out <= rom_array(15193);
		when "0011101101011010" => data_out <= rom_array(15194);
		when "0011101101011011" => data_out <= rom_array(15195);
		when "0011101101011100" => data_out <= rom_array(15196);
		when "0011101101011101" => data_out <= rom_array(15197);
		when "0011101101011110" => data_out <= rom_array(15198);
		when "0011101101011111" => data_out <= rom_array(15199);
		when "0011101101100000" => data_out <= rom_array(15200);
		when "0011101101100001" => data_out <= rom_array(15201);
		when "0011101101100010" => data_out <= rom_array(15202);
		when "0011101101100011" => data_out <= rom_array(15203);
		when "0011101101100100" => data_out <= rom_array(15204);
		when "0011101101100101" => data_out <= rom_array(15205);
		when "0011101101100110" => data_out <= rom_array(15206);
		when "0011101101100111" => data_out <= rom_array(15207);
		when "0011101101101000" => data_out <= rom_array(15208);
		when "0011101101101001" => data_out <= rom_array(15209);
		when "0011101101101010" => data_out <= rom_array(15210);
		when "0011101101101011" => data_out <= rom_array(15211);
		when "0011101101101100" => data_out <= rom_array(15212);
		when "0011101101101101" => data_out <= rom_array(15213);
		when "0011101101101110" => data_out <= rom_array(15214);
		when "0011101101101111" => data_out <= rom_array(15215);
		when "0011101101110000" => data_out <= rom_array(15216);
		when "0011101101110001" => data_out <= rom_array(15217);
		when "0011101101110010" => data_out <= rom_array(15218);
		when "0011101101110011" => data_out <= rom_array(15219);
		when "0011101101110100" => data_out <= rom_array(15220);
		when "0011101101110101" => data_out <= rom_array(15221);
		when "0011101101110110" => data_out <= rom_array(15222);
		when "0011101101110111" => data_out <= rom_array(15223);
		when "0011101101111000" => data_out <= rom_array(15224);
		when "0011101101111001" => data_out <= rom_array(15225);
		when "0011101101111010" => data_out <= rom_array(15226);
		when "0011101101111011" => data_out <= rom_array(15227);
		when "0011101101111100" => data_out <= rom_array(15228);
		when "0011101101111101" => data_out <= rom_array(15229);
		when "0011101101111110" => data_out <= rom_array(15230);
		when "0011101101111111" => data_out <= rom_array(15231);
		when "0011101110000000" => data_out <= rom_array(15232);
		when "0011101110000001" => data_out <= rom_array(15233);
		when "0011101110000010" => data_out <= rom_array(15234);
		when "0011101110000011" => data_out <= rom_array(15235);
		when "0011101110000100" => data_out <= rom_array(15236);
		when "0011101110000101" => data_out <= rom_array(15237);
		when "0011101110000110" => data_out <= rom_array(15238);
		when "0011101110000111" => data_out <= rom_array(15239);
		when "0011101110001000" => data_out <= rom_array(15240);
		when "0011101110001001" => data_out <= rom_array(15241);
		when "0011101110001010" => data_out <= rom_array(15242);
		when "0011101110001011" => data_out <= rom_array(15243);
		when "0011101110001100" => data_out <= rom_array(15244);
		when "0011101110001101" => data_out <= rom_array(15245);
		when "0011101110001110" => data_out <= rom_array(15246);
		when "0011101110001111" => data_out <= rom_array(15247);
		when "0011101110010000" => data_out <= rom_array(15248);
		when "0011101110010001" => data_out <= rom_array(15249);
		when "0011101110010010" => data_out <= rom_array(15250);
		when "0011101110010011" => data_out <= rom_array(15251);
		when "0011101110010100" => data_out <= rom_array(15252);
		when "0011101110010101" => data_out <= rom_array(15253);
		when "0011101110010110" => data_out <= rom_array(15254);
		when "0011101110010111" => data_out <= rom_array(15255);
		when "0011101110011000" => data_out <= rom_array(15256);
		when "0011101110011001" => data_out <= rom_array(15257);
		when "0011101110011010" => data_out <= rom_array(15258);
		when "0011101110011011" => data_out <= rom_array(15259);
		when "0011101110011100" => data_out <= rom_array(15260);
		when "0011101110011101" => data_out <= rom_array(15261);
		when "0011101110011110" => data_out <= rom_array(15262);
		when "0011101110011111" => data_out <= rom_array(15263);
		when "0011101110100000" => data_out <= rom_array(15264);
		when "0011101110100001" => data_out <= rom_array(15265);
		when "0011101110100010" => data_out <= rom_array(15266);
		when "0011101110100011" => data_out <= rom_array(15267);
		when "0011101110100100" => data_out <= rom_array(15268);
		when "0011101110100101" => data_out <= rom_array(15269);
		when "0011101110100110" => data_out <= rom_array(15270);
		when "0011101110100111" => data_out <= rom_array(15271);
		when "0011101110101000" => data_out <= rom_array(15272);
		when "0011101110101001" => data_out <= rom_array(15273);
		when "0011101110101010" => data_out <= rom_array(15274);
		when "0011101110101011" => data_out <= rom_array(15275);
		when "0011101110101100" => data_out <= rom_array(15276);
		when "0011101110101101" => data_out <= rom_array(15277);
		when "0011101110101110" => data_out <= rom_array(15278);
		when "0011101110101111" => data_out <= rom_array(15279);
		when "0011101110110000" => data_out <= rom_array(15280);
		when "0011101110110001" => data_out <= rom_array(15281);
		when "0011101110110010" => data_out <= rom_array(15282);
		when "0011101110110011" => data_out <= rom_array(15283);
		when "0011101110110100" => data_out <= rom_array(15284);
		when "0011101110110101" => data_out <= rom_array(15285);
		when "0011101110110110" => data_out <= rom_array(15286);
		when "0011101110110111" => data_out <= rom_array(15287);
		when "0011101110111000" => data_out <= rom_array(15288);
		when "0011101110111001" => data_out <= rom_array(15289);
		when "0011101110111010" => data_out <= rom_array(15290);
		when "0011101110111011" => data_out <= rom_array(15291);
		when "0011101110111100" => data_out <= rom_array(15292);
		when "0011101110111101" => data_out <= rom_array(15293);
		when "0011101110111110" => data_out <= rom_array(15294);
		when "0011101110111111" => data_out <= rom_array(15295);
		when "0011101111000000" => data_out <= rom_array(15296);
		when "0011101111000001" => data_out <= rom_array(15297);
		when "0011101111000010" => data_out <= rom_array(15298);
		when "0011101111000011" => data_out <= rom_array(15299);
		when "0011101111000100" => data_out <= rom_array(15300);
		when "0011101111000101" => data_out <= rom_array(15301);
		when "0011101111000110" => data_out <= rom_array(15302);
		when "0011101111000111" => data_out <= rom_array(15303);
		when "0011101111001000" => data_out <= rom_array(15304);
		when "0011101111001001" => data_out <= rom_array(15305);
		when "0011101111001010" => data_out <= rom_array(15306);
		when "0011101111001011" => data_out <= rom_array(15307);
		when "0011101111001100" => data_out <= rom_array(15308);
		when "0011101111001101" => data_out <= rom_array(15309);
		when "0011101111001110" => data_out <= rom_array(15310);
		when "0011101111001111" => data_out <= rom_array(15311);
		when "0011101111010000" => data_out <= rom_array(15312);
		when "0011101111010001" => data_out <= rom_array(15313);
		when "0011101111010010" => data_out <= rom_array(15314);
		when "0011101111010011" => data_out <= rom_array(15315);
		when "0011101111010100" => data_out <= rom_array(15316);
		when "0011101111010101" => data_out <= rom_array(15317);
		when "0011101111010110" => data_out <= rom_array(15318);
		when "0011101111010111" => data_out <= rom_array(15319);
		when "0011101111011000" => data_out <= rom_array(15320);
		when "0011101111011001" => data_out <= rom_array(15321);
		when "0011101111011010" => data_out <= rom_array(15322);
		when "0011101111011011" => data_out <= rom_array(15323);
		when "0011101111011100" => data_out <= rom_array(15324);
		when "0011101111011101" => data_out <= rom_array(15325);
		when "0011101111011110" => data_out <= rom_array(15326);
		when "0011101111011111" => data_out <= rom_array(15327);
		when "0011101111100000" => data_out <= rom_array(15328);
		when "0011101111100001" => data_out <= rom_array(15329);
		when "0011101111100010" => data_out <= rom_array(15330);
		when "0011101111100011" => data_out <= rom_array(15331);
		when "0011101111100100" => data_out <= rom_array(15332);
		when "0011101111100101" => data_out <= rom_array(15333);
		when "0011101111100110" => data_out <= rom_array(15334);
		when "0011101111100111" => data_out <= rom_array(15335);
		when "0011101111101000" => data_out <= rom_array(15336);
		when "0011101111101001" => data_out <= rom_array(15337);
		when "0011101111101010" => data_out <= rom_array(15338);
		when "0011101111101011" => data_out <= rom_array(15339);
		when "0011101111101100" => data_out <= rom_array(15340);
		when "0011101111101101" => data_out <= rom_array(15341);
		when "0011101111101110" => data_out <= rom_array(15342);
		when "0011101111101111" => data_out <= rom_array(15343);
		when "0011101111110000" => data_out <= rom_array(15344);
		when "0011101111110001" => data_out <= rom_array(15345);
		when "0011101111110010" => data_out <= rom_array(15346);
		when "0011101111110011" => data_out <= rom_array(15347);
		when "0011101111110100" => data_out <= rom_array(15348);
		when "0011101111110101" => data_out <= rom_array(15349);
		when "0011101111110110" => data_out <= rom_array(15350);
		when "0011101111110111" => data_out <= rom_array(15351);
		when "0011101111111000" => data_out <= rom_array(15352);
		when "0011101111111001" => data_out <= rom_array(15353);
		when "0011101111111010" => data_out <= rom_array(15354);
		when "0011101111111011" => data_out <= rom_array(15355);
		when "0011101111111100" => data_out <= rom_array(15356);
		when "0011101111111101" => data_out <= rom_array(15357);
		when "0011101111111110" => data_out <= rom_array(15358);
		when "0011101111111111" => data_out <= rom_array(15359);
		when "0011110000000000" => data_out <= rom_array(15360);
		when "0011110000000001" => data_out <= rom_array(15361);
		when "0011110000000010" => data_out <= rom_array(15362);
		when "0011110000000011" => data_out <= rom_array(15363);
		when "0011110000000100" => data_out <= rom_array(15364);
		when "0011110000000101" => data_out <= rom_array(15365);
		when "0011110000000110" => data_out <= rom_array(15366);
		when "0011110000000111" => data_out <= rom_array(15367);
		when "0011110000001000" => data_out <= rom_array(15368);
		when "0011110000001001" => data_out <= rom_array(15369);
		when "0011110000001010" => data_out <= rom_array(15370);
		when "0011110000001011" => data_out <= rom_array(15371);
		when "0011110000001100" => data_out <= rom_array(15372);
		when "0011110000001101" => data_out <= rom_array(15373);
		when "0011110000001110" => data_out <= rom_array(15374);
		when "0011110000001111" => data_out <= rom_array(15375);
		when "0011110000010000" => data_out <= rom_array(15376);
		when "0011110000010001" => data_out <= rom_array(15377);
		when "0011110000010010" => data_out <= rom_array(15378);
		when "0011110000010011" => data_out <= rom_array(15379);
		when "0011110000010100" => data_out <= rom_array(15380);
		when "0011110000010101" => data_out <= rom_array(15381);
		when "0011110000010110" => data_out <= rom_array(15382);
		when "0011110000010111" => data_out <= rom_array(15383);
		when "0011110000011000" => data_out <= rom_array(15384);
		when "0011110000011001" => data_out <= rom_array(15385);
		when "0011110000011010" => data_out <= rom_array(15386);
		when "0011110000011011" => data_out <= rom_array(15387);
		when "0011110000011100" => data_out <= rom_array(15388);
		when "0011110000011101" => data_out <= rom_array(15389);
		when "0011110000011110" => data_out <= rom_array(15390);
		when "0011110000011111" => data_out <= rom_array(15391);
		when "0011110000100000" => data_out <= rom_array(15392);
		when "0011110000100001" => data_out <= rom_array(15393);
		when "0011110000100010" => data_out <= rom_array(15394);
		when "0011110000100011" => data_out <= rom_array(15395);
		when "0011110000100100" => data_out <= rom_array(15396);
		when "0011110000100101" => data_out <= rom_array(15397);
		when "0011110000100110" => data_out <= rom_array(15398);
		when "0011110000100111" => data_out <= rom_array(15399);
		when "0011110000101000" => data_out <= rom_array(15400);
		when "0011110000101001" => data_out <= rom_array(15401);
		when "0011110000101010" => data_out <= rom_array(15402);
		when "0011110000101011" => data_out <= rom_array(15403);
		when "0011110000101100" => data_out <= rom_array(15404);
		when "0011110000101101" => data_out <= rom_array(15405);
		when "0011110000101110" => data_out <= rom_array(15406);
		when "0011110000101111" => data_out <= rom_array(15407);
		when "0011110000110000" => data_out <= rom_array(15408);
		when "0011110000110001" => data_out <= rom_array(15409);
		when "0011110000110010" => data_out <= rom_array(15410);
		when "0011110000110011" => data_out <= rom_array(15411);
		when "0011110000110100" => data_out <= rom_array(15412);
		when "0011110000110101" => data_out <= rom_array(15413);
		when "0011110000110110" => data_out <= rom_array(15414);
		when "0011110000110111" => data_out <= rom_array(15415);
		when "0011110000111000" => data_out <= rom_array(15416);
		when "0011110000111001" => data_out <= rom_array(15417);
		when "0011110000111010" => data_out <= rom_array(15418);
		when "0011110000111011" => data_out <= rom_array(15419);
		when "0011110000111100" => data_out <= rom_array(15420);
		when "0011110000111101" => data_out <= rom_array(15421);
		when "0011110000111110" => data_out <= rom_array(15422);
		when "0011110000111111" => data_out <= rom_array(15423);
		when "0011110001000000" => data_out <= rom_array(15424);
		when "0011110001000001" => data_out <= rom_array(15425);
		when "0011110001000010" => data_out <= rom_array(15426);
		when "0011110001000011" => data_out <= rom_array(15427);
		when "0011110001000100" => data_out <= rom_array(15428);
		when "0011110001000101" => data_out <= rom_array(15429);
		when "0011110001000110" => data_out <= rom_array(15430);
		when "0011110001000111" => data_out <= rom_array(15431);
		when "0011110001001000" => data_out <= rom_array(15432);
		when "0011110001001001" => data_out <= rom_array(15433);
		when "0011110001001010" => data_out <= rom_array(15434);
		when "0011110001001011" => data_out <= rom_array(15435);
		when "0011110001001100" => data_out <= rom_array(15436);
		when "0011110001001101" => data_out <= rom_array(15437);
		when "0011110001001110" => data_out <= rom_array(15438);
		when "0011110001001111" => data_out <= rom_array(15439);
		when "0011110001010000" => data_out <= rom_array(15440);
		when "0011110001010001" => data_out <= rom_array(15441);
		when "0011110001010010" => data_out <= rom_array(15442);
		when "0011110001010011" => data_out <= rom_array(15443);
		when "0011110001010100" => data_out <= rom_array(15444);
		when "0011110001010101" => data_out <= rom_array(15445);
		when "0011110001010110" => data_out <= rom_array(15446);
		when "0011110001010111" => data_out <= rom_array(15447);
		when "0011110001011000" => data_out <= rom_array(15448);
		when "0011110001011001" => data_out <= rom_array(15449);
		when "0011110001011010" => data_out <= rom_array(15450);
		when "0011110001011011" => data_out <= rom_array(15451);
		when "0011110001011100" => data_out <= rom_array(15452);
		when "0011110001011101" => data_out <= rom_array(15453);
		when "0011110001011110" => data_out <= rom_array(15454);
		when "0011110001011111" => data_out <= rom_array(15455);
		when "0011110001100000" => data_out <= rom_array(15456);
		when "0011110001100001" => data_out <= rom_array(15457);
		when "0011110001100010" => data_out <= rom_array(15458);
		when "0011110001100011" => data_out <= rom_array(15459);
		when "0011110001100100" => data_out <= rom_array(15460);
		when "0011110001100101" => data_out <= rom_array(15461);
		when "0011110001100110" => data_out <= rom_array(15462);
		when "0011110001100111" => data_out <= rom_array(15463);
		when "0011110001101000" => data_out <= rom_array(15464);
		when "0011110001101001" => data_out <= rom_array(15465);
		when "0011110001101010" => data_out <= rom_array(15466);
		when "0011110001101011" => data_out <= rom_array(15467);
		when "0011110001101100" => data_out <= rom_array(15468);
		when "0011110001101101" => data_out <= rom_array(15469);
		when "0011110001101110" => data_out <= rom_array(15470);
		when "0011110001101111" => data_out <= rom_array(15471);
		when "0011110001110000" => data_out <= rom_array(15472);
		when "0011110001110001" => data_out <= rom_array(15473);
		when "0011110001110010" => data_out <= rom_array(15474);
		when "0011110001110011" => data_out <= rom_array(15475);
		when "0011110001110100" => data_out <= rom_array(15476);
		when "0011110001110101" => data_out <= rom_array(15477);
		when "0011110001110110" => data_out <= rom_array(15478);
		when "0011110001110111" => data_out <= rom_array(15479);
		when "0011110001111000" => data_out <= rom_array(15480);
		when "0011110001111001" => data_out <= rom_array(15481);
		when "0011110001111010" => data_out <= rom_array(15482);
		when "0011110001111011" => data_out <= rom_array(15483);
		when "0011110001111100" => data_out <= rom_array(15484);
		when "0011110001111101" => data_out <= rom_array(15485);
		when "0011110001111110" => data_out <= rom_array(15486);
		when "0011110001111111" => data_out <= rom_array(15487);
		when "0011110010000000" => data_out <= rom_array(15488);
		when "0011110010000001" => data_out <= rom_array(15489);
		when "0011110010000010" => data_out <= rom_array(15490);
		when "0011110010000011" => data_out <= rom_array(15491);
		when "0011110010000100" => data_out <= rom_array(15492);
		when "0011110010000101" => data_out <= rom_array(15493);
		when "0011110010000110" => data_out <= rom_array(15494);
		when "0011110010000111" => data_out <= rom_array(15495);
		when "0011110010001000" => data_out <= rom_array(15496);
		when "0011110010001001" => data_out <= rom_array(15497);
		when "0011110010001010" => data_out <= rom_array(15498);
		when "0011110010001011" => data_out <= rom_array(15499);
		when "0011110010001100" => data_out <= rom_array(15500);
		when "0011110010001101" => data_out <= rom_array(15501);
		when "0011110010001110" => data_out <= rom_array(15502);
		when "0011110010001111" => data_out <= rom_array(15503);
		when "0011110010010000" => data_out <= rom_array(15504);
		when "0011110010010001" => data_out <= rom_array(15505);
		when "0011110010010010" => data_out <= rom_array(15506);
		when "0011110010010011" => data_out <= rom_array(15507);
		when "0011110010010100" => data_out <= rom_array(15508);
		when "0011110010010101" => data_out <= rom_array(15509);
		when "0011110010010110" => data_out <= rom_array(15510);
		when "0011110010010111" => data_out <= rom_array(15511);
		when "0011110010011000" => data_out <= rom_array(15512);
		when "0011110010011001" => data_out <= rom_array(15513);
		when "0011110010011010" => data_out <= rom_array(15514);
		when "0011110010011011" => data_out <= rom_array(15515);
		when "0011110010011100" => data_out <= rom_array(15516);
		when "0011110010011101" => data_out <= rom_array(15517);
		when "0011110010011110" => data_out <= rom_array(15518);
		when "0011110010011111" => data_out <= rom_array(15519);
		when "0011110010100000" => data_out <= rom_array(15520);
		when "0011110010100001" => data_out <= rom_array(15521);
		when "0011110010100010" => data_out <= rom_array(15522);
		when "0011110010100011" => data_out <= rom_array(15523);
		when "0011110010100100" => data_out <= rom_array(15524);
		when "0011110010100101" => data_out <= rom_array(15525);
		when "0011110010100110" => data_out <= rom_array(15526);
		when "0011110010100111" => data_out <= rom_array(15527);
		when "0011110010101000" => data_out <= rom_array(15528);
		when "0011110010101001" => data_out <= rom_array(15529);
		when "0011110010101010" => data_out <= rom_array(15530);
		when "0011110010101011" => data_out <= rom_array(15531);
		when "0011110010101100" => data_out <= rom_array(15532);
		when "0011110010101101" => data_out <= rom_array(15533);
		when "0011110010101110" => data_out <= rom_array(15534);
		when "0011110010101111" => data_out <= rom_array(15535);
		when "0011110010110000" => data_out <= rom_array(15536);
		when "0011110010110001" => data_out <= rom_array(15537);
		when "0011110010110010" => data_out <= rom_array(15538);
		when "0011110010110011" => data_out <= rom_array(15539);
		when "0011110010110100" => data_out <= rom_array(15540);
		when "0011110010110101" => data_out <= rom_array(15541);
		when "0011110010110110" => data_out <= rom_array(15542);
		when "0011110010110111" => data_out <= rom_array(15543);
		when "0011110010111000" => data_out <= rom_array(15544);
		when "0011110010111001" => data_out <= rom_array(15545);
		when "0011110010111010" => data_out <= rom_array(15546);
		when "0011110010111011" => data_out <= rom_array(15547);
		when "0011110010111100" => data_out <= rom_array(15548);
		when "0011110010111101" => data_out <= rom_array(15549);
		when "0011110010111110" => data_out <= rom_array(15550);
		when "0011110010111111" => data_out <= rom_array(15551);
		when "0011110011000000" => data_out <= rom_array(15552);
		when "0011110011000001" => data_out <= rom_array(15553);
		when "0011110011000010" => data_out <= rom_array(15554);
		when "0011110011000011" => data_out <= rom_array(15555);
		when "0011110011000100" => data_out <= rom_array(15556);
		when "0011110011000101" => data_out <= rom_array(15557);
		when "0011110011000110" => data_out <= rom_array(15558);
		when "0011110011000111" => data_out <= rom_array(15559);
		when "0011110011001000" => data_out <= rom_array(15560);
		when "0011110011001001" => data_out <= rom_array(15561);
		when "0011110011001010" => data_out <= rom_array(15562);
		when "0011110011001011" => data_out <= rom_array(15563);
		when "0011110011001100" => data_out <= rom_array(15564);
		when "0011110011001101" => data_out <= rom_array(15565);
		when "0011110011001110" => data_out <= rom_array(15566);
		when "0011110011001111" => data_out <= rom_array(15567);
		when "0011110011010000" => data_out <= rom_array(15568);
		when "0011110011010001" => data_out <= rom_array(15569);
		when "0011110011010010" => data_out <= rom_array(15570);
		when "0011110011010011" => data_out <= rom_array(15571);
		when "0011110011010100" => data_out <= rom_array(15572);
		when "0011110011010101" => data_out <= rom_array(15573);
		when "0011110011010110" => data_out <= rom_array(15574);
		when "0011110011010111" => data_out <= rom_array(15575);
		when "0011110011011000" => data_out <= rom_array(15576);
		when "0011110011011001" => data_out <= rom_array(15577);
		when "0011110011011010" => data_out <= rom_array(15578);
		when "0011110011011011" => data_out <= rom_array(15579);
		when "0011110011011100" => data_out <= rom_array(15580);
		when "0011110011011101" => data_out <= rom_array(15581);
		when "0011110011011110" => data_out <= rom_array(15582);
		when "0011110011011111" => data_out <= rom_array(15583);
		when "0011110011100000" => data_out <= rom_array(15584);
		when "0011110011100001" => data_out <= rom_array(15585);
		when "0011110011100010" => data_out <= rom_array(15586);
		when "0011110011100011" => data_out <= rom_array(15587);
		when "0011110011100100" => data_out <= rom_array(15588);
		when "0011110011100101" => data_out <= rom_array(15589);
		when "0011110011100110" => data_out <= rom_array(15590);
		when "0011110011100111" => data_out <= rom_array(15591);
		when "0011110011101000" => data_out <= rom_array(15592);
		when "0011110011101001" => data_out <= rom_array(15593);
		when "0011110011101010" => data_out <= rom_array(15594);
		when "0011110011101011" => data_out <= rom_array(15595);
		when "0011110011101100" => data_out <= rom_array(15596);
		when "0011110011101101" => data_out <= rom_array(15597);
		when "0011110011101110" => data_out <= rom_array(15598);
		when "0011110011101111" => data_out <= rom_array(15599);
		when "0011110011110000" => data_out <= rom_array(15600);
		when "0011110011110001" => data_out <= rom_array(15601);
		when "0011110011110010" => data_out <= rom_array(15602);
		when "0011110011110011" => data_out <= rom_array(15603);
		when "0011110011110100" => data_out <= rom_array(15604);
		when "0011110011110101" => data_out <= rom_array(15605);
		when "0011110011110110" => data_out <= rom_array(15606);
		when "0011110011110111" => data_out <= rom_array(15607);
		when "0011110011111000" => data_out <= rom_array(15608);
		when "0011110011111001" => data_out <= rom_array(15609);
		when "0011110011111010" => data_out <= rom_array(15610);
		when "0011110011111011" => data_out <= rom_array(15611);
		when "0011110011111100" => data_out <= rom_array(15612);
		when "0011110011111101" => data_out <= rom_array(15613);
		when "0011110011111110" => data_out <= rom_array(15614);
		when "0011110011111111" => data_out <= rom_array(15615);
		when "0011110100000000" => data_out <= rom_array(15616);
		when "0011110100000001" => data_out <= rom_array(15617);
		when "0011110100000010" => data_out <= rom_array(15618);
		when "0011110100000011" => data_out <= rom_array(15619);
		when "0011110100000100" => data_out <= rom_array(15620);
		when "0011110100000101" => data_out <= rom_array(15621);
		when "0011110100000110" => data_out <= rom_array(15622);
		when "0011110100000111" => data_out <= rom_array(15623);
		when "0011110100001000" => data_out <= rom_array(15624);
		when "0011110100001001" => data_out <= rom_array(15625);
		when "0011110100001010" => data_out <= rom_array(15626);
		when "0011110100001011" => data_out <= rom_array(15627);
		when "0011110100001100" => data_out <= rom_array(15628);
		when "0011110100001101" => data_out <= rom_array(15629);
		when "0011110100001110" => data_out <= rom_array(15630);
		when "0011110100001111" => data_out <= rom_array(15631);
		when "0011110100010000" => data_out <= rom_array(15632);
		when "0011110100010001" => data_out <= rom_array(15633);
		when "0011110100010010" => data_out <= rom_array(15634);
		when "0011110100010011" => data_out <= rom_array(15635);
		when "0011110100010100" => data_out <= rom_array(15636);
		when "0011110100010101" => data_out <= rom_array(15637);
		when "0011110100010110" => data_out <= rom_array(15638);
		when "0011110100010111" => data_out <= rom_array(15639);
		when "0011110100011000" => data_out <= rom_array(15640);
		when "0011110100011001" => data_out <= rom_array(15641);
		when "0011110100011010" => data_out <= rom_array(15642);
		when "0011110100011011" => data_out <= rom_array(15643);
		when "0011110100011100" => data_out <= rom_array(15644);
		when "0011110100011101" => data_out <= rom_array(15645);
		when "0011110100011110" => data_out <= rom_array(15646);
		when "0011110100011111" => data_out <= rom_array(15647);
		when "0011110100100000" => data_out <= rom_array(15648);
		when "0011110100100001" => data_out <= rom_array(15649);
		when "0011110100100010" => data_out <= rom_array(15650);
		when "0011110100100011" => data_out <= rom_array(15651);
		when "0011110100100100" => data_out <= rom_array(15652);
		when "0011110100100101" => data_out <= rom_array(15653);
		when "0011110100100110" => data_out <= rom_array(15654);
		when "0011110100100111" => data_out <= rom_array(15655);
		when "0011110100101000" => data_out <= rom_array(15656);
		when "0011110100101001" => data_out <= rom_array(15657);
		when "0011110100101010" => data_out <= rom_array(15658);
		when "0011110100101011" => data_out <= rom_array(15659);
		when "0011110100101100" => data_out <= rom_array(15660);
		when "0011110100101101" => data_out <= rom_array(15661);
		when "0011110100101110" => data_out <= rom_array(15662);
		when "0011110100101111" => data_out <= rom_array(15663);
		when "0011110100110000" => data_out <= rom_array(15664);
		when "0011110100110001" => data_out <= rom_array(15665);
		when "0011110100110010" => data_out <= rom_array(15666);
		when "0011110100110011" => data_out <= rom_array(15667);
		when "0011110100110100" => data_out <= rom_array(15668);
		when "0011110100110101" => data_out <= rom_array(15669);
		when "0011110100110110" => data_out <= rom_array(15670);
		when "0011110100110111" => data_out <= rom_array(15671);
		when "0011110100111000" => data_out <= rom_array(15672);
		when "0011110100111001" => data_out <= rom_array(15673);
		when "0011110100111010" => data_out <= rom_array(15674);
		when "0011110100111011" => data_out <= rom_array(15675);
		when "0011110100111100" => data_out <= rom_array(15676);
		when "0011110100111101" => data_out <= rom_array(15677);
		when "0011110100111110" => data_out <= rom_array(15678);
		when "0011110100111111" => data_out <= rom_array(15679);
		when "0011110101000000" => data_out <= rom_array(15680);
		when "0011110101000001" => data_out <= rom_array(15681);
		when "0011110101000010" => data_out <= rom_array(15682);
		when "0011110101000011" => data_out <= rom_array(15683);
		when "0011110101000100" => data_out <= rom_array(15684);
		when "0011110101000101" => data_out <= rom_array(15685);
		when "0011110101000110" => data_out <= rom_array(15686);
		when "0011110101000111" => data_out <= rom_array(15687);
		when "0011110101001000" => data_out <= rom_array(15688);
		when "0011110101001001" => data_out <= rom_array(15689);
		when "0011110101001010" => data_out <= rom_array(15690);
		when "0011110101001011" => data_out <= rom_array(15691);
		when "0011110101001100" => data_out <= rom_array(15692);
		when "0011110101001101" => data_out <= rom_array(15693);
		when "0011110101001110" => data_out <= rom_array(15694);
		when "0011110101001111" => data_out <= rom_array(15695);
		when "0011110101010000" => data_out <= rom_array(15696);
		when "0011110101010001" => data_out <= rom_array(15697);
		when "0011110101010010" => data_out <= rom_array(15698);
		when "0011110101010011" => data_out <= rom_array(15699);
		when "0011110101010100" => data_out <= rom_array(15700);
		when "0011110101010101" => data_out <= rom_array(15701);
		when "0011110101010110" => data_out <= rom_array(15702);
		when "0011110101010111" => data_out <= rom_array(15703);
		when "0011110101011000" => data_out <= rom_array(15704);
		when "0011110101011001" => data_out <= rom_array(15705);
		when "0011110101011010" => data_out <= rom_array(15706);
		when "0011110101011011" => data_out <= rom_array(15707);
		when "0011110101011100" => data_out <= rom_array(15708);
		when "0011110101011101" => data_out <= rom_array(15709);
		when "0011110101011110" => data_out <= rom_array(15710);
		when "0011110101011111" => data_out <= rom_array(15711);
		when "0011110101100000" => data_out <= rom_array(15712);
		when "0011110101100001" => data_out <= rom_array(15713);
		when "0011110101100010" => data_out <= rom_array(15714);
		when "0011110101100011" => data_out <= rom_array(15715);
		when "0011110101100100" => data_out <= rom_array(15716);
		when "0011110101100101" => data_out <= rom_array(15717);
		when "0011110101100110" => data_out <= rom_array(15718);
		when "0011110101100111" => data_out <= rom_array(15719);
		when "0011110101101000" => data_out <= rom_array(15720);
		when "0011110101101001" => data_out <= rom_array(15721);
		when "0011110101101010" => data_out <= rom_array(15722);
		when "0011110101101011" => data_out <= rom_array(15723);
		when "0011110101101100" => data_out <= rom_array(15724);
		when "0011110101101101" => data_out <= rom_array(15725);
		when "0011110101101110" => data_out <= rom_array(15726);
		when "0011110101101111" => data_out <= rom_array(15727);
		when "0011110101110000" => data_out <= rom_array(15728);
		when "0011110101110001" => data_out <= rom_array(15729);
		when "0011110101110010" => data_out <= rom_array(15730);
		when "0011110101110011" => data_out <= rom_array(15731);
		when "0011110101110100" => data_out <= rom_array(15732);
		when "0011110101110101" => data_out <= rom_array(15733);
		when "0011110101110110" => data_out <= rom_array(15734);
		when "0011110101110111" => data_out <= rom_array(15735);
		when "0011110101111000" => data_out <= rom_array(15736);
		when "0011110101111001" => data_out <= rom_array(15737);
		when "0011110101111010" => data_out <= rom_array(15738);
		when "0011110101111011" => data_out <= rom_array(15739);
		when "0011110101111100" => data_out <= rom_array(15740);
		when "0011110101111101" => data_out <= rom_array(15741);
		when "0011110101111110" => data_out <= rom_array(15742);
		when "0011110101111111" => data_out <= rom_array(15743);
		when "0011110110000000" => data_out <= rom_array(15744);
		when "0011110110000001" => data_out <= rom_array(15745);
		when "0011110110000010" => data_out <= rom_array(15746);
		when "0011110110000011" => data_out <= rom_array(15747);
		when "0011110110000100" => data_out <= rom_array(15748);
		when "0011110110000101" => data_out <= rom_array(15749);
		when "0011110110000110" => data_out <= rom_array(15750);
		when "0011110110000111" => data_out <= rom_array(15751);
		when "0011110110001000" => data_out <= rom_array(15752);
		when "0011110110001001" => data_out <= rom_array(15753);
		when "0011110110001010" => data_out <= rom_array(15754);
		when "0011110110001011" => data_out <= rom_array(15755);
		when "0011110110001100" => data_out <= rom_array(15756);
		when "0011110110001101" => data_out <= rom_array(15757);
		when "0011110110001110" => data_out <= rom_array(15758);
		when "0011110110001111" => data_out <= rom_array(15759);
		when "0011110110010000" => data_out <= rom_array(15760);
		when "0011110110010001" => data_out <= rom_array(15761);
		when "0011110110010010" => data_out <= rom_array(15762);
		when "0011110110010011" => data_out <= rom_array(15763);
		when "0011110110010100" => data_out <= rom_array(15764);
		when "0011110110010101" => data_out <= rom_array(15765);
		when "0011110110010110" => data_out <= rom_array(15766);
		when "0011110110010111" => data_out <= rom_array(15767);
		when "0011110110011000" => data_out <= rom_array(15768);
		when "0011110110011001" => data_out <= rom_array(15769);
		when "0011110110011010" => data_out <= rom_array(15770);
		when "0011110110011011" => data_out <= rom_array(15771);
		when "0011110110011100" => data_out <= rom_array(15772);
		when "0011110110011101" => data_out <= rom_array(15773);
		when "0011110110011110" => data_out <= rom_array(15774);
		when "0011110110011111" => data_out <= rom_array(15775);
		when "0011110110100000" => data_out <= rom_array(15776);
		when "0011110110100001" => data_out <= rom_array(15777);
		when "0011110110100010" => data_out <= rom_array(15778);
		when "0011110110100011" => data_out <= rom_array(15779);
		when "0011110110100100" => data_out <= rom_array(15780);
		when "0011110110100101" => data_out <= rom_array(15781);
		when "0011110110100110" => data_out <= rom_array(15782);
		when "0011110110100111" => data_out <= rom_array(15783);
		when "0011110110101000" => data_out <= rom_array(15784);
		when "0011110110101001" => data_out <= rom_array(15785);
		when "0011110110101010" => data_out <= rom_array(15786);
		when "0011110110101011" => data_out <= rom_array(15787);
		when "0011110110101100" => data_out <= rom_array(15788);
		when "0011110110101101" => data_out <= rom_array(15789);
		when "0011110110101110" => data_out <= rom_array(15790);
		when "0011110110101111" => data_out <= rom_array(15791);
		when "0011110110110000" => data_out <= rom_array(15792);
		when "0011110110110001" => data_out <= rom_array(15793);
		when "0011110110110010" => data_out <= rom_array(15794);
		when "0011110110110011" => data_out <= rom_array(15795);
		when "0011110110110100" => data_out <= rom_array(15796);
		when "0011110110110101" => data_out <= rom_array(15797);
		when "0011110110110110" => data_out <= rom_array(15798);
		when "0011110110110111" => data_out <= rom_array(15799);
		when "0011110110111000" => data_out <= rom_array(15800);
		when "0011110110111001" => data_out <= rom_array(15801);
		when "0011110110111010" => data_out <= rom_array(15802);
		when "0011110110111011" => data_out <= rom_array(15803);
		when "0011110110111100" => data_out <= rom_array(15804);
		when "0011110110111101" => data_out <= rom_array(15805);
		when "0011110110111110" => data_out <= rom_array(15806);
		when "0011110110111111" => data_out <= rom_array(15807);
		when "0011110111000000" => data_out <= rom_array(15808);
		when "0011110111000001" => data_out <= rom_array(15809);
		when "0011110111000010" => data_out <= rom_array(15810);
		when "0011110111000011" => data_out <= rom_array(15811);
		when "0011110111000100" => data_out <= rom_array(15812);
		when "0011110111000101" => data_out <= rom_array(15813);
		when "0011110111000110" => data_out <= rom_array(15814);
		when "0011110111000111" => data_out <= rom_array(15815);
		when "0011110111001000" => data_out <= rom_array(15816);
		when "0011110111001001" => data_out <= rom_array(15817);
		when "0011110111001010" => data_out <= rom_array(15818);
		when "0011110111001011" => data_out <= rom_array(15819);
		when "0011110111001100" => data_out <= rom_array(15820);
		when "0011110111001101" => data_out <= rom_array(15821);
		when "0011110111001110" => data_out <= rom_array(15822);
		when "0011110111001111" => data_out <= rom_array(15823);
		when "0011110111010000" => data_out <= rom_array(15824);
		when "0011110111010001" => data_out <= rom_array(15825);
		when "0011110111010010" => data_out <= rom_array(15826);
		when "0011110111010011" => data_out <= rom_array(15827);
		when "0011110111010100" => data_out <= rom_array(15828);
		when "0011110111010101" => data_out <= rom_array(15829);
		when "0011110111010110" => data_out <= rom_array(15830);
		when "0011110111010111" => data_out <= rom_array(15831);
		when "0011110111011000" => data_out <= rom_array(15832);
		when "0011110111011001" => data_out <= rom_array(15833);
		when "0011110111011010" => data_out <= rom_array(15834);
		when "0011110111011011" => data_out <= rom_array(15835);
		when "0011110111011100" => data_out <= rom_array(15836);
		when "0011110111011101" => data_out <= rom_array(15837);
		when "0011110111011110" => data_out <= rom_array(15838);
		when "0011110111011111" => data_out <= rom_array(15839);
		when "0011110111100000" => data_out <= rom_array(15840);
		when "0011110111100001" => data_out <= rom_array(15841);
		when "0011110111100010" => data_out <= rom_array(15842);
		when "0011110111100011" => data_out <= rom_array(15843);
		when "0011110111100100" => data_out <= rom_array(15844);
		when "0011110111100101" => data_out <= rom_array(15845);
		when "0011110111100110" => data_out <= rom_array(15846);
		when "0011110111100111" => data_out <= rom_array(15847);
		when "0011110111101000" => data_out <= rom_array(15848);
		when "0011110111101001" => data_out <= rom_array(15849);
		when "0011110111101010" => data_out <= rom_array(15850);
		when "0011110111101011" => data_out <= rom_array(15851);
		when "0011110111101100" => data_out <= rom_array(15852);
		when "0011110111101101" => data_out <= rom_array(15853);
		when "0011110111101110" => data_out <= rom_array(15854);
		when "0011110111101111" => data_out <= rom_array(15855);
		when "0011110111110000" => data_out <= rom_array(15856);
		when "0011110111110001" => data_out <= rom_array(15857);
		when "0011110111110010" => data_out <= rom_array(15858);
		when "0011110111110011" => data_out <= rom_array(15859);
		when "0011110111110100" => data_out <= rom_array(15860);
		when "0011110111110101" => data_out <= rom_array(15861);
		when "0011110111110110" => data_out <= rom_array(15862);
		when "0011110111110111" => data_out <= rom_array(15863);
		when "0011110111111000" => data_out <= rom_array(15864);
		when "0011110111111001" => data_out <= rom_array(15865);
		when "0011110111111010" => data_out <= rom_array(15866);
		when "0011110111111011" => data_out <= rom_array(15867);
		when "0011110111111100" => data_out <= rom_array(15868);
		when "0011110111111101" => data_out <= rom_array(15869);
		when "0011110111111110" => data_out <= rom_array(15870);
		when "0011110111111111" => data_out <= rom_array(15871);
		when "0011111000000000" => data_out <= rom_array(15872);
		when "0011111000000001" => data_out <= rom_array(15873);
		when "0011111000000010" => data_out <= rom_array(15874);
		when "0011111000000011" => data_out <= rom_array(15875);
		when "0011111000000100" => data_out <= rom_array(15876);
		when "0011111000000101" => data_out <= rom_array(15877);
		when "0011111000000110" => data_out <= rom_array(15878);
		when "0011111000000111" => data_out <= rom_array(15879);
		when "0011111000001000" => data_out <= rom_array(15880);
		when "0011111000001001" => data_out <= rom_array(15881);
		when "0011111000001010" => data_out <= rom_array(15882);
		when "0011111000001011" => data_out <= rom_array(15883);
		when "0011111000001100" => data_out <= rom_array(15884);
		when "0011111000001101" => data_out <= rom_array(15885);
		when "0011111000001110" => data_out <= rom_array(15886);
		when "0011111000001111" => data_out <= rom_array(15887);
		when "0011111000010000" => data_out <= rom_array(15888);
		when "0011111000010001" => data_out <= rom_array(15889);
		when "0011111000010010" => data_out <= rom_array(15890);
		when "0011111000010011" => data_out <= rom_array(15891);
		when "0011111000010100" => data_out <= rom_array(15892);
		when "0011111000010101" => data_out <= rom_array(15893);
		when "0011111000010110" => data_out <= rom_array(15894);
		when "0011111000010111" => data_out <= rom_array(15895);
		when "0011111000011000" => data_out <= rom_array(15896);
		when "0011111000011001" => data_out <= rom_array(15897);
		when "0011111000011010" => data_out <= rom_array(15898);
		when "0011111000011011" => data_out <= rom_array(15899);
		when "0011111000011100" => data_out <= rom_array(15900);
		when "0011111000011101" => data_out <= rom_array(15901);
		when "0011111000011110" => data_out <= rom_array(15902);
		when "0011111000011111" => data_out <= rom_array(15903);
		when "0011111000100000" => data_out <= rom_array(15904);
		when "0011111000100001" => data_out <= rom_array(15905);
		when "0011111000100010" => data_out <= rom_array(15906);
		when "0011111000100011" => data_out <= rom_array(15907);
		when "0011111000100100" => data_out <= rom_array(15908);
		when "0011111000100101" => data_out <= rom_array(15909);
		when "0011111000100110" => data_out <= rom_array(15910);
		when "0011111000100111" => data_out <= rom_array(15911);
		when "0011111000101000" => data_out <= rom_array(15912);
		when "0011111000101001" => data_out <= rom_array(15913);
		when "0011111000101010" => data_out <= rom_array(15914);
		when "0011111000101011" => data_out <= rom_array(15915);
		when "0011111000101100" => data_out <= rom_array(15916);
		when "0011111000101101" => data_out <= rom_array(15917);
		when "0011111000101110" => data_out <= rom_array(15918);
		when "0011111000101111" => data_out <= rom_array(15919);
		when "0011111000110000" => data_out <= rom_array(15920);
		when "0011111000110001" => data_out <= rom_array(15921);
		when "0011111000110010" => data_out <= rom_array(15922);
		when "0011111000110011" => data_out <= rom_array(15923);
		when "0011111000110100" => data_out <= rom_array(15924);
		when "0011111000110101" => data_out <= rom_array(15925);
		when "0011111000110110" => data_out <= rom_array(15926);
		when "0011111000110111" => data_out <= rom_array(15927);
		when "0011111000111000" => data_out <= rom_array(15928);
		when "0011111000111001" => data_out <= rom_array(15929);
		when "0011111000111010" => data_out <= rom_array(15930);
		when "0011111000111011" => data_out <= rom_array(15931);
		when "0011111000111100" => data_out <= rom_array(15932);
		when "0011111000111101" => data_out <= rom_array(15933);
		when "0011111000111110" => data_out <= rom_array(15934);
		when "0011111000111111" => data_out <= rom_array(15935);
		when "0011111001000000" => data_out <= rom_array(15936);
		when "0011111001000001" => data_out <= rom_array(15937);
		when "0011111001000010" => data_out <= rom_array(15938);
		when "0011111001000011" => data_out <= rom_array(15939);
		when "0011111001000100" => data_out <= rom_array(15940);
		when "0011111001000101" => data_out <= rom_array(15941);
		when "0011111001000110" => data_out <= rom_array(15942);
		when "0011111001000111" => data_out <= rom_array(15943);
		when "0011111001001000" => data_out <= rom_array(15944);
		when "0011111001001001" => data_out <= rom_array(15945);
		when "0011111001001010" => data_out <= rom_array(15946);
		when "0011111001001011" => data_out <= rom_array(15947);
		when "0011111001001100" => data_out <= rom_array(15948);
		when "0011111001001101" => data_out <= rom_array(15949);
		when "0011111001001110" => data_out <= rom_array(15950);
		when "0011111001001111" => data_out <= rom_array(15951);
		when "0011111001010000" => data_out <= rom_array(15952);
		when "0011111001010001" => data_out <= rom_array(15953);
		when "0011111001010010" => data_out <= rom_array(15954);
		when "0011111001010011" => data_out <= rom_array(15955);
		when "0011111001010100" => data_out <= rom_array(15956);
		when "0011111001010101" => data_out <= rom_array(15957);
		when "0011111001010110" => data_out <= rom_array(15958);
		when "0011111001010111" => data_out <= rom_array(15959);
		when "0011111001011000" => data_out <= rom_array(15960);
		when "0011111001011001" => data_out <= rom_array(15961);
		when "0011111001011010" => data_out <= rom_array(15962);
		when "0011111001011011" => data_out <= rom_array(15963);
		when "0011111001011100" => data_out <= rom_array(15964);
		when "0011111001011101" => data_out <= rom_array(15965);
		when "0011111001011110" => data_out <= rom_array(15966);
		when "0011111001011111" => data_out <= rom_array(15967);
		when "0011111001100000" => data_out <= rom_array(15968);
		when "0011111001100001" => data_out <= rom_array(15969);
		when "0011111001100010" => data_out <= rom_array(15970);
		when "0011111001100011" => data_out <= rom_array(15971);
		when "0011111001100100" => data_out <= rom_array(15972);
		when "0011111001100101" => data_out <= rom_array(15973);
		when "0011111001100110" => data_out <= rom_array(15974);
		when "0011111001100111" => data_out <= rom_array(15975);
		when "0011111001101000" => data_out <= rom_array(15976);
		when "0011111001101001" => data_out <= rom_array(15977);
		when "0011111001101010" => data_out <= rom_array(15978);
		when "0011111001101011" => data_out <= rom_array(15979);
		when "0011111001101100" => data_out <= rom_array(15980);
		when "0011111001101101" => data_out <= rom_array(15981);
		when "0011111001101110" => data_out <= rom_array(15982);
		when "0011111001101111" => data_out <= rom_array(15983);
		when "0011111001110000" => data_out <= rom_array(15984);
		when "0011111001110001" => data_out <= rom_array(15985);
		when "0011111001110010" => data_out <= rom_array(15986);
		when "0011111001110011" => data_out <= rom_array(15987);
		when "0011111001110100" => data_out <= rom_array(15988);
		when "0011111001110101" => data_out <= rom_array(15989);
		when "0011111001110110" => data_out <= rom_array(15990);
		when "0011111001110111" => data_out <= rom_array(15991);
		when "0011111001111000" => data_out <= rom_array(15992);
		when "0011111001111001" => data_out <= rom_array(15993);
		when "0011111001111010" => data_out <= rom_array(15994);
		when "0011111001111011" => data_out <= rom_array(15995);
		when "0011111001111100" => data_out <= rom_array(15996);
		when "0011111001111101" => data_out <= rom_array(15997);
		when "0011111001111110" => data_out <= rom_array(15998);
		when "0011111001111111" => data_out <= rom_array(15999);
		when "0011111010000000" => data_out <= rom_array(16000);
		when "0011111010000001" => data_out <= rom_array(16001);
		when "0011111010000010" => data_out <= rom_array(16002);
		when "0011111010000011" => data_out <= rom_array(16003);
		when "0011111010000100" => data_out <= rom_array(16004);
		when "0011111010000101" => data_out <= rom_array(16005);
		when "0011111010000110" => data_out <= rom_array(16006);
		when "0011111010000111" => data_out <= rom_array(16007);
		when "0011111010001000" => data_out <= rom_array(16008);
		when "0011111010001001" => data_out <= rom_array(16009);
		when "0011111010001010" => data_out <= rom_array(16010);
		when "0011111010001011" => data_out <= rom_array(16011);
		when "0011111010001100" => data_out <= rom_array(16012);
		when "0011111010001101" => data_out <= rom_array(16013);
		when "0011111010001110" => data_out <= rom_array(16014);
		when "0011111010001111" => data_out <= rom_array(16015);
		when "0011111010010000" => data_out <= rom_array(16016);
		when "0011111010010001" => data_out <= rom_array(16017);
		when "0011111010010010" => data_out <= rom_array(16018);
		when "0011111010010011" => data_out <= rom_array(16019);
		when "0011111010010100" => data_out <= rom_array(16020);
		when "0011111010010101" => data_out <= rom_array(16021);
		when "0011111010010110" => data_out <= rom_array(16022);
		when "0011111010010111" => data_out <= rom_array(16023);
		when "0011111010011000" => data_out <= rom_array(16024);
		when "0011111010011001" => data_out <= rom_array(16025);
		when "0011111010011010" => data_out <= rom_array(16026);
		when "0011111010011011" => data_out <= rom_array(16027);
		when "0011111010011100" => data_out <= rom_array(16028);
		when "0011111010011101" => data_out <= rom_array(16029);
		when "0011111010011110" => data_out <= rom_array(16030);
		when "0011111010011111" => data_out <= rom_array(16031);
		when "0011111010100000" => data_out <= rom_array(16032);
		when "0011111010100001" => data_out <= rom_array(16033);
		when "0011111010100010" => data_out <= rom_array(16034);
		when "0011111010100011" => data_out <= rom_array(16035);
		when "0011111010100100" => data_out <= rom_array(16036);
		when "0011111010100101" => data_out <= rom_array(16037);
		when "0011111010100110" => data_out <= rom_array(16038);
		when "0011111010100111" => data_out <= rom_array(16039);
		when "0011111010101000" => data_out <= rom_array(16040);
		when "0011111010101001" => data_out <= rom_array(16041);
		when "0011111010101010" => data_out <= rom_array(16042);
		when "0011111010101011" => data_out <= rom_array(16043);
		when "0011111010101100" => data_out <= rom_array(16044);
		when "0011111010101101" => data_out <= rom_array(16045);
		when "0011111010101110" => data_out <= rom_array(16046);
		when "0011111010101111" => data_out <= rom_array(16047);
		when "0011111010110000" => data_out <= rom_array(16048);
		when "0011111010110001" => data_out <= rom_array(16049);
		when "0011111010110010" => data_out <= rom_array(16050);
		when "0011111010110011" => data_out <= rom_array(16051);
		when "0011111010110100" => data_out <= rom_array(16052);
		when "0011111010110101" => data_out <= rom_array(16053);
		when "0011111010110110" => data_out <= rom_array(16054);
		when "0011111010110111" => data_out <= rom_array(16055);
		when "0011111010111000" => data_out <= rom_array(16056);
		when "0011111010111001" => data_out <= rom_array(16057);
		when "0011111010111010" => data_out <= rom_array(16058);
		when "0011111010111011" => data_out <= rom_array(16059);
		when "0011111010111100" => data_out <= rom_array(16060);
		when "0011111010111101" => data_out <= rom_array(16061);
		when "0011111010111110" => data_out <= rom_array(16062);
		when "0011111010111111" => data_out <= rom_array(16063);
		when "0011111011000000" => data_out <= rom_array(16064);
		when "0011111011000001" => data_out <= rom_array(16065);
		when "0011111011000010" => data_out <= rom_array(16066);
		when "0011111011000011" => data_out <= rom_array(16067);
		when "0011111011000100" => data_out <= rom_array(16068);
		when "0011111011000101" => data_out <= rom_array(16069);
		when "0011111011000110" => data_out <= rom_array(16070);
		when "0011111011000111" => data_out <= rom_array(16071);
		when "0011111011001000" => data_out <= rom_array(16072);
		when "0011111011001001" => data_out <= rom_array(16073);
		when "0011111011001010" => data_out <= rom_array(16074);
		when "0011111011001011" => data_out <= rom_array(16075);
		when "0011111011001100" => data_out <= rom_array(16076);
		when "0011111011001101" => data_out <= rom_array(16077);
		when "0011111011001110" => data_out <= rom_array(16078);
		when "0011111011001111" => data_out <= rom_array(16079);
		when "0011111011010000" => data_out <= rom_array(16080);
		when "0011111011010001" => data_out <= rom_array(16081);
		when "0011111011010010" => data_out <= rom_array(16082);
		when "0011111011010011" => data_out <= rom_array(16083);
		when "0011111011010100" => data_out <= rom_array(16084);
		when "0011111011010101" => data_out <= rom_array(16085);
		when "0011111011010110" => data_out <= rom_array(16086);
		when "0011111011010111" => data_out <= rom_array(16087);
		when "0011111011011000" => data_out <= rom_array(16088);
		when "0011111011011001" => data_out <= rom_array(16089);
		when "0011111011011010" => data_out <= rom_array(16090);
		when "0011111011011011" => data_out <= rom_array(16091);
		when "0011111011011100" => data_out <= rom_array(16092);
		when "0011111011011101" => data_out <= rom_array(16093);
		when "0011111011011110" => data_out <= rom_array(16094);
		when "0011111011011111" => data_out <= rom_array(16095);
		when "0011111011100000" => data_out <= rom_array(16096);
		when "0011111011100001" => data_out <= rom_array(16097);
		when "0011111011100010" => data_out <= rom_array(16098);
		when "0011111011100011" => data_out <= rom_array(16099);
		when "0011111011100100" => data_out <= rom_array(16100);
		when "0011111011100101" => data_out <= rom_array(16101);
		when "0011111011100110" => data_out <= rom_array(16102);
		when "0011111011100111" => data_out <= rom_array(16103);
		when "0011111011101000" => data_out <= rom_array(16104);
		when "0011111011101001" => data_out <= rom_array(16105);
		when "0011111011101010" => data_out <= rom_array(16106);
		when "0011111011101011" => data_out <= rom_array(16107);
		when "0011111011101100" => data_out <= rom_array(16108);
		when "0011111011101101" => data_out <= rom_array(16109);
		when "0011111011101110" => data_out <= rom_array(16110);
		when "0011111011101111" => data_out <= rom_array(16111);
		when "0011111011110000" => data_out <= rom_array(16112);
		when "0011111011110001" => data_out <= rom_array(16113);
		when "0011111011110010" => data_out <= rom_array(16114);
		when "0011111011110011" => data_out <= rom_array(16115);
		when "0011111011110100" => data_out <= rom_array(16116);
		when "0011111011110101" => data_out <= rom_array(16117);
		when "0011111011110110" => data_out <= rom_array(16118);
		when "0011111011110111" => data_out <= rom_array(16119);
		when "0011111011111000" => data_out <= rom_array(16120);
		when "0011111011111001" => data_out <= rom_array(16121);
		when "0011111011111010" => data_out <= rom_array(16122);
		when "0011111011111011" => data_out <= rom_array(16123);
		when "0011111011111100" => data_out <= rom_array(16124);
		when "0011111011111101" => data_out <= rom_array(16125);
		when "0011111011111110" => data_out <= rom_array(16126);
		when "0011111011111111" => data_out <= rom_array(16127);
		when "0011111100000000" => data_out <= rom_array(16128);
		when "0011111100000001" => data_out <= rom_array(16129);
		when "0011111100000010" => data_out <= rom_array(16130);
		when "0011111100000011" => data_out <= rom_array(16131);
		when "0011111100000100" => data_out <= rom_array(16132);
		when "0011111100000101" => data_out <= rom_array(16133);
		when "0011111100000110" => data_out <= rom_array(16134);
		when "0011111100000111" => data_out <= rom_array(16135);
		when "0011111100001000" => data_out <= rom_array(16136);
		when "0011111100001001" => data_out <= rom_array(16137);
		when "0011111100001010" => data_out <= rom_array(16138);
		when "0011111100001011" => data_out <= rom_array(16139);
		when "0011111100001100" => data_out <= rom_array(16140);
		when "0011111100001101" => data_out <= rom_array(16141);
		when "0011111100001110" => data_out <= rom_array(16142);
		when "0011111100001111" => data_out <= rom_array(16143);
		when "0011111100010000" => data_out <= rom_array(16144);
		when "0011111100010001" => data_out <= rom_array(16145);
		when "0011111100010010" => data_out <= rom_array(16146);
		when "0011111100010011" => data_out <= rom_array(16147);
		when "0011111100010100" => data_out <= rom_array(16148);
		when "0011111100010101" => data_out <= rom_array(16149);
		when "0011111100010110" => data_out <= rom_array(16150);
		when "0011111100010111" => data_out <= rom_array(16151);
		when "0011111100011000" => data_out <= rom_array(16152);
		when "0011111100011001" => data_out <= rom_array(16153);
		when "0011111100011010" => data_out <= rom_array(16154);
		when "0011111100011011" => data_out <= rom_array(16155);
		when "0011111100011100" => data_out <= rom_array(16156);
		when "0011111100011101" => data_out <= rom_array(16157);
		when "0011111100011110" => data_out <= rom_array(16158);
		when "0011111100011111" => data_out <= rom_array(16159);
		when "0011111100100000" => data_out <= rom_array(16160);
		when "0011111100100001" => data_out <= rom_array(16161);
		when "0011111100100010" => data_out <= rom_array(16162);
		when "0011111100100011" => data_out <= rom_array(16163);
		when "0011111100100100" => data_out <= rom_array(16164);
		when "0011111100100101" => data_out <= rom_array(16165);
		when "0011111100100110" => data_out <= rom_array(16166);
		when "0011111100100111" => data_out <= rom_array(16167);
		when "0011111100101000" => data_out <= rom_array(16168);
		when "0011111100101001" => data_out <= rom_array(16169);
		when "0011111100101010" => data_out <= rom_array(16170);
		when "0011111100101011" => data_out <= rom_array(16171);
		when "0011111100101100" => data_out <= rom_array(16172);
		when "0011111100101101" => data_out <= rom_array(16173);
		when "0011111100101110" => data_out <= rom_array(16174);
		when "0011111100101111" => data_out <= rom_array(16175);
		when "0011111100110000" => data_out <= rom_array(16176);
		when "0011111100110001" => data_out <= rom_array(16177);
		when "0011111100110010" => data_out <= rom_array(16178);
		when "0011111100110011" => data_out <= rom_array(16179);
		when "0011111100110100" => data_out <= rom_array(16180);
		when "0011111100110101" => data_out <= rom_array(16181);
		when "0011111100110110" => data_out <= rom_array(16182);
		when "0011111100110111" => data_out <= rom_array(16183);
		when "0011111100111000" => data_out <= rom_array(16184);
		when "0011111100111001" => data_out <= rom_array(16185);
		when "0011111100111010" => data_out <= rom_array(16186);
		when "0011111100111011" => data_out <= rom_array(16187);
		when "0011111100111100" => data_out <= rom_array(16188);
		when "0011111100111101" => data_out <= rom_array(16189);
		when "0011111100111110" => data_out <= rom_array(16190);
		when "0011111100111111" => data_out <= rom_array(16191);
		when "0011111101000000" => data_out <= rom_array(16192);
		when "0011111101000001" => data_out <= rom_array(16193);
		when "0011111101000010" => data_out <= rom_array(16194);
		when "0011111101000011" => data_out <= rom_array(16195);
		when "0011111101000100" => data_out <= rom_array(16196);
		when "0011111101000101" => data_out <= rom_array(16197);
		when "0011111101000110" => data_out <= rom_array(16198);
		when "0011111101000111" => data_out <= rom_array(16199);
		when "0011111101001000" => data_out <= rom_array(16200);
		when "0011111101001001" => data_out <= rom_array(16201);
		when "0011111101001010" => data_out <= rom_array(16202);
		when "0011111101001011" => data_out <= rom_array(16203);
		when "0011111101001100" => data_out <= rom_array(16204);
		when "0011111101001101" => data_out <= rom_array(16205);
		when "0011111101001110" => data_out <= rom_array(16206);
		when "0011111101001111" => data_out <= rom_array(16207);
		when "0011111101010000" => data_out <= rom_array(16208);
		when "0011111101010001" => data_out <= rom_array(16209);
		when "0011111101010010" => data_out <= rom_array(16210);
		when "0011111101010011" => data_out <= rom_array(16211);
		when "0011111101010100" => data_out <= rom_array(16212);
		when "0011111101010101" => data_out <= rom_array(16213);
		when "0011111101010110" => data_out <= rom_array(16214);
		when "0011111101010111" => data_out <= rom_array(16215);
		when "0011111101011000" => data_out <= rom_array(16216);
		when "0011111101011001" => data_out <= rom_array(16217);
		when "0011111101011010" => data_out <= rom_array(16218);
		when "0011111101011011" => data_out <= rom_array(16219);
		when "0011111101011100" => data_out <= rom_array(16220);
		when "0011111101011101" => data_out <= rom_array(16221);
		when "0011111101011110" => data_out <= rom_array(16222);
		when "0011111101011111" => data_out <= rom_array(16223);
		when "0011111101100000" => data_out <= rom_array(16224);
		when "0011111101100001" => data_out <= rom_array(16225);
		when "0011111101100010" => data_out <= rom_array(16226);
		when "0011111101100011" => data_out <= rom_array(16227);
		when "0011111101100100" => data_out <= rom_array(16228);
		when "0011111101100101" => data_out <= rom_array(16229);
		when "0011111101100110" => data_out <= rom_array(16230);
		when "0011111101100111" => data_out <= rom_array(16231);
		when "0011111101101000" => data_out <= rom_array(16232);
		when "0011111101101001" => data_out <= rom_array(16233);
		when "0011111101101010" => data_out <= rom_array(16234);
		when "0011111101101011" => data_out <= rom_array(16235);
		when "0011111101101100" => data_out <= rom_array(16236);
		when "0011111101101101" => data_out <= rom_array(16237);
		when "0011111101101110" => data_out <= rom_array(16238);
		when "0011111101101111" => data_out <= rom_array(16239);
		when "0011111101110000" => data_out <= rom_array(16240);
		when "0011111101110001" => data_out <= rom_array(16241);
		when "0011111101110010" => data_out <= rom_array(16242);
		when "0011111101110011" => data_out <= rom_array(16243);
		when "0011111101110100" => data_out <= rom_array(16244);
		when "0011111101110101" => data_out <= rom_array(16245);
		when "0011111101110110" => data_out <= rom_array(16246);
		when "0011111101110111" => data_out <= rom_array(16247);
		when "0011111101111000" => data_out <= rom_array(16248);
		when "0011111101111001" => data_out <= rom_array(16249);
		when "0011111101111010" => data_out <= rom_array(16250);
		when "0011111101111011" => data_out <= rom_array(16251);
		when "0011111101111100" => data_out <= rom_array(16252);
		when "0011111101111101" => data_out <= rom_array(16253);
		when "0011111101111110" => data_out <= rom_array(16254);
		when "0011111101111111" => data_out <= rom_array(16255);
		when "0011111110000000" => data_out <= rom_array(16256);
		when "0011111110000001" => data_out <= rom_array(16257);
		when "0011111110000010" => data_out <= rom_array(16258);
		when "0011111110000011" => data_out <= rom_array(16259);
		when "0011111110000100" => data_out <= rom_array(16260);
		when "0011111110000101" => data_out <= rom_array(16261);
		when "0011111110000110" => data_out <= rom_array(16262);
		when "0011111110000111" => data_out <= rom_array(16263);
		when "0011111110001000" => data_out <= rom_array(16264);
		when "0011111110001001" => data_out <= rom_array(16265);
		when "0011111110001010" => data_out <= rom_array(16266);
		when "0011111110001011" => data_out <= rom_array(16267);
		when "0011111110001100" => data_out <= rom_array(16268);
		when "0011111110001101" => data_out <= rom_array(16269);
		when "0011111110001110" => data_out <= rom_array(16270);
		when "0011111110001111" => data_out <= rom_array(16271);
		when "0011111110010000" => data_out <= rom_array(16272);
		when "0011111110010001" => data_out <= rom_array(16273);
		when "0011111110010010" => data_out <= rom_array(16274);
		when "0011111110010011" => data_out <= rom_array(16275);
		when "0011111110010100" => data_out <= rom_array(16276);
		when "0011111110010101" => data_out <= rom_array(16277);
		when "0011111110010110" => data_out <= rom_array(16278);
		when "0011111110010111" => data_out <= rom_array(16279);
		when "0011111110011000" => data_out <= rom_array(16280);
		when "0011111110011001" => data_out <= rom_array(16281);
		when "0011111110011010" => data_out <= rom_array(16282);
		when "0011111110011011" => data_out <= rom_array(16283);
		when "0011111110011100" => data_out <= rom_array(16284);
		when "0011111110011101" => data_out <= rom_array(16285);
		when "0011111110011110" => data_out <= rom_array(16286);
		when "0011111110011111" => data_out <= rom_array(16287);
		when "0011111110100000" => data_out <= rom_array(16288);
		when "0011111110100001" => data_out <= rom_array(16289);
		when "0011111110100010" => data_out <= rom_array(16290);
		when "0011111110100011" => data_out <= rom_array(16291);
		when "0011111110100100" => data_out <= rom_array(16292);
		when "0011111110100101" => data_out <= rom_array(16293);
		when "0011111110100110" => data_out <= rom_array(16294);
		when "0011111110100111" => data_out <= rom_array(16295);
		when "0011111110101000" => data_out <= rom_array(16296);
		when "0011111110101001" => data_out <= rom_array(16297);
		when "0011111110101010" => data_out <= rom_array(16298);
		when "0011111110101011" => data_out <= rom_array(16299);
		when "0011111110101100" => data_out <= rom_array(16300);
		when "0011111110101101" => data_out <= rom_array(16301);
		when "0011111110101110" => data_out <= rom_array(16302);
		when "0011111110101111" => data_out <= rom_array(16303);
		when "0011111110110000" => data_out <= rom_array(16304);
		when "0011111110110001" => data_out <= rom_array(16305);
		when "0011111110110010" => data_out <= rom_array(16306);
		when "0011111110110011" => data_out <= rom_array(16307);
		when "0011111110110100" => data_out <= rom_array(16308);
		when "0011111110110101" => data_out <= rom_array(16309);
		when "0011111110110110" => data_out <= rom_array(16310);
		when "0011111110110111" => data_out <= rom_array(16311);
		when "0011111110111000" => data_out <= rom_array(16312);
		when "0011111110111001" => data_out <= rom_array(16313);
		when "0011111110111010" => data_out <= rom_array(16314);
		when "0011111110111011" => data_out <= rom_array(16315);
		when "0011111110111100" => data_out <= rom_array(16316);
		when "0011111110111101" => data_out <= rom_array(16317);
		when "0011111110111110" => data_out <= rom_array(16318);
		when "0011111110111111" => data_out <= rom_array(16319);
		when "0011111111000000" => data_out <= rom_array(16320);
		when "0011111111000001" => data_out <= rom_array(16321);
		when "0011111111000010" => data_out <= rom_array(16322);
		when "0011111111000011" => data_out <= rom_array(16323);
		when "0011111111000100" => data_out <= rom_array(16324);
		when "0011111111000101" => data_out <= rom_array(16325);
		when "0011111111000110" => data_out <= rom_array(16326);
		when "0011111111000111" => data_out <= rom_array(16327);
		when "0011111111001000" => data_out <= rom_array(16328);
		when "0011111111001001" => data_out <= rom_array(16329);
		when "0011111111001010" => data_out <= rom_array(16330);
		when "0011111111001011" => data_out <= rom_array(16331);
		when "0011111111001100" => data_out <= rom_array(16332);
		when "0011111111001101" => data_out <= rom_array(16333);
		when "0011111111001110" => data_out <= rom_array(16334);
		when "0011111111001111" => data_out <= rom_array(16335);
		when "0011111111010000" => data_out <= rom_array(16336);
		when "0011111111010001" => data_out <= rom_array(16337);
		when "0011111111010010" => data_out <= rom_array(16338);
		when "0011111111010011" => data_out <= rom_array(16339);
		when "0011111111010100" => data_out <= rom_array(16340);
		when "0011111111010101" => data_out <= rom_array(16341);
		when "0011111111010110" => data_out <= rom_array(16342);
		when "0011111111010111" => data_out <= rom_array(16343);
		when "0011111111011000" => data_out <= rom_array(16344);
		when "0011111111011001" => data_out <= rom_array(16345);
		when "0011111111011010" => data_out <= rom_array(16346);
		when "0011111111011011" => data_out <= rom_array(16347);
		when "0011111111011100" => data_out <= rom_array(16348);
		when "0011111111011101" => data_out <= rom_array(16349);
		when "0011111111011110" => data_out <= rom_array(16350);
		when "0011111111011111" => data_out <= rom_array(16351);
		when "0011111111100000" => data_out <= rom_array(16352);
		when "0011111111100001" => data_out <= rom_array(16353);
		when "0011111111100010" => data_out <= rom_array(16354);
		when "0011111111100011" => data_out <= rom_array(16355);
		when "0011111111100100" => data_out <= rom_array(16356);
		when "0011111111100101" => data_out <= rom_array(16357);
		when "0011111111100110" => data_out <= rom_array(16358);
		when "0011111111100111" => data_out <= rom_array(16359);
		when "0011111111101000" => data_out <= rom_array(16360);
		when "0011111111101001" => data_out <= rom_array(16361);
		when "0011111111101010" => data_out <= rom_array(16362);
		when "0011111111101011" => data_out <= rom_array(16363);
		when "0011111111101100" => data_out <= rom_array(16364);
		when "0011111111101101" => data_out <= rom_array(16365);
		when "0011111111101110" => data_out <= rom_array(16366);
		when "0011111111101111" => data_out <= rom_array(16367);
		when "0011111111110000" => data_out <= rom_array(16368);
		when "0011111111110001" => data_out <= rom_array(16369);
		when "0011111111110010" => data_out <= rom_array(16370);
		when "0011111111110011" => data_out <= rom_array(16371);
		when "0011111111110100" => data_out <= rom_array(16372);
		when "0011111111110101" => data_out <= rom_array(16373);
		when "0011111111110110" => data_out <= rom_array(16374);
		when "0011111111110111" => data_out <= rom_array(16375);
		when "0011111111111000" => data_out <= rom_array(16376);
		when "0011111111111001" => data_out <= rom_array(16377);
		when "0011111111111010" => data_out <= rom_array(16378);
		when "0011111111111011" => data_out <= rom_array(16379);
		when "0011111111111100" => data_out <= rom_array(16380);
		when "0011111111111101" => data_out <= rom_array(16381);
		when "0011111111111110" => data_out <= rom_array(16382);
		when "0011111111111111" => data_out <= rom_array(16383);
		when "0100000000000000" => data_out <= rom_array(16384);
		when "0100000000000001" => data_out <= rom_array(16385);
		when "0100000000000010" => data_out <= rom_array(16386);
		when "0100000000000011" => data_out <= rom_array(16387);
		when "0100000000000100" => data_out <= rom_array(16388);
		when "0100000000000101" => data_out <= rom_array(16389);
		when "0100000000000110" => data_out <= rom_array(16390);
		when "0100000000000111" => data_out <= rom_array(16391);
		when "0100000000001000" => data_out <= rom_array(16392);
		when "0100000000001001" => data_out <= rom_array(16393);
		when "0100000000001010" => data_out <= rom_array(16394);
		when "0100000000001011" => data_out <= rom_array(16395);
		when "0100000000001100" => data_out <= rom_array(16396);
		when "0100000000001101" => data_out <= rom_array(16397);
		when "0100000000001110" => data_out <= rom_array(16398);
		when "0100000000001111" => data_out <= rom_array(16399);
		when "0100000000010000" => data_out <= rom_array(16400);
		when "0100000000010001" => data_out <= rom_array(16401);
		when "0100000000010010" => data_out <= rom_array(16402);
		when "0100000000010011" => data_out <= rom_array(16403);
		when "0100000000010100" => data_out <= rom_array(16404);
		when "0100000000010101" => data_out <= rom_array(16405);
		when "0100000000010110" => data_out <= rom_array(16406);
		when "0100000000010111" => data_out <= rom_array(16407);
		when "0100000000011000" => data_out <= rom_array(16408);
		when "0100000000011001" => data_out <= rom_array(16409);
		when "0100000000011010" => data_out <= rom_array(16410);
		when "0100000000011011" => data_out <= rom_array(16411);
		when "0100000000011100" => data_out <= rom_array(16412);
		when "0100000000011101" => data_out <= rom_array(16413);
		when "0100000000011110" => data_out <= rom_array(16414);
		when "0100000000011111" => data_out <= rom_array(16415);
		when "0100000000100000" => data_out <= rom_array(16416);
		when "0100000000100001" => data_out <= rom_array(16417);
		when "0100000000100010" => data_out <= rom_array(16418);
		when "0100000000100011" => data_out <= rom_array(16419);
		when "0100000000100100" => data_out <= rom_array(16420);
		when "0100000000100101" => data_out <= rom_array(16421);
		when "0100000000100110" => data_out <= rom_array(16422);
		when "0100000000100111" => data_out <= rom_array(16423);
		when "0100000000101000" => data_out <= rom_array(16424);
		when "0100000000101001" => data_out <= rom_array(16425);
		when "0100000000101010" => data_out <= rom_array(16426);
		when "0100000000101011" => data_out <= rom_array(16427);
		when "0100000000101100" => data_out <= rom_array(16428);
		when "0100000000101101" => data_out <= rom_array(16429);
		when "0100000000101110" => data_out <= rom_array(16430);
		when "0100000000101111" => data_out <= rom_array(16431);
		when "0100000000110000" => data_out <= rom_array(16432);
		when "0100000000110001" => data_out <= rom_array(16433);
		when "0100000000110010" => data_out <= rom_array(16434);
		when "0100000000110011" => data_out <= rom_array(16435);
		when "0100000000110100" => data_out <= rom_array(16436);
		when "0100000000110101" => data_out <= rom_array(16437);
		when "0100000000110110" => data_out <= rom_array(16438);
		when "0100000000110111" => data_out <= rom_array(16439);
		when "0100000000111000" => data_out <= rom_array(16440);
		when "0100000000111001" => data_out <= rom_array(16441);
		when "0100000000111010" => data_out <= rom_array(16442);
		when "0100000000111011" => data_out <= rom_array(16443);
		when "0100000000111100" => data_out <= rom_array(16444);
		when "0100000000111101" => data_out <= rom_array(16445);
		when "0100000000111110" => data_out <= rom_array(16446);
		when "0100000000111111" => data_out <= rom_array(16447);
		when "0100000001000000" => data_out <= rom_array(16448);
		when "0100000001000001" => data_out <= rom_array(16449);
		when "0100000001000010" => data_out <= rom_array(16450);
		when "0100000001000011" => data_out <= rom_array(16451);
		when "0100000001000100" => data_out <= rom_array(16452);
		when "0100000001000101" => data_out <= rom_array(16453);
		when "0100000001000110" => data_out <= rom_array(16454);
		when "0100000001000111" => data_out <= rom_array(16455);
		when "0100000001001000" => data_out <= rom_array(16456);
		when "0100000001001001" => data_out <= rom_array(16457);
		when "0100000001001010" => data_out <= rom_array(16458);
		when "0100000001001011" => data_out <= rom_array(16459);
		when "0100000001001100" => data_out <= rom_array(16460);
		when "0100000001001101" => data_out <= rom_array(16461);
		when "0100000001001110" => data_out <= rom_array(16462);
		when "0100000001001111" => data_out <= rom_array(16463);
		when "0100000001010000" => data_out <= rom_array(16464);
		when "0100000001010001" => data_out <= rom_array(16465);
		when "0100000001010010" => data_out <= rom_array(16466);
		when "0100000001010011" => data_out <= rom_array(16467);
		when "0100000001010100" => data_out <= rom_array(16468);
		when "0100000001010101" => data_out <= rom_array(16469);
		when "0100000001010110" => data_out <= rom_array(16470);
		when "0100000001010111" => data_out <= rom_array(16471);
		when "0100000001011000" => data_out <= rom_array(16472);
		when "0100000001011001" => data_out <= rom_array(16473);
		when "0100000001011010" => data_out <= rom_array(16474);
		when "0100000001011011" => data_out <= rom_array(16475);
		when "0100000001011100" => data_out <= rom_array(16476);
		when "0100000001011101" => data_out <= rom_array(16477);
		when "0100000001011110" => data_out <= rom_array(16478);
		when "0100000001011111" => data_out <= rom_array(16479);
		when "0100000001100000" => data_out <= rom_array(16480);
		when "0100000001100001" => data_out <= rom_array(16481);
		when "0100000001100010" => data_out <= rom_array(16482);
		when "0100000001100011" => data_out <= rom_array(16483);
		when "0100000001100100" => data_out <= rom_array(16484);
		when "0100000001100101" => data_out <= rom_array(16485);
		when "0100000001100110" => data_out <= rom_array(16486);
		when "0100000001100111" => data_out <= rom_array(16487);
		when "0100000001101000" => data_out <= rom_array(16488);
		when "0100000001101001" => data_out <= rom_array(16489);
		when "0100000001101010" => data_out <= rom_array(16490);
		when "0100000001101011" => data_out <= rom_array(16491);
		when "0100000001101100" => data_out <= rom_array(16492);
		when "0100000001101101" => data_out <= rom_array(16493);
		when "0100000001101110" => data_out <= rom_array(16494);
		when "0100000001101111" => data_out <= rom_array(16495);
		when "0100000001110000" => data_out <= rom_array(16496);
		when "0100000001110001" => data_out <= rom_array(16497);
		when "0100000001110010" => data_out <= rom_array(16498);
		when "0100000001110011" => data_out <= rom_array(16499);
		when "0100000001110100" => data_out <= rom_array(16500);
		when "0100000001110101" => data_out <= rom_array(16501);
		when "0100000001110110" => data_out <= rom_array(16502);
		when "0100000001110111" => data_out <= rom_array(16503);
		when "0100000001111000" => data_out <= rom_array(16504);
		when "0100000001111001" => data_out <= rom_array(16505);
		when "0100000001111010" => data_out <= rom_array(16506);
		when "0100000001111011" => data_out <= rom_array(16507);
		when "0100000001111100" => data_out <= rom_array(16508);
		when "0100000001111101" => data_out <= rom_array(16509);
		when "0100000001111110" => data_out <= rom_array(16510);
		when "0100000001111111" => data_out <= rom_array(16511);
		when "0100000010000000" => data_out <= rom_array(16512);
		when "0100000010000001" => data_out <= rom_array(16513);
		when "0100000010000010" => data_out <= rom_array(16514);
		when "0100000010000011" => data_out <= rom_array(16515);
		when "0100000010000100" => data_out <= rom_array(16516);
		when "0100000010000101" => data_out <= rom_array(16517);
		when "0100000010000110" => data_out <= rom_array(16518);
		when "0100000010000111" => data_out <= rom_array(16519);
		when "0100000010001000" => data_out <= rom_array(16520);
		when "0100000010001001" => data_out <= rom_array(16521);
		when "0100000010001010" => data_out <= rom_array(16522);
		when "0100000010001011" => data_out <= rom_array(16523);
		when "0100000010001100" => data_out <= rom_array(16524);
		when "0100000010001101" => data_out <= rom_array(16525);
		when "0100000010001110" => data_out <= rom_array(16526);
		when "0100000010001111" => data_out <= rom_array(16527);
		when "0100000010010000" => data_out <= rom_array(16528);
		when "0100000010010001" => data_out <= rom_array(16529);
		when "0100000010010010" => data_out <= rom_array(16530);
		when "0100000010010011" => data_out <= rom_array(16531);
		when "0100000010010100" => data_out <= rom_array(16532);
		when "0100000010010101" => data_out <= rom_array(16533);
		when "0100000010010110" => data_out <= rom_array(16534);
		when "0100000010010111" => data_out <= rom_array(16535);
		when "0100000010011000" => data_out <= rom_array(16536);
		when "0100000010011001" => data_out <= rom_array(16537);
		when "0100000010011010" => data_out <= rom_array(16538);
		when "0100000010011011" => data_out <= rom_array(16539);
		when "0100000010011100" => data_out <= rom_array(16540);
		when "0100000010011101" => data_out <= rom_array(16541);
		when "0100000010011110" => data_out <= rom_array(16542);
		when "0100000010011111" => data_out <= rom_array(16543);
		when "0100000010100000" => data_out <= rom_array(16544);
		when "0100000010100001" => data_out <= rom_array(16545);
		when "0100000010100010" => data_out <= rom_array(16546);
		when "0100000010100011" => data_out <= rom_array(16547);
		when "0100000010100100" => data_out <= rom_array(16548);
		when "0100000010100101" => data_out <= rom_array(16549);
		when "0100000010100110" => data_out <= rom_array(16550);
		when "0100000010100111" => data_out <= rom_array(16551);
		when "0100000010101000" => data_out <= rom_array(16552);
		when "0100000010101001" => data_out <= rom_array(16553);
		when "0100000010101010" => data_out <= rom_array(16554);
		when "0100000010101011" => data_out <= rom_array(16555);
		when "0100000010101100" => data_out <= rom_array(16556);
		when "0100000010101101" => data_out <= rom_array(16557);
		when "0100000010101110" => data_out <= rom_array(16558);
		when "0100000010101111" => data_out <= rom_array(16559);
		when "0100000010110000" => data_out <= rom_array(16560);
		when "0100000010110001" => data_out <= rom_array(16561);
		when "0100000010110010" => data_out <= rom_array(16562);
		when "0100000010110011" => data_out <= rom_array(16563);
		when "0100000010110100" => data_out <= rom_array(16564);
		when "0100000010110101" => data_out <= rom_array(16565);
		when "0100000010110110" => data_out <= rom_array(16566);
		when "0100000010110111" => data_out <= rom_array(16567);
		when "0100000010111000" => data_out <= rom_array(16568);
		when "0100000010111001" => data_out <= rom_array(16569);
		when "0100000010111010" => data_out <= rom_array(16570);
		when "0100000010111011" => data_out <= rom_array(16571);
		when "0100000010111100" => data_out <= rom_array(16572);
		when "0100000010111101" => data_out <= rom_array(16573);
		when "0100000010111110" => data_out <= rom_array(16574);
		when "0100000010111111" => data_out <= rom_array(16575);
		when "0100000011000000" => data_out <= rom_array(16576);
		when "0100000011000001" => data_out <= rom_array(16577);
		when "0100000011000010" => data_out <= rom_array(16578);
		when "0100000011000011" => data_out <= rom_array(16579);
		when "0100000011000100" => data_out <= rom_array(16580);
		when "0100000011000101" => data_out <= rom_array(16581);
		when "0100000011000110" => data_out <= rom_array(16582);
		when "0100000011000111" => data_out <= rom_array(16583);
		when "0100000011001000" => data_out <= rom_array(16584);
		when "0100000011001001" => data_out <= rom_array(16585);
		when "0100000011001010" => data_out <= rom_array(16586);
		when "0100000011001011" => data_out <= rom_array(16587);
		when "0100000011001100" => data_out <= rom_array(16588);
		when "0100000011001101" => data_out <= rom_array(16589);
		when "0100000011001110" => data_out <= rom_array(16590);
		when "0100000011001111" => data_out <= rom_array(16591);
		when "0100000011010000" => data_out <= rom_array(16592);
		when "0100000011010001" => data_out <= rom_array(16593);
		when "0100000011010010" => data_out <= rom_array(16594);
		when "0100000011010011" => data_out <= rom_array(16595);
		when "0100000011010100" => data_out <= rom_array(16596);
		when "0100000011010101" => data_out <= rom_array(16597);
		when "0100000011010110" => data_out <= rom_array(16598);
		when "0100000011010111" => data_out <= rom_array(16599);
		when "0100000011011000" => data_out <= rom_array(16600);
		when "0100000011011001" => data_out <= rom_array(16601);
		when "0100000011011010" => data_out <= rom_array(16602);
		when "0100000011011011" => data_out <= rom_array(16603);
		when "0100000011011100" => data_out <= rom_array(16604);
		when "0100000011011101" => data_out <= rom_array(16605);
		when "0100000011011110" => data_out <= rom_array(16606);
		when "0100000011011111" => data_out <= rom_array(16607);
		when "0100000011100000" => data_out <= rom_array(16608);
		when "0100000011100001" => data_out <= rom_array(16609);
		when "0100000011100010" => data_out <= rom_array(16610);
		when "0100000011100011" => data_out <= rom_array(16611);
		when "0100000011100100" => data_out <= rom_array(16612);
		when "0100000011100101" => data_out <= rom_array(16613);
		when "0100000011100110" => data_out <= rom_array(16614);
		when "0100000011100111" => data_out <= rom_array(16615);
		when "0100000011101000" => data_out <= rom_array(16616);
		when "0100000011101001" => data_out <= rom_array(16617);
		when "0100000011101010" => data_out <= rom_array(16618);
		when "0100000011101011" => data_out <= rom_array(16619);
		when "0100000011101100" => data_out <= rom_array(16620);
		when "0100000011101101" => data_out <= rom_array(16621);
		when "0100000011101110" => data_out <= rom_array(16622);
		when "0100000011101111" => data_out <= rom_array(16623);
		when "0100000011110000" => data_out <= rom_array(16624);
		when "0100000011110001" => data_out <= rom_array(16625);
		when "0100000011110010" => data_out <= rom_array(16626);
		when "0100000011110011" => data_out <= rom_array(16627);
		when "0100000011110100" => data_out <= rom_array(16628);
		when "0100000011110101" => data_out <= rom_array(16629);
		when "0100000011110110" => data_out <= rom_array(16630);
		when "0100000011110111" => data_out <= rom_array(16631);
		when "0100000011111000" => data_out <= rom_array(16632);
		when "0100000011111001" => data_out <= rom_array(16633);
		when "0100000011111010" => data_out <= rom_array(16634);
		when "0100000011111011" => data_out <= rom_array(16635);
		when "0100000011111100" => data_out <= rom_array(16636);
		when "0100000011111101" => data_out <= rom_array(16637);
		when "0100000011111110" => data_out <= rom_array(16638);
		when "0100000011111111" => data_out <= rom_array(16639);
		when "0100000100000000" => data_out <= rom_array(16640);
		when "0100000100000001" => data_out <= rom_array(16641);
		when "0100000100000010" => data_out <= rom_array(16642);
		when "0100000100000011" => data_out <= rom_array(16643);
		when "0100000100000100" => data_out <= rom_array(16644);
		when "0100000100000101" => data_out <= rom_array(16645);
		when "0100000100000110" => data_out <= rom_array(16646);
		when "0100000100000111" => data_out <= rom_array(16647);
		when "0100000100001000" => data_out <= rom_array(16648);
		when "0100000100001001" => data_out <= rom_array(16649);
		when "0100000100001010" => data_out <= rom_array(16650);
		when "0100000100001011" => data_out <= rom_array(16651);
		when "0100000100001100" => data_out <= rom_array(16652);
		when "0100000100001101" => data_out <= rom_array(16653);
		when "0100000100001110" => data_out <= rom_array(16654);
		when "0100000100001111" => data_out <= rom_array(16655);
		when "0100000100010000" => data_out <= rom_array(16656);
		when "0100000100010001" => data_out <= rom_array(16657);
		when "0100000100010010" => data_out <= rom_array(16658);
		when "0100000100010011" => data_out <= rom_array(16659);
		when "0100000100010100" => data_out <= rom_array(16660);
		when "0100000100010101" => data_out <= rom_array(16661);
		when "0100000100010110" => data_out <= rom_array(16662);
		when "0100000100010111" => data_out <= rom_array(16663);
		when "0100000100011000" => data_out <= rom_array(16664);
		when "0100000100011001" => data_out <= rom_array(16665);
		when "0100000100011010" => data_out <= rom_array(16666);
		when "0100000100011011" => data_out <= rom_array(16667);
		when "0100000100011100" => data_out <= rom_array(16668);
		when "0100000100011101" => data_out <= rom_array(16669);
		when "0100000100011110" => data_out <= rom_array(16670);
		when "0100000100011111" => data_out <= rom_array(16671);
		when "0100000100100000" => data_out <= rom_array(16672);
		when "0100000100100001" => data_out <= rom_array(16673);
		when "0100000100100010" => data_out <= rom_array(16674);
		when "0100000100100011" => data_out <= rom_array(16675);
		when "0100000100100100" => data_out <= rom_array(16676);
		when "0100000100100101" => data_out <= rom_array(16677);
		when "0100000100100110" => data_out <= rom_array(16678);
		when "0100000100100111" => data_out <= rom_array(16679);
		when "0100000100101000" => data_out <= rom_array(16680);
		when "0100000100101001" => data_out <= rom_array(16681);
		when "0100000100101010" => data_out <= rom_array(16682);
		when "0100000100101011" => data_out <= rom_array(16683);
		when "0100000100101100" => data_out <= rom_array(16684);
		when "0100000100101101" => data_out <= rom_array(16685);
		when "0100000100101110" => data_out <= rom_array(16686);
		when "0100000100101111" => data_out <= rom_array(16687);
		when "0100000100110000" => data_out <= rom_array(16688);
		when "0100000100110001" => data_out <= rom_array(16689);
		when "0100000100110010" => data_out <= rom_array(16690);
		when "0100000100110011" => data_out <= rom_array(16691);
		when "0100000100110100" => data_out <= rom_array(16692);
		when "0100000100110101" => data_out <= rom_array(16693);
		when "0100000100110110" => data_out <= rom_array(16694);
		when "0100000100110111" => data_out <= rom_array(16695);
		when "0100000100111000" => data_out <= rom_array(16696);
		when "0100000100111001" => data_out <= rom_array(16697);
		when "0100000100111010" => data_out <= rom_array(16698);
		when "0100000100111011" => data_out <= rom_array(16699);
		when "0100000100111100" => data_out <= rom_array(16700);
		when "0100000100111101" => data_out <= rom_array(16701);
		when "0100000100111110" => data_out <= rom_array(16702);
		when "0100000100111111" => data_out <= rom_array(16703);
		when "0100000101000000" => data_out <= rom_array(16704);
		when "0100000101000001" => data_out <= rom_array(16705);
		when "0100000101000010" => data_out <= rom_array(16706);
		when "0100000101000011" => data_out <= rom_array(16707);
		when "0100000101000100" => data_out <= rom_array(16708);
		when "0100000101000101" => data_out <= rom_array(16709);
		when "0100000101000110" => data_out <= rom_array(16710);
		when "0100000101000111" => data_out <= rom_array(16711);
		when "0100000101001000" => data_out <= rom_array(16712);
		when "0100000101001001" => data_out <= rom_array(16713);
		when "0100000101001010" => data_out <= rom_array(16714);
		when "0100000101001011" => data_out <= rom_array(16715);
		when "0100000101001100" => data_out <= rom_array(16716);
		when "0100000101001101" => data_out <= rom_array(16717);
		when "0100000101001110" => data_out <= rom_array(16718);
		when "0100000101001111" => data_out <= rom_array(16719);
		when "0100000101010000" => data_out <= rom_array(16720);
		when "0100000101010001" => data_out <= rom_array(16721);
		when "0100000101010010" => data_out <= rom_array(16722);
		when "0100000101010011" => data_out <= rom_array(16723);
		when "0100000101010100" => data_out <= rom_array(16724);
		when "0100000101010101" => data_out <= rom_array(16725);
		when "0100000101010110" => data_out <= rom_array(16726);
		when "0100000101010111" => data_out <= rom_array(16727);
		when "0100000101011000" => data_out <= rom_array(16728);
		when "0100000101011001" => data_out <= rom_array(16729);
		when "0100000101011010" => data_out <= rom_array(16730);
		when "0100000101011011" => data_out <= rom_array(16731);
		when "0100000101011100" => data_out <= rom_array(16732);
		when "0100000101011101" => data_out <= rom_array(16733);
		when "0100000101011110" => data_out <= rom_array(16734);
		when "0100000101011111" => data_out <= rom_array(16735);
		when "0100000101100000" => data_out <= rom_array(16736);
		when "0100000101100001" => data_out <= rom_array(16737);
		when "0100000101100010" => data_out <= rom_array(16738);
		when "0100000101100011" => data_out <= rom_array(16739);
		when "0100000101100100" => data_out <= rom_array(16740);
		when "0100000101100101" => data_out <= rom_array(16741);
		when "0100000101100110" => data_out <= rom_array(16742);
		when "0100000101100111" => data_out <= rom_array(16743);
		when "0100000101101000" => data_out <= rom_array(16744);
		when "0100000101101001" => data_out <= rom_array(16745);
		when "0100000101101010" => data_out <= rom_array(16746);
		when "0100000101101011" => data_out <= rom_array(16747);
		when "0100000101101100" => data_out <= rom_array(16748);
		when "0100000101101101" => data_out <= rom_array(16749);
		when "0100000101101110" => data_out <= rom_array(16750);
		when "0100000101101111" => data_out <= rom_array(16751);
		when "0100000101110000" => data_out <= rom_array(16752);
		when "0100000101110001" => data_out <= rom_array(16753);
		when "0100000101110010" => data_out <= rom_array(16754);
		when "0100000101110011" => data_out <= rom_array(16755);
		when "0100000101110100" => data_out <= rom_array(16756);
		when "0100000101110101" => data_out <= rom_array(16757);
		when "0100000101110110" => data_out <= rom_array(16758);
		when "0100000101110111" => data_out <= rom_array(16759);
		when "0100000101111000" => data_out <= rom_array(16760);
		when "0100000101111001" => data_out <= rom_array(16761);
		when "0100000101111010" => data_out <= rom_array(16762);
		when "0100000101111011" => data_out <= rom_array(16763);
		when "0100000101111100" => data_out <= rom_array(16764);
		when "0100000101111101" => data_out <= rom_array(16765);
		when "0100000101111110" => data_out <= rom_array(16766);
		when "0100000101111111" => data_out <= rom_array(16767);
		when "0100000110000000" => data_out <= rom_array(16768);
		when "0100000110000001" => data_out <= rom_array(16769);
		when "0100000110000010" => data_out <= rom_array(16770);
		when "0100000110000011" => data_out <= rom_array(16771);
		when "0100000110000100" => data_out <= rom_array(16772);
		when "0100000110000101" => data_out <= rom_array(16773);
		when "0100000110000110" => data_out <= rom_array(16774);
		when "0100000110000111" => data_out <= rom_array(16775);
		when "0100000110001000" => data_out <= rom_array(16776);
		when "0100000110001001" => data_out <= rom_array(16777);
		when "0100000110001010" => data_out <= rom_array(16778);
		when "0100000110001011" => data_out <= rom_array(16779);
		when "0100000110001100" => data_out <= rom_array(16780);
		when "0100000110001101" => data_out <= rom_array(16781);
		when "0100000110001110" => data_out <= rom_array(16782);
		when "0100000110001111" => data_out <= rom_array(16783);
		when "0100000110010000" => data_out <= rom_array(16784);
		when "0100000110010001" => data_out <= rom_array(16785);
		when "0100000110010010" => data_out <= rom_array(16786);
		when "0100000110010011" => data_out <= rom_array(16787);
		when "0100000110010100" => data_out <= rom_array(16788);
		when "0100000110010101" => data_out <= rom_array(16789);
		when "0100000110010110" => data_out <= rom_array(16790);
		when "0100000110010111" => data_out <= rom_array(16791);
		when "0100000110011000" => data_out <= rom_array(16792);
		when "0100000110011001" => data_out <= rom_array(16793);
		when "0100000110011010" => data_out <= rom_array(16794);
		when "0100000110011011" => data_out <= rom_array(16795);
		when "0100000110011100" => data_out <= rom_array(16796);
		when "0100000110011101" => data_out <= rom_array(16797);
		when "0100000110011110" => data_out <= rom_array(16798);
		when "0100000110011111" => data_out <= rom_array(16799);
		when "0100000110100000" => data_out <= rom_array(16800);
		when "0100000110100001" => data_out <= rom_array(16801);
		when "0100000110100010" => data_out <= rom_array(16802);
		when "0100000110100011" => data_out <= rom_array(16803);
		when "0100000110100100" => data_out <= rom_array(16804);
		when "0100000110100101" => data_out <= rom_array(16805);
		when "0100000110100110" => data_out <= rom_array(16806);
		when "0100000110100111" => data_out <= rom_array(16807);
		when "0100000110101000" => data_out <= rom_array(16808);
		when "0100000110101001" => data_out <= rom_array(16809);
		when "0100000110101010" => data_out <= rom_array(16810);
		when "0100000110101011" => data_out <= rom_array(16811);
		when "0100000110101100" => data_out <= rom_array(16812);
		when "0100000110101101" => data_out <= rom_array(16813);
		when "0100000110101110" => data_out <= rom_array(16814);
		when "0100000110101111" => data_out <= rom_array(16815);
		when "0100000110110000" => data_out <= rom_array(16816);
		when "0100000110110001" => data_out <= rom_array(16817);
		when "0100000110110010" => data_out <= rom_array(16818);
		when "0100000110110011" => data_out <= rom_array(16819);
		when "0100000110110100" => data_out <= rom_array(16820);
		when "0100000110110101" => data_out <= rom_array(16821);
		when "0100000110110110" => data_out <= rom_array(16822);
		when "0100000110110111" => data_out <= rom_array(16823);
		when "0100000110111000" => data_out <= rom_array(16824);
		when "0100000110111001" => data_out <= rom_array(16825);
		when "0100000110111010" => data_out <= rom_array(16826);
		when "0100000110111011" => data_out <= rom_array(16827);
		when "0100000110111100" => data_out <= rom_array(16828);
		when "0100000110111101" => data_out <= rom_array(16829);
		when "0100000110111110" => data_out <= rom_array(16830);
		when "0100000110111111" => data_out <= rom_array(16831);
		when "0100000111000000" => data_out <= rom_array(16832);
		when "0100000111000001" => data_out <= rom_array(16833);
		when "0100000111000010" => data_out <= rom_array(16834);
		when "0100000111000011" => data_out <= rom_array(16835);
		when "0100000111000100" => data_out <= rom_array(16836);
		when "0100000111000101" => data_out <= rom_array(16837);
		when "0100000111000110" => data_out <= rom_array(16838);
		when "0100000111000111" => data_out <= rom_array(16839);
		when "0100000111001000" => data_out <= rom_array(16840);
		when "0100000111001001" => data_out <= rom_array(16841);
		when "0100000111001010" => data_out <= rom_array(16842);
		when "0100000111001011" => data_out <= rom_array(16843);
		when "0100000111001100" => data_out <= rom_array(16844);
		when "0100000111001101" => data_out <= rom_array(16845);
		when "0100000111001110" => data_out <= rom_array(16846);
		when "0100000111001111" => data_out <= rom_array(16847);
		when "0100000111010000" => data_out <= rom_array(16848);
		when "0100000111010001" => data_out <= rom_array(16849);
		when "0100000111010010" => data_out <= rom_array(16850);
		when "0100000111010011" => data_out <= rom_array(16851);
		when "0100000111010100" => data_out <= rom_array(16852);
		when "0100000111010101" => data_out <= rom_array(16853);
		when "0100000111010110" => data_out <= rom_array(16854);
		when "0100000111010111" => data_out <= rom_array(16855);
		when "0100000111011000" => data_out <= rom_array(16856);
		when "0100000111011001" => data_out <= rom_array(16857);
		when "0100000111011010" => data_out <= rom_array(16858);
		when "0100000111011011" => data_out <= rom_array(16859);
		when "0100000111011100" => data_out <= rom_array(16860);
		when "0100000111011101" => data_out <= rom_array(16861);
		when "0100000111011110" => data_out <= rom_array(16862);
		when "0100000111011111" => data_out <= rom_array(16863);
		when "0100000111100000" => data_out <= rom_array(16864);
		when "0100000111100001" => data_out <= rom_array(16865);
		when "0100000111100010" => data_out <= rom_array(16866);
		when "0100000111100011" => data_out <= rom_array(16867);
		when "0100000111100100" => data_out <= rom_array(16868);
		when "0100000111100101" => data_out <= rom_array(16869);
		when "0100000111100110" => data_out <= rom_array(16870);
		when "0100000111100111" => data_out <= rom_array(16871);
		when "0100000111101000" => data_out <= rom_array(16872);
		when "0100000111101001" => data_out <= rom_array(16873);
		when "0100000111101010" => data_out <= rom_array(16874);
		when "0100000111101011" => data_out <= rom_array(16875);
		when "0100000111101100" => data_out <= rom_array(16876);
		when "0100000111101101" => data_out <= rom_array(16877);
		when "0100000111101110" => data_out <= rom_array(16878);
		when "0100000111101111" => data_out <= rom_array(16879);
		when "0100000111110000" => data_out <= rom_array(16880);
		when "0100000111110001" => data_out <= rom_array(16881);
		when "0100000111110010" => data_out <= rom_array(16882);
		when "0100000111110011" => data_out <= rom_array(16883);
		when "0100000111110100" => data_out <= rom_array(16884);
		when "0100000111110101" => data_out <= rom_array(16885);
		when "0100000111110110" => data_out <= rom_array(16886);
		when "0100000111110111" => data_out <= rom_array(16887);
		when "0100000111111000" => data_out <= rom_array(16888);
		when "0100000111111001" => data_out <= rom_array(16889);
		when "0100000111111010" => data_out <= rom_array(16890);
		when "0100000111111011" => data_out <= rom_array(16891);
		when "0100000111111100" => data_out <= rom_array(16892);
		when "0100000111111101" => data_out <= rom_array(16893);
		when "0100000111111110" => data_out <= rom_array(16894);
		when "0100000111111111" => data_out <= rom_array(16895);
		when "0100001000000000" => data_out <= rom_array(16896);
		when "0100001000000001" => data_out <= rom_array(16897);
		when "0100001000000010" => data_out <= rom_array(16898);
		when "0100001000000011" => data_out <= rom_array(16899);
		when "0100001000000100" => data_out <= rom_array(16900);
		when "0100001000000101" => data_out <= rom_array(16901);
		when "0100001000000110" => data_out <= rom_array(16902);
		when "0100001000000111" => data_out <= rom_array(16903);
		when "0100001000001000" => data_out <= rom_array(16904);
		when "0100001000001001" => data_out <= rom_array(16905);
		when "0100001000001010" => data_out <= rom_array(16906);
		when "0100001000001011" => data_out <= rom_array(16907);
		when "0100001000001100" => data_out <= rom_array(16908);
		when "0100001000001101" => data_out <= rom_array(16909);
		when "0100001000001110" => data_out <= rom_array(16910);
		when "0100001000001111" => data_out <= rom_array(16911);
		when "0100001000010000" => data_out <= rom_array(16912);
		when "0100001000010001" => data_out <= rom_array(16913);
		when "0100001000010010" => data_out <= rom_array(16914);
		when "0100001000010011" => data_out <= rom_array(16915);
		when "0100001000010100" => data_out <= rom_array(16916);
		when "0100001000010101" => data_out <= rom_array(16917);
		when "0100001000010110" => data_out <= rom_array(16918);
		when "0100001000010111" => data_out <= rom_array(16919);
		when "0100001000011000" => data_out <= rom_array(16920);
		when "0100001000011001" => data_out <= rom_array(16921);
		when "0100001000011010" => data_out <= rom_array(16922);
		when "0100001000011011" => data_out <= rom_array(16923);
		when "0100001000011100" => data_out <= rom_array(16924);
		when "0100001000011101" => data_out <= rom_array(16925);
		when "0100001000011110" => data_out <= rom_array(16926);
		when "0100001000011111" => data_out <= rom_array(16927);
		when "0100001000100000" => data_out <= rom_array(16928);
		when "0100001000100001" => data_out <= rom_array(16929);
		when "0100001000100010" => data_out <= rom_array(16930);
		when "0100001000100011" => data_out <= rom_array(16931);
		when "0100001000100100" => data_out <= rom_array(16932);
		when "0100001000100101" => data_out <= rom_array(16933);
		when "0100001000100110" => data_out <= rom_array(16934);
		when "0100001000100111" => data_out <= rom_array(16935);
		when "0100001000101000" => data_out <= rom_array(16936);
		when "0100001000101001" => data_out <= rom_array(16937);
		when "0100001000101010" => data_out <= rom_array(16938);
		when "0100001000101011" => data_out <= rom_array(16939);
		when "0100001000101100" => data_out <= rom_array(16940);
		when "0100001000101101" => data_out <= rom_array(16941);
		when "0100001000101110" => data_out <= rom_array(16942);
		when "0100001000101111" => data_out <= rom_array(16943);
		when "0100001000110000" => data_out <= rom_array(16944);
		when "0100001000110001" => data_out <= rom_array(16945);
		when "0100001000110010" => data_out <= rom_array(16946);
		when "0100001000110011" => data_out <= rom_array(16947);
		when "0100001000110100" => data_out <= rom_array(16948);
		when "0100001000110101" => data_out <= rom_array(16949);
		when "0100001000110110" => data_out <= rom_array(16950);
		when "0100001000110111" => data_out <= rom_array(16951);
		when "0100001000111000" => data_out <= rom_array(16952);
		when "0100001000111001" => data_out <= rom_array(16953);
		when "0100001000111010" => data_out <= rom_array(16954);
		when "0100001000111011" => data_out <= rom_array(16955);
		when "0100001000111100" => data_out <= rom_array(16956);
		when "0100001000111101" => data_out <= rom_array(16957);
		when "0100001000111110" => data_out <= rom_array(16958);
		when "0100001000111111" => data_out <= rom_array(16959);
		when "0100001001000000" => data_out <= rom_array(16960);
		when "0100001001000001" => data_out <= rom_array(16961);
		when "0100001001000010" => data_out <= rom_array(16962);
		when "0100001001000011" => data_out <= rom_array(16963);
		when "0100001001000100" => data_out <= rom_array(16964);
		when "0100001001000101" => data_out <= rom_array(16965);
		when "0100001001000110" => data_out <= rom_array(16966);
		when "0100001001000111" => data_out <= rom_array(16967);
		when "0100001001001000" => data_out <= rom_array(16968);
		when "0100001001001001" => data_out <= rom_array(16969);
		when "0100001001001010" => data_out <= rom_array(16970);
		when "0100001001001011" => data_out <= rom_array(16971);
		when "0100001001001100" => data_out <= rom_array(16972);
		when "0100001001001101" => data_out <= rom_array(16973);
		when "0100001001001110" => data_out <= rom_array(16974);
		when "0100001001001111" => data_out <= rom_array(16975);
		when "0100001001010000" => data_out <= rom_array(16976);
		when "0100001001010001" => data_out <= rom_array(16977);
		when "0100001001010010" => data_out <= rom_array(16978);
		when "0100001001010011" => data_out <= rom_array(16979);
		when "0100001001010100" => data_out <= rom_array(16980);
		when "0100001001010101" => data_out <= rom_array(16981);
		when "0100001001010110" => data_out <= rom_array(16982);
		when "0100001001010111" => data_out <= rom_array(16983);
		when "0100001001011000" => data_out <= rom_array(16984);
		when "0100001001011001" => data_out <= rom_array(16985);
		when "0100001001011010" => data_out <= rom_array(16986);
		when "0100001001011011" => data_out <= rom_array(16987);
		when "0100001001011100" => data_out <= rom_array(16988);
		when "0100001001011101" => data_out <= rom_array(16989);
		when "0100001001011110" => data_out <= rom_array(16990);
		when "0100001001011111" => data_out <= rom_array(16991);
		when "0100001001100000" => data_out <= rom_array(16992);
		when "0100001001100001" => data_out <= rom_array(16993);
		when "0100001001100010" => data_out <= rom_array(16994);
		when "0100001001100011" => data_out <= rom_array(16995);
		when "0100001001100100" => data_out <= rom_array(16996);
		when "0100001001100101" => data_out <= rom_array(16997);
		when "0100001001100110" => data_out <= rom_array(16998);
		when "0100001001100111" => data_out <= rom_array(16999);
		when "0100001001101000" => data_out <= rom_array(17000);
		when "0100001001101001" => data_out <= rom_array(17001);
		when "0100001001101010" => data_out <= rom_array(17002);
		when "0100001001101011" => data_out <= rom_array(17003);
		when "0100001001101100" => data_out <= rom_array(17004);
		when "0100001001101101" => data_out <= rom_array(17005);
		when "0100001001101110" => data_out <= rom_array(17006);
		when "0100001001101111" => data_out <= rom_array(17007);
		when "0100001001110000" => data_out <= rom_array(17008);
		when "0100001001110001" => data_out <= rom_array(17009);
		when "0100001001110010" => data_out <= rom_array(17010);
		when "0100001001110011" => data_out <= rom_array(17011);
		when "0100001001110100" => data_out <= rom_array(17012);
		when "0100001001110101" => data_out <= rom_array(17013);
		when "0100001001110110" => data_out <= rom_array(17014);
		when "0100001001110111" => data_out <= rom_array(17015);
		when "0100001001111000" => data_out <= rom_array(17016);
		when "0100001001111001" => data_out <= rom_array(17017);
		when "0100001001111010" => data_out <= rom_array(17018);
		when "0100001001111011" => data_out <= rom_array(17019);
		when "0100001001111100" => data_out <= rom_array(17020);
		when "0100001001111101" => data_out <= rom_array(17021);
		when "0100001001111110" => data_out <= rom_array(17022);
		when "0100001001111111" => data_out <= rom_array(17023);
		when "0100001010000000" => data_out <= rom_array(17024);
		when "0100001010000001" => data_out <= rom_array(17025);
		when "0100001010000010" => data_out <= rom_array(17026);
		when "0100001010000011" => data_out <= rom_array(17027);
		when "0100001010000100" => data_out <= rom_array(17028);
		when "0100001010000101" => data_out <= rom_array(17029);
		when "0100001010000110" => data_out <= rom_array(17030);
		when "0100001010000111" => data_out <= rom_array(17031);
		when "0100001010001000" => data_out <= rom_array(17032);
		when "0100001010001001" => data_out <= rom_array(17033);
		when "0100001010001010" => data_out <= rom_array(17034);
		when "0100001010001011" => data_out <= rom_array(17035);
		when "0100001010001100" => data_out <= rom_array(17036);
		when "0100001010001101" => data_out <= rom_array(17037);
		when "0100001010001110" => data_out <= rom_array(17038);
		when "0100001010001111" => data_out <= rom_array(17039);
		when "0100001010010000" => data_out <= rom_array(17040);
		when "0100001010010001" => data_out <= rom_array(17041);
		when "0100001010010010" => data_out <= rom_array(17042);
		when "0100001010010011" => data_out <= rom_array(17043);
		when "0100001010010100" => data_out <= rom_array(17044);
		when "0100001010010101" => data_out <= rom_array(17045);
		when "0100001010010110" => data_out <= rom_array(17046);
		when "0100001010010111" => data_out <= rom_array(17047);
		when "0100001010011000" => data_out <= rom_array(17048);
		when "0100001010011001" => data_out <= rom_array(17049);
		when "0100001010011010" => data_out <= rom_array(17050);
		when "0100001010011011" => data_out <= rom_array(17051);
		when "0100001010011100" => data_out <= rom_array(17052);
		when "0100001010011101" => data_out <= rom_array(17053);
		when "0100001010011110" => data_out <= rom_array(17054);
		when "0100001010011111" => data_out <= rom_array(17055);
		when "0100001010100000" => data_out <= rom_array(17056);
		when "0100001010100001" => data_out <= rom_array(17057);
		when "0100001010100010" => data_out <= rom_array(17058);
		when "0100001010100011" => data_out <= rom_array(17059);
		when "0100001010100100" => data_out <= rom_array(17060);
		when "0100001010100101" => data_out <= rom_array(17061);
		when "0100001010100110" => data_out <= rom_array(17062);
		when "0100001010100111" => data_out <= rom_array(17063);
		when "0100001010101000" => data_out <= rom_array(17064);
		when "0100001010101001" => data_out <= rom_array(17065);
		when "0100001010101010" => data_out <= rom_array(17066);
		when "0100001010101011" => data_out <= rom_array(17067);
		when "0100001010101100" => data_out <= rom_array(17068);
		when "0100001010101101" => data_out <= rom_array(17069);
		when "0100001010101110" => data_out <= rom_array(17070);
		when "0100001010101111" => data_out <= rom_array(17071);
		when "0100001010110000" => data_out <= rom_array(17072);
		when "0100001010110001" => data_out <= rom_array(17073);
		when "0100001010110010" => data_out <= rom_array(17074);
		when "0100001010110011" => data_out <= rom_array(17075);
		when "0100001010110100" => data_out <= rom_array(17076);
		when "0100001010110101" => data_out <= rom_array(17077);
		when "0100001010110110" => data_out <= rom_array(17078);
		when "0100001010110111" => data_out <= rom_array(17079);
		when "0100001010111000" => data_out <= rom_array(17080);
		when "0100001010111001" => data_out <= rom_array(17081);
		when "0100001010111010" => data_out <= rom_array(17082);
		when "0100001010111011" => data_out <= rom_array(17083);
		when "0100001010111100" => data_out <= rom_array(17084);
		when "0100001010111101" => data_out <= rom_array(17085);
		when "0100001010111110" => data_out <= rom_array(17086);
		when "0100001010111111" => data_out <= rom_array(17087);
		when "0100001011000000" => data_out <= rom_array(17088);
		when "0100001011000001" => data_out <= rom_array(17089);
		when "0100001011000010" => data_out <= rom_array(17090);
		when "0100001011000011" => data_out <= rom_array(17091);
		when "0100001011000100" => data_out <= rom_array(17092);
		when "0100001011000101" => data_out <= rom_array(17093);
		when "0100001011000110" => data_out <= rom_array(17094);
		when "0100001011000111" => data_out <= rom_array(17095);
		when "0100001011001000" => data_out <= rom_array(17096);
		when "0100001011001001" => data_out <= rom_array(17097);
		when "0100001011001010" => data_out <= rom_array(17098);
		when "0100001011001011" => data_out <= rom_array(17099);
		when "0100001011001100" => data_out <= rom_array(17100);
		when "0100001011001101" => data_out <= rom_array(17101);
		when "0100001011001110" => data_out <= rom_array(17102);
		when "0100001011001111" => data_out <= rom_array(17103);
		when "0100001011010000" => data_out <= rom_array(17104);
		when "0100001011010001" => data_out <= rom_array(17105);
		when "0100001011010010" => data_out <= rom_array(17106);
		when "0100001011010011" => data_out <= rom_array(17107);
		when "0100001011010100" => data_out <= rom_array(17108);
		when "0100001011010101" => data_out <= rom_array(17109);
		when "0100001011010110" => data_out <= rom_array(17110);
		when "0100001011010111" => data_out <= rom_array(17111);
		when "0100001011011000" => data_out <= rom_array(17112);
		when "0100001011011001" => data_out <= rom_array(17113);
		when "0100001011011010" => data_out <= rom_array(17114);
		when "0100001011011011" => data_out <= rom_array(17115);
		when "0100001011011100" => data_out <= rom_array(17116);
		when "0100001011011101" => data_out <= rom_array(17117);
		when "0100001011011110" => data_out <= rom_array(17118);
		when "0100001011011111" => data_out <= rom_array(17119);
		when "0100001011100000" => data_out <= rom_array(17120);
		when "0100001011100001" => data_out <= rom_array(17121);
		when "0100001011100010" => data_out <= rom_array(17122);
		when "0100001011100011" => data_out <= rom_array(17123);
		when "0100001011100100" => data_out <= rom_array(17124);
		when "0100001011100101" => data_out <= rom_array(17125);
		when "0100001011100110" => data_out <= rom_array(17126);
		when "0100001011100111" => data_out <= rom_array(17127);
		when "0100001011101000" => data_out <= rom_array(17128);
		when "0100001011101001" => data_out <= rom_array(17129);
		when "0100001011101010" => data_out <= rom_array(17130);
		when "0100001011101011" => data_out <= rom_array(17131);
		when "0100001011101100" => data_out <= rom_array(17132);
		when "0100001011101101" => data_out <= rom_array(17133);
		when "0100001011101110" => data_out <= rom_array(17134);
		when "0100001011101111" => data_out <= rom_array(17135);
		when "0100001011110000" => data_out <= rom_array(17136);
		when "0100001011110001" => data_out <= rom_array(17137);
		when "0100001011110010" => data_out <= rom_array(17138);
		when "0100001011110011" => data_out <= rom_array(17139);
		when "0100001011110100" => data_out <= rom_array(17140);
		when "0100001011110101" => data_out <= rom_array(17141);
		when "0100001011110110" => data_out <= rom_array(17142);
		when "0100001011110111" => data_out <= rom_array(17143);
		when "0100001011111000" => data_out <= rom_array(17144);
		when "0100001011111001" => data_out <= rom_array(17145);
		when "0100001011111010" => data_out <= rom_array(17146);
		when "0100001011111011" => data_out <= rom_array(17147);
		when "0100001011111100" => data_out <= rom_array(17148);
		when "0100001011111101" => data_out <= rom_array(17149);
		when "0100001011111110" => data_out <= rom_array(17150);
		when "0100001011111111" => data_out <= rom_array(17151);
		when "0100001100000000" => data_out <= rom_array(17152);
		when "0100001100000001" => data_out <= rom_array(17153);
		when "0100001100000010" => data_out <= rom_array(17154);
		when "0100001100000011" => data_out <= rom_array(17155);
		when "0100001100000100" => data_out <= rom_array(17156);
		when "0100001100000101" => data_out <= rom_array(17157);
		when "0100001100000110" => data_out <= rom_array(17158);
		when "0100001100000111" => data_out <= rom_array(17159);
		when "0100001100001000" => data_out <= rom_array(17160);
		when "0100001100001001" => data_out <= rom_array(17161);
		when "0100001100001010" => data_out <= rom_array(17162);
		when "0100001100001011" => data_out <= rom_array(17163);
		when "0100001100001100" => data_out <= rom_array(17164);
		when "0100001100001101" => data_out <= rom_array(17165);
		when "0100001100001110" => data_out <= rom_array(17166);
		when "0100001100001111" => data_out <= rom_array(17167);
		when "0100001100010000" => data_out <= rom_array(17168);
		when "0100001100010001" => data_out <= rom_array(17169);
		when "0100001100010010" => data_out <= rom_array(17170);
		when "0100001100010011" => data_out <= rom_array(17171);
		when "0100001100010100" => data_out <= rom_array(17172);
		when "0100001100010101" => data_out <= rom_array(17173);
		when "0100001100010110" => data_out <= rom_array(17174);
		when "0100001100010111" => data_out <= rom_array(17175);
		when "0100001100011000" => data_out <= rom_array(17176);
		when "0100001100011001" => data_out <= rom_array(17177);
		when "0100001100011010" => data_out <= rom_array(17178);
		when "0100001100011011" => data_out <= rom_array(17179);
		when "0100001100011100" => data_out <= rom_array(17180);
		when "0100001100011101" => data_out <= rom_array(17181);
		when "0100001100011110" => data_out <= rom_array(17182);
		when "0100001100011111" => data_out <= rom_array(17183);
		when "0100001100100000" => data_out <= rom_array(17184);
		when "0100001100100001" => data_out <= rom_array(17185);
		when "0100001100100010" => data_out <= rom_array(17186);
		when "0100001100100011" => data_out <= rom_array(17187);
		when "0100001100100100" => data_out <= rom_array(17188);
		when "0100001100100101" => data_out <= rom_array(17189);
		when "0100001100100110" => data_out <= rom_array(17190);
		when "0100001100100111" => data_out <= rom_array(17191);
		when "0100001100101000" => data_out <= rom_array(17192);
		when "0100001100101001" => data_out <= rom_array(17193);
		when "0100001100101010" => data_out <= rom_array(17194);
		when "0100001100101011" => data_out <= rom_array(17195);
		when "0100001100101100" => data_out <= rom_array(17196);
		when "0100001100101101" => data_out <= rom_array(17197);
		when "0100001100101110" => data_out <= rom_array(17198);
		when "0100001100101111" => data_out <= rom_array(17199);
		when "0100001100110000" => data_out <= rom_array(17200);
		when "0100001100110001" => data_out <= rom_array(17201);
		when "0100001100110010" => data_out <= rom_array(17202);
		when "0100001100110011" => data_out <= rom_array(17203);
		when "0100001100110100" => data_out <= rom_array(17204);
		when "0100001100110101" => data_out <= rom_array(17205);
		when "0100001100110110" => data_out <= rom_array(17206);
		when "0100001100110111" => data_out <= rom_array(17207);
		when "0100001100111000" => data_out <= rom_array(17208);
		when "0100001100111001" => data_out <= rom_array(17209);
		when "0100001100111010" => data_out <= rom_array(17210);
		when "0100001100111011" => data_out <= rom_array(17211);
		when "0100001100111100" => data_out <= rom_array(17212);
		when "0100001100111101" => data_out <= rom_array(17213);
		when "0100001100111110" => data_out <= rom_array(17214);
		when "0100001100111111" => data_out <= rom_array(17215);
		when "0100001101000000" => data_out <= rom_array(17216);
		when "0100001101000001" => data_out <= rom_array(17217);
		when "0100001101000010" => data_out <= rom_array(17218);
		when "0100001101000011" => data_out <= rom_array(17219);
		when "0100001101000100" => data_out <= rom_array(17220);
		when "0100001101000101" => data_out <= rom_array(17221);
		when "0100001101000110" => data_out <= rom_array(17222);
		when "0100001101000111" => data_out <= rom_array(17223);
		when "0100001101001000" => data_out <= rom_array(17224);
		when "0100001101001001" => data_out <= rom_array(17225);
		when "0100001101001010" => data_out <= rom_array(17226);
		when "0100001101001011" => data_out <= rom_array(17227);
		when "0100001101001100" => data_out <= rom_array(17228);
		when "0100001101001101" => data_out <= rom_array(17229);
		when "0100001101001110" => data_out <= rom_array(17230);
		when "0100001101001111" => data_out <= rom_array(17231);
		when "0100001101010000" => data_out <= rom_array(17232);
		when "0100001101010001" => data_out <= rom_array(17233);
		when "0100001101010010" => data_out <= rom_array(17234);
		when "0100001101010011" => data_out <= rom_array(17235);
		when "0100001101010100" => data_out <= rom_array(17236);
		when "0100001101010101" => data_out <= rom_array(17237);
		when "0100001101010110" => data_out <= rom_array(17238);
		when "0100001101010111" => data_out <= rom_array(17239);
		when "0100001101011000" => data_out <= rom_array(17240);
		when "0100001101011001" => data_out <= rom_array(17241);
		when "0100001101011010" => data_out <= rom_array(17242);
		when "0100001101011011" => data_out <= rom_array(17243);
		when "0100001101011100" => data_out <= rom_array(17244);
		when "0100001101011101" => data_out <= rom_array(17245);
		when "0100001101011110" => data_out <= rom_array(17246);
		when "0100001101011111" => data_out <= rom_array(17247);
		when "0100001101100000" => data_out <= rom_array(17248);
		when "0100001101100001" => data_out <= rom_array(17249);
		when "0100001101100010" => data_out <= rom_array(17250);
		when "0100001101100011" => data_out <= rom_array(17251);
		when "0100001101100100" => data_out <= rom_array(17252);
		when "0100001101100101" => data_out <= rom_array(17253);
		when "0100001101100110" => data_out <= rom_array(17254);
		when "0100001101100111" => data_out <= rom_array(17255);
		when "0100001101101000" => data_out <= rom_array(17256);
		when "0100001101101001" => data_out <= rom_array(17257);
		when "0100001101101010" => data_out <= rom_array(17258);
		when "0100001101101011" => data_out <= rom_array(17259);
		when "0100001101101100" => data_out <= rom_array(17260);
		when "0100001101101101" => data_out <= rom_array(17261);
		when "0100001101101110" => data_out <= rom_array(17262);
		when "0100001101101111" => data_out <= rom_array(17263);
		when "0100001101110000" => data_out <= rom_array(17264);
		when "0100001101110001" => data_out <= rom_array(17265);
		when "0100001101110010" => data_out <= rom_array(17266);
		when "0100001101110011" => data_out <= rom_array(17267);
		when "0100001101110100" => data_out <= rom_array(17268);
		when "0100001101110101" => data_out <= rom_array(17269);
		when "0100001101110110" => data_out <= rom_array(17270);
		when "0100001101110111" => data_out <= rom_array(17271);
		when "0100001101111000" => data_out <= rom_array(17272);
		when "0100001101111001" => data_out <= rom_array(17273);
		when "0100001101111010" => data_out <= rom_array(17274);
		when "0100001101111011" => data_out <= rom_array(17275);
		when "0100001101111100" => data_out <= rom_array(17276);
		when "0100001101111101" => data_out <= rom_array(17277);
		when "0100001101111110" => data_out <= rom_array(17278);
		when "0100001101111111" => data_out <= rom_array(17279);
		when "0100001110000000" => data_out <= rom_array(17280);
		when "0100001110000001" => data_out <= rom_array(17281);
		when "0100001110000010" => data_out <= rom_array(17282);
		when "0100001110000011" => data_out <= rom_array(17283);
		when "0100001110000100" => data_out <= rom_array(17284);
		when "0100001110000101" => data_out <= rom_array(17285);
		when "0100001110000110" => data_out <= rom_array(17286);
		when "0100001110000111" => data_out <= rom_array(17287);
		when "0100001110001000" => data_out <= rom_array(17288);
		when "0100001110001001" => data_out <= rom_array(17289);
		when "0100001110001010" => data_out <= rom_array(17290);
		when "0100001110001011" => data_out <= rom_array(17291);
		when "0100001110001100" => data_out <= rom_array(17292);
		when "0100001110001101" => data_out <= rom_array(17293);
		when "0100001110001110" => data_out <= rom_array(17294);
		when "0100001110001111" => data_out <= rom_array(17295);
		when "0100001110010000" => data_out <= rom_array(17296);
		when "0100001110010001" => data_out <= rom_array(17297);
		when "0100001110010010" => data_out <= rom_array(17298);
		when "0100001110010011" => data_out <= rom_array(17299);
		when "0100001110010100" => data_out <= rom_array(17300);
		when "0100001110010101" => data_out <= rom_array(17301);
		when "0100001110010110" => data_out <= rom_array(17302);
		when "0100001110010111" => data_out <= rom_array(17303);
		when "0100001110011000" => data_out <= rom_array(17304);
		when "0100001110011001" => data_out <= rom_array(17305);
		when "0100001110011010" => data_out <= rom_array(17306);
		when "0100001110011011" => data_out <= rom_array(17307);
		when "0100001110011100" => data_out <= rom_array(17308);
		when "0100001110011101" => data_out <= rom_array(17309);
		when "0100001110011110" => data_out <= rom_array(17310);
		when "0100001110011111" => data_out <= rom_array(17311);
		when "0100001110100000" => data_out <= rom_array(17312);
		when "0100001110100001" => data_out <= rom_array(17313);
		when "0100001110100010" => data_out <= rom_array(17314);
		when "0100001110100011" => data_out <= rom_array(17315);
		when "0100001110100100" => data_out <= rom_array(17316);
		when "0100001110100101" => data_out <= rom_array(17317);
		when "0100001110100110" => data_out <= rom_array(17318);
		when "0100001110100111" => data_out <= rom_array(17319);
		when "0100001110101000" => data_out <= rom_array(17320);
		when "0100001110101001" => data_out <= rom_array(17321);
		when "0100001110101010" => data_out <= rom_array(17322);
		when "0100001110101011" => data_out <= rom_array(17323);
		when "0100001110101100" => data_out <= rom_array(17324);
		when "0100001110101101" => data_out <= rom_array(17325);
		when "0100001110101110" => data_out <= rom_array(17326);
		when "0100001110101111" => data_out <= rom_array(17327);
		when "0100001110110000" => data_out <= rom_array(17328);
		when "0100001110110001" => data_out <= rom_array(17329);
		when "0100001110110010" => data_out <= rom_array(17330);
		when "0100001110110011" => data_out <= rom_array(17331);
		when "0100001110110100" => data_out <= rom_array(17332);
		when "0100001110110101" => data_out <= rom_array(17333);
		when "0100001110110110" => data_out <= rom_array(17334);
		when "0100001110110111" => data_out <= rom_array(17335);
		when "0100001110111000" => data_out <= rom_array(17336);
		when "0100001110111001" => data_out <= rom_array(17337);
		when "0100001110111010" => data_out <= rom_array(17338);
		when "0100001110111011" => data_out <= rom_array(17339);
		when "0100001110111100" => data_out <= rom_array(17340);
		when "0100001110111101" => data_out <= rom_array(17341);
		when "0100001110111110" => data_out <= rom_array(17342);
		when "0100001110111111" => data_out <= rom_array(17343);
		when "0100001111000000" => data_out <= rom_array(17344);
		when "0100001111000001" => data_out <= rom_array(17345);
		when "0100001111000010" => data_out <= rom_array(17346);
		when "0100001111000011" => data_out <= rom_array(17347);
		when "0100001111000100" => data_out <= rom_array(17348);
		when "0100001111000101" => data_out <= rom_array(17349);
		when "0100001111000110" => data_out <= rom_array(17350);
		when "0100001111000111" => data_out <= rom_array(17351);
		when "0100001111001000" => data_out <= rom_array(17352);
		when "0100001111001001" => data_out <= rom_array(17353);
		when "0100001111001010" => data_out <= rom_array(17354);
		when "0100001111001011" => data_out <= rom_array(17355);
		when "0100001111001100" => data_out <= rom_array(17356);
		when "0100001111001101" => data_out <= rom_array(17357);
		when "0100001111001110" => data_out <= rom_array(17358);
		when "0100001111001111" => data_out <= rom_array(17359);
		when "0100001111010000" => data_out <= rom_array(17360);
		when "0100001111010001" => data_out <= rom_array(17361);
		when "0100001111010010" => data_out <= rom_array(17362);
		when "0100001111010011" => data_out <= rom_array(17363);
		when "0100001111010100" => data_out <= rom_array(17364);
		when "0100001111010101" => data_out <= rom_array(17365);
		when "0100001111010110" => data_out <= rom_array(17366);
		when "0100001111010111" => data_out <= rom_array(17367);
		when "0100001111011000" => data_out <= rom_array(17368);
		when "0100001111011001" => data_out <= rom_array(17369);
		when "0100001111011010" => data_out <= rom_array(17370);
		when "0100001111011011" => data_out <= rom_array(17371);
		when "0100001111011100" => data_out <= rom_array(17372);
		when "0100001111011101" => data_out <= rom_array(17373);
		when "0100001111011110" => data_out <= rom_array(17374);
		when "0100001111011111" => data_out <= rom_array(17375);
		when "0100001111100000" => data_out <= rom_array(17376);
		when "0100001111100001" => data_out <= rom_array(17377);
		when "0100001111100010" => data_out <= rom_array(17378);
		when "0100001111100011" => data_out <= rom_array(17379);
		when "0100001111100100" => data_out <= rom_array(17380);
		when "0100001111100101" => data_out <= rom_array(17381);
		when "0100001111100110" => data_out <= rom_array(17382);
		when "0100001111100111" => data_out <= rom_array(17383);
		when "0100001111101000" => data_out <= rom_array(17384);
		when "0100001111101001" => data_out <= rom_array(17385);
		when "0100001111101010" => data_out <= rom_array(17386);
		when "0100001111101011" => data_out <= rom_array(17387);
		when "0100001111101100" => data_out <= rom_array(17388);
		when "0100001111101101" => data_out <= rom_array(17389);
		when "0100001111101110" => data_out <= rom_array(17390);
		when "0100001111101111" => data_out <= rom_array(17391);
		when "0100001111110000" => data_out <= rom_array(17392);
		when "0100001111110001" => data_out <= rom_array(17393);
		when "0100001111110010" => data_out <= rom_array(17394);
		when "0100001111110011" => data_out <= rom_array(17395);
		when "0100001111110100" => data_out <= rom_array(17396);
		when "0100001111110101" => data_out <= rom_array(17397);
		when "0100001111110110" => data_out <= rom_array(17398);
		when "0100001111110111" => data_out <= rom_array(17399);
		when "0100001111111000" => data_out <= rom_array(17400);
		when "0100001111111001" => data_out <= rom_array(17401);
		when "0100001111111010" => data_out <= rom_array(17402);
		when "0100001111111011" => data_out <= rom_array(17403);
		when "0100001111111100" => data_out <= rom_array(17404);
		when "0100001111111101" => data_out <= rom_array(17405);
		when "0100001111111110" => data_out <= rom_array(17406);
		when "0100001111111111" => data_out <= rom_array(17407);
		when "0100010000000000" => data_out <= rom_array(17408);
		when "0100010000000001" => data_out <= rom_array(17409);
		when "0100010000000010" => data_out <= rom_array(17410);
		when "0100010000000011" => data_out <= rom_array(17411);
		when "0100010000000100" => data_out <= rom_array(17412);
		when "0100010000000101" => data_out <= rom_array(17413);
		when "0100010000000110" => data_out <= rom_array(17414);
		when "0100010000000111" => data_out <= rom_array(17415);
		when "0100010000001000" => data_out <= rom_array(17416);
		when "0100010000001001" => data_out <= rom_array(17417);
		when "0100010000001010" => data_out <= rom_array(17418);
		when "0100010000001011" => data_out <= rom_array(17419);
		when "0100010000001100" => data_out <= rom_array(17420);
		when "0100010000001101" => data_out <= rom_array(17421);
		when "0100010000001110" => data_out <= rom_array(17422);
		when "0100010000001111" => data_out <= rom_array(17423);
		when "0100010000010000" => data_out <= rom_array(17424);
		when "0100010000010001" => data_out <= rom_array(17425);
		when "0100010000010010" => data_out <= rom_array(17426);
		when "0100010000010011" => data_out <= rom_array(17427);
		when "0100010000010100" => data_out <= rom_array(17428);
		when "0100010000010101" => data_out <= rom_array(17429);
		when "0100010000010110" => data_out <= rom_array(17430);
		when "0100010000010111" => data_out <= rom_array(17431);
		when "0100010000011000" => data_out <= rom_array(17432);
		when "0100010000011001" => data_out <= rom_array(17433);
		when "0100010000011010" => data_out <= rom_array(17434);
		when "0100010000011011" => data_out <= rom_array(17435);
		when "0100010000011100" => data_out <= rom_array(17436);
		when "0100010000011101" => data_out <= rom_array(17437);
		when "0100010000011110" => data_out <= rom_array(17438);
		when "0100010000011111" => data_out <= rom_array(17439);
		when "0100010000100000" => data_out <= rom_array(17440);
		when "0100010000100001" => data_out <= rom_array(17441);
		when "0100010000100010" => data_out <= rom_array(17442);
		when "0100010000100011" => data_out <= rom_array(17443);
		when "0100010000100100" => data_out <= rom_array(17444);
		when "0100010000100101" => data_out <= rom_array(17445);
		when "0100010000100110" => data_out <= rom_array(17446);
		when "0100010000100111" => data_out <= rom_array(17447);
		when "0100010000101000" => data_out <= rom_array(17448);
		when "0100010000101001" => data_out <= rom_array(17449);
		when "0100010000101010" => data_out <= rom_array(17450);
		when "0100010000101011" => data_out <= rom_array(17451);
		when "0100010000101100" => data_out <= rom_array(17452);
		when "0100010000101101" => data_out <= rom_array(17453);
		when "0100010000101110" => data_out <= rom_array(17454);
		when "0100010000101111" => data_out <= rom_array(17455);
		when "0100010000110000" => data_out <= rom_array(17456);
		when "0100010000110001" => data_out <= rom_array(17457);
		when "0100010000110010" => data_out <= rom_array(17458);
		when "0100010000110011" => data_out <= rom_array(17459);
		when "0100010000110100" => data_out <= rom_array(17460);
		when "0100010000110101" => data_out <= rom_array(17461);
		when "0100010000110110" => data_out <= rom_array(17462);
		when "0100010000110111" => data_out <= rom_array(17463);
		when "0100010000111000" => data_out <= rom_array(17464);
		when "0100010000111001" => data_out <= rom_array(17465);
		when "0100010000111010" => data_out <= rom_array(17466);
		when "0100010000111011" => data_out <= rom_array(17467);
		when "0100010000111100" => data_out <= rom_array(17468);
		when "0100010000111101" => data_out <= rom_array(17469);
		when "0100010000111110" => data_out <= rom_array(17470);
		when "0100010000111111" => data_out <= rom_array(17471);
		when "0100010001000000" => data_out <= rom_array(17472);
		when "0100010001000001" => data_out <= rom_array(17473);
		when "0100010001000010" => data_out <= rom_array(17474);
		when "0100010001000011" => data_out <= rom_array(17475);
		when "0100010001000100" => data_out <= rom_array(17476);
		when "0100010001000101" => data_out <= rom_array(17477);
		when "0100010001000110" => data_out <= rom_array(17478);
		when "0100010001000111" => data_out <= rom_array(17479);
		when "0100010001001000" => data_out <= rom_array(17480);
		when "0100010001001001" => data_out <= rom_array(17481);
		when "0100010001001010" => data_out <= rom_array(17482);
		when "0100010001001011" => data_out <= rom_array(17483);
		when "0100010001001100" => data_out <= rom_array(17484);
		when "0100010001001101" => data_out <= rom_array(17485);
		when "0100010001001110" => data_out <= rom_array(17486);
		when "0100010001001111" => data_out <= rom_array(17487);
		when "0100010001010000" => data_out <= rom_array(17488);
		when "0100010001010001" => data_out <= rom_array(17489);
		when "0100010001010010" => data_out <= rom_array(17490);
		when "0100010001010011" => data_out <= rom_array(17491);
		when "0100010001010100" => data_out <= rom_array(17492);
		when "0100010001010101" => data_out <= rom_array(17493);
		when "0100010001010110" => data_out <= rom_array(17494);
		when "0100010001010111" => data_out <= rom_array(17495);
		when "0100010001011000" => data_out <= rom_array(17496);
		when "0100010001011001" => data_out <= rom_array(17497);
		when "0100010001011010" => data_out <= rom_array(17498);
		when "0100010001011011" => data_out <= rom_array(17499);
		when "0100010001011100" => data_out <= rom_array(17500);
		when "0100010001011101" => data_out <= rom_array(17501);
		when "0100010001011110" => data_out <= rom_array(17502);
		when "0100010001011111" => data_out <= rom_array(17503);
		when "0100010001100000" => data_out <= rom_array(17504);
		when "0100010001100001" => data_out <= rom_array(17505);
		when "0100010001100010" => data_out <= rom_array(17506);
		when "0100010001100011" => data_out <= rom_array(17507);
		when "0100010001100100" => data_out <= rom_array(17508);
		when "0100010001100101" => data_out <= rom_array(17509);
		when "0100010001100110" => data_out <= rom_array(17510);
		when "0100010001100111" => data_out <= rom_array(17511);
		when "0100010001101000" => data_out <= rom_array(17512);
		when "0100010001101001" => data_out <= rom_array(17513);
		when "0100010001101010" => data_out <= rom_array(17514);
		when "0100010001101011" => data_out <= rom_array(17515);
		when "0100010001101100" => data_out <= rom_array(17516);
		when "0100010001101101" => data_out <= rom_array(17517);
		when "0100010001101110" => data_out <= rom_array(17518);
		when "0100010001101111" => data_out <= rom_array(17519);
		when "0100010001110000" => data_out <= rom_array(17520);
		when "0100010001110001" => data_out <= rom_array(17521);
		when "0100010001110010" => data_out <= rom_array(17522);
		when "0100010001110011" => data_out <= rom_array(17523);
		when "0100010001110100" => data_out <= rom_array(17524);
		when "0100010001110101" => data_out <= rom_array(17525);
		when "0100010001110110" => data_out <= rom_array(17526);
		when "0100010001110111" => data_out <= rom_array(17527);
		when "0100010001111000" => data_out <= rom_array(17528);
		when "0100010001111001" => data_out <= rom_array(17529);
		when "0100010001111010" => data_out <= rom_array(17530);
		when "0100010001111011" => data_out <= rom_array(17531);
		when "0100010001111100" => data_out <= rom_array(17532);
		when "0100010001111101" => data_out <= rom_array(17533);
		when "0100010001111110" => data_out <= rom_array(17534);
		when "0100010001111111" => data_out <= rom_array(17535);
		when "0100010010000000" => data_out <= rom_array(17536);
		when "0100010010000001" => data_out <= rom_array(17537);
		when "0100010010000010" => data_out <= rom_array(17538);
		when "0100010010000011" => data_out <= rom_array(17539);
		when "0100010010000100" => data_out <= rom_array(17540);
		when "0100010010000101" => data_out <= rom_array(17541);
		when "0100010010000110" => data_out <= rom_array(17542);
		when "0100010010000111" => data_out <= rom_array(17543);
		when "0100010010001000" => data_out <= rom_array(17544);
		when "0100010010001001" => data_out <= rom_array(17545);
		when "0100010010001010" => data_out <= rom_array(17546);
		when "0100010010001011" => data_out <= rom_array(17547);
		when "0100010010001100" => data_out <= rom_array(17548);
		when "0100010010001101" => data_out <= rom_array(17549);
		when "0100010010001110" => data_out <= rom_array(17550);
		when "0100010010001111" => data_out <= rom_array(17551);
		when "0100010010010000" => data_out <= rom_array(17552);
		when "0100010010010001" => data_out <= rom_array(17553);
		when "0100010010010010" => data_out <= rom_array(17554);
		when "0100010010010011" => data_out <= rom_array(17555);
		when "0100010010010100" => data_out <= rom_array(17556);
		when "0100010010010101" => data_out <= rom_array(17557);
		when "0100010010010110" => data_out <= rom_array(17558);
		when "0100010010010111" => data_out <= rom_array(17559);
		when "0100010010011000" => data_out <= rom_array(17560);
		when "0100010010011001" => data_out <= rom_array(17561);
		when "0100010010011010" => data_out <= rom_array(17562);
		when "0100010010011011" => data_out <= rom_array(17563);
		when "0100010010011100" => data_out <= rom_array(17564);
		when "0100010010011101" => data_out <= rom_array(17565);
		when "0100010010011110" => data_out <= rom_array(17566);
		when "0100010010011111" => data_out <= rom_array(17567);
		when "0100010010100000" => data_out <= rom_array(17568);
		when "0100010010100001" => data_out <= rom_array(17569);
		when "0100010010100010" => data_out <= rom_array(17570);
		when "0100010010100011" => data_out <= rom_array(17571);
		when "0100010010100100" => data_out <= rom_array(17572);
		when "0100010010100101" => data_out <= rom_array(17573);
		when "0100010010100110" => data_out <= rom_array(17574);
		when "0100010010100111" => data_out <= rom_array(17575);
		when "0100010010101000" => data_out <= rom_array(17576);
		when "0100010010101001" => data_out <= rom_array(17577);
		when "0100010010101010" => data_out <= rom_array(17578);
		when "0100010010101011" => data_out <= rom_array(17579);
		when "0100010010101100" => data_out <= rom_array(17580);
		when "0100010010101101" => data_out <= rom_array(17581);
		when "0100010010101110" => data_out <= rom_array(17582);
		when "0100010010101111" => data_out <= rom_array(17583);
		when "0100010010110000" => data_out <= rom_array(17584);
		when "0100010010110001" => data_out <= rom_array(17585);
		when "0100010010110010" => data_out <= rom_array(17586);
		when "0100010010110011" => data_out <= rom_array(17587);
		when "0100010010110100" => data_out <= rom_array(17588);
		when "0100010010110101" => data_out <= rom_array(17589);
		when "0100010010110110" => data_out <= rom_array(17590);
		when "0100010010110111" => data_out <= rom_array(17591);
		when "0100010010111000" => data_out <= rom_array(17592);
		when "0100010010111001" => data_out <= rom_array(17593);
		when "0100010010111010" => data_out <= rom_array(17594);
		when "0100010010111011" => data_out <= rom_array(17595);
		when "0100010010111100" => data_out <= rom_array(17596);
		when "0100010010111101" => data_out <= rom_array(17597);
		when "0100010010111110" => data_out <= rom_array(17598);
		when "0100010010111111" => data_out <= rom_array(17599);
		when "0100010011000000" => data_out <= rom_array(17600);
		when "0100010011000001" => data_out <= rom_array(17601);
		when "0100010011000010" => data_out <= rom_array(17602);
		when "0100010011000011" => data_out <= rom_array(17603);
		when "0100010011000100" => data_out <= rom_array(17604);
		when "0100010011000101" => data_out <= rom_array(17605);
		when "0100010011000110" => data_out <= rom_array(17606);
		when "0100010011000111" => data_out <= rom_array(17607);
		when "0100010011001000" => data_out <= rom_array(17608);
		when "0100010011001001" => data_out <= rom_array(17609);
		when "0100010011001010" => data_out <= rom_array(17610);
		when "0100010011001011" => data_out <= rom_array(17611);
		when "0100010011001100" => data_out <= rom_array(17612);
		when "0100010011001101" => data_out <= rom_array(17613);
		when "0100010011001110" => data_out <= rom_array(17614);
		when "0100010011001111" => data_out <= rom_array(17615);
		when "0100010011010000" => data_out <= rom_array(17616);
		when "0100010011010001" => data_out <= rom_array(17617);
		when "0100010011010010" => data_out <= rom_array(17618);
		when "0100010011010011" => data_out <= rom_array(17619);
		when "0100010011010100" => data_out <= rom_array(17620);
		when "0100010011010101" => data_out <= rom_array(17621);
		when "0100010011010110" => data_out <= rom_array(17622);
		when "0100010011010111" => data_out <= rom_array(17623);
		when "0100010011011000" => data_out <= rom_array(17624);
		when "0100010011011001" => data_out <= rom_array(17625);
		when "0100010011011010" => data_out <= rom_array(17626);
		when "0100010011011011" => data_out <= rom_array(17627);
		when "0100010011011100" => data_out <= rom_array(17628);
		when "0100010011011101" => data_out <= rom_array(17629);
		when "0100010011011110" => data_out <= rom_array(17630);
		when "0100010011011111" => data_out <= rom_array(17631);
		when "0100010011100000" => data_out <= rom_array(17632);
		when "0100010011100001" => data_out <= rom_array(17633);
		when "0100010011100010" => data_out <= rom_array(17634);
		when "0100010011100011" => data_out <= rom_array(17635);
		when "0100010011100100" => data_out <= rom_array(17636);
		when "0100010011100101" => data_out <= rom_array(17637);
		when "0100010011100110" => data_out <= rom_array(17638);
		when "0100010011100111" => data_out <= rom_array(17639);
		when "0100010011101000" => data_out <= rom_array(17640);
		when "0100010011101001" => data_out <= rom_array(17641);
		when "0100010011101010" => data_out <= rom_array(17642);
		when "0100010011101011" => data_out <= rom_array(17643);
		when "0100010011101100" => data_out <= rom_array(17644);
		when "0100010011101101" => data_out <= rom_array(17645);
		when "0100010011101110" => data_out <= rom_array(17646);
		when "0100010011101111" => data_out <= rom_array(17647);
		when "0100010011110000" => data_out <= rom_array(17648);
		when "0100010011110001" => data_out <= rom_array(17649);
		when "0100010011110010" => data_out <= rom_array(17650);
		when "0100010011110011" => data_out <= rom_array(17651);
		when "0100010011110100" => data_out <= rom_array(17652);
		when "0100010011110101" => data_out <= rom_array(17653);
		when "0100010011110110" => data_out <= rom_array(17654);
		when "0100010011110111" => data_out <= rom_array(17655);
		when "0100010011111000" => data_out <= rom_array(17656);
		when "0100010011111001" => data_out <= rom_array(17657);
		when "0100010011111010" => data_out <= rom_array(17658);
		when "0100010011111011" => data_out <= rom_array(17659);
		when "0100010011111100" => data_out <= rom_array(17660);
		when "0100010011111101" => data_out <= rom_array(17661);
		when "0100010011111110" => data_out <= rom_array(17662);
		when "0100010011111111" => data_out <= rom_array(17663);
		when "0100010100000000" => data_out <= rom_array(17664);
		when "0100010100000001" => data_out <= rom_array(17665);
		when "0100010100000010" => data_out <= rom_array(17666);
		when "0100010100000011" => data_out <= rom_array(17667);
		when "0100010100000100" => data_out <= rom_array(17668);
		when "0100010100000101" => data_out <= rom_array(17669);
		when "0100010100000110" => data_out <= rom_array(17670);
		when "0100010100000111" => data_out <= rom_array(17671);
		when "0100010100001000" => data_out <= rom_array(17672);
		when "0100010100001001" => data_out <= rom_array(17673);
		when "0100010100001010" => data_out <= rom_array(17674);
		when "0100010100001011" => data_out <= rom_array(17675);
		when "0100010100001100" => data_out <= rom_array(17676);
		when "0100010100001101" => data_out <= rom_array(17677);
		when "0100010100001110" => data_out <= rom_array(17678);
		when "0100010100001111" => data_out <= rom_array(17679);
		when "0100010100010000" => data_out <= rom_array(17680);
		when "0100010100010001" => data_out <= rom_array(17681);
		when "0100010100010010" => data_out <= rom_array(17682);
		when "0100010100010011" => data_out <= rom_array(17683);
		when "0100010100010100" => data_out <= rom_array(17684);
		when "0100010100010101" => data_out <= rom_array(17685);
		when "0100010100010110" => data_out <= rom_array(17686);
		when "0100010100010111" => data_out <= rom_array(17687);
		when "0100010100011000" => data_out <= rom_array(17688);
		when "0100010100011001" => data_out <= rom_array(17689);
		when "0100010100011010" => data_out <= rom_array(17690);
		when "0100010100011011" => data_out <= rom_array(17691);
		when "0100010100011100" => data_out <= rom_array(17692);
		when "0100010100011101" => data_out <= rom_array(17693);
		when "0100010100011110" => data_out <= rom_array(17694);
		when "0100010100011111" => data_out <= rom_array(17695);
		when "0100010100100000" => data_out <= rom_array(17696);
		when "0100010100100001" => data_out <= rom_array(17697);
		when "0100010100100010" => data_out <= rom_array(17698);
		when "0100010100100011" => data_out <= rom_array(17699);
		when "0100010100100100" => data_out <= rom_array(17700);
		when "0100010100100101" => data_out <= rom_array(17701);
		when "0100010100100110" => data_out <= rom_array(17702);
		when "0100010100100111" => data_out <= rom_array(17703);
		when "0100010100101000" => data_out <= rom_array(17704);
		when "0100010100101001" => data_out <= rom_array(17705);
		when "0100010100101010" => data_out <= rom_array(17706);
		when "0100010100101011" => data_out <= rom_array(17707);
		when "0100010100101100" => data_out <= rom_array(17708);
		when "0100010100101101" => data_out <= rom_array(17709);
		when "0100010100101110" => data_out <= rom_array(17710);
		when "0100010100101111" => data_out <= rom_array(17711);
		when "0100010100110000" => data_out <= rom_array(17712);
		when "0100010100110001" => data_out <= rom_array(17713);
		when "0100010100110010" => data_out <= rom_array(17714);
		when "0100010100110011" => data_out <= rom_array(17715);
		when "0100010100110100" => data_out <= rom_array(17716);
		when "0100010100110101" => data_out <= rom_array(17717);
		when "0100010100110110" => data_out <= rom_array(17718);
		when "0100010100110111" => data_out <= rom_array(17719);
		when "0100010100111000" => data_out <= rom_array(17720);
		when "0100010100111001" => data_out <= rom_array(17721);
		when "0100010100111010" => data_out <= rom_array(17722);
		when "0100010100111011" => data_out <= rom_array(17723);
		when "0100010100111100" => data_out <= rom_array(17724);
		when "0100010100111101" => data_out <= rom_array(17725);
		when "0100010100111110" => data_out <= rom_array(17726);
		when "0100010100111111" => data_out <= rom_array(17727);
		when "0100010101000000" => data_out <= rom_array(17728);
		when "0100010101000001" => data_out <= rom_array(17729);
		when "0100010101000010" => data_out <= rom_array(17730);
		when "0100010101000011" => data_out <= rom_array(17731);
		when "0100010101000100" => data_out <= rom_array(17732);
		when "0100010101000101" => data_out <= rom_array(17733);
		when "0100010101000110" => data_out <= rom_array(17734);
		when "0100010101000111" => data_out <= rom_array(17735);
		when "0100010101001000" => data_out <= rom_array(17736);
		when "0100010101001001" => data_out <= rom_array(17737);
		when "0100010101001010" => data_out <= rom_array(17738);
		when "0100010101001011" => data_out <= rom_array(17739);
		when "0100010101001100" => data_out <= rom_array(17740);
		when "0100010101001101" => data_out <= rom_array(17741);
		when "0100010101001110" => data_out <= rom_array(17742);
		when "0100010101001111" => data_out <= rom_array(17743);
		when "0100010101010000" => data_out <= rom_array(17744);
		when "0100010101010001" => data_out <= rom_array(17745);
		when "0100010101010010" => data_out <= rom_array(17746);
		when "0100010101010011" => data_out <= rom_array(17747);
		when "0100010101010100" => data_out <= rom_array(17748);
		when "0100010101010101" => data_out <= rom_array(17749);
		when "0100010101010110" => data_out <= rom_array(17750);
		when "0100010101010111" => data_out <= rom_array(17751);
		when "0100010101011000" => data_out <= rom_array(17752);
		when "0100010101011001" => data_out <= rom_array(17753);
		when "0100010101011010" => data_out <= rom_array(17754);
		when "0100010101011011" => data_out <= rom_array(17755);
		when "0100010101011100" => data_out <= rom_array(17756);
		when "0100010101011101" => data_out <= rom_array(17757);
		when "0100010101011110" => data_out <= rom_array(17758);
		when "0100010101011111" => data_out <= rom_array(17759);
		when "0100010101100000" => data_out <= rom_array(17760);
		when "0100010101100001" => data_out <= rom_array(17761);
		when "0100010101100010" => data_out <= rom_array(17762);
		when "0100010101100011" => data_out <= rom_array(17763);
		when "0100010101100100" => data_out <= rom_array(17764);
		when "0100010101100101" => data_out <= rom_array(17765);
		when "0100010101100110" => data_out <= rom_array(17766);
		when "0100010101100111" => data_out <= rom_array(17767);
		when "0100010101101000" => data_out <= rom_array(17768);
		when "0100010101101001" => data_out <= rom_array(17769);
		when "0100010101101010" => data_out <= rom_array(17770);
		when "0100010101101011" => data_out <= rom_array(17771);
		when "0100010101101100" => data_out <= rom_array(17772);
		when "0100010101101101" => data_out <= rom_array(17773);
		when "0100010101101110" => data_out <= rom_array(17774);
		when "0100010101101111" => data_out <= rom_array(17775);
		when "0100010101110000" => data_out <= rom_array(17776);
		when "0100010101110001" => data_out <= rom_array(17777);
		when "0100010101110010" => data_out <= rom_array(17778);
		when "0100010101110011" => data_out <= rom_array(17779);
		when "0100010101110100" => data_out <= rom_array(17780);
		when "0100010101110101" => data_out <= rom_array(17781);
		when "0100010101110110" => data_out <= rom_array(17782);
		when "0100010101110111" => data_out <= rom_array(17783);
		when "0100010101111000" => data_out <= rom_array(17784);
		when "0100010101111001" => data_out <= rom_array(17785);
		when "0100010101111010" => data_out <= rom_array(17786);
		when "0100010101111011" => data_out <= rom_array(17787);
		when "0100010101111100" => data_out <= rom_array(17788);
		when "0100010101111101" => data_out <= rom_array(17789);
		when "0100010101111110" => data_out <= rom_array(17790);
		when "0100010101111111" => data_out <= rom_array(17791);
		when "0100010110000000" => data_out <= rom_array(17792);
		when "0100010110000001" => data_out <= rom_array(17793);
		when "0100010110000010" => data_out <= rom_array(17794);
		when "0100010110000011" => data_out <= rom_array(17795);
		when "0100010110000100" => data_out <= rom_array(17796);
		when "0100010110000101" => data_out <= rom_array(17797);
		when "0100010110000110" => data_out <= rom_array(17798);
		when "0100010110000111" => data_out <= rom_array(17799);
		when "0100010110001000" => data_out <= rom_array(17800);
		when "0100010110001001" => data_out <= rom_array(17801);
		when "0100010110001010" => data_out <= rom_array(17802);
		when "0100010110001011" => data_out <= rom_array(17803);
		when "0100010110001100" => data_out <= rom_array(17804);
		when "0100010110001101" => data_out <= rom_array(17805);
		when "0100010110001110" => data_out <= rom_array(17806);
		when "0100010110001111" => data_out <= rom_array(17807);
		when "0100010110010000" => data_out <= rom_array(17808);
		when "0100010110010001" => data_out <= rom_array(17809);
		when "0100010110010010" => data_out <= rom_array(17810);
		when "0100010110010011" => data_out <= rom_array(17811);
		when "0100010110010100" => data_out <= rom_array(17812);
		when "0100010110010101" => data_out <= rom_array(17813);
		when "0100010110010110" => data_out <= rom_array(17814);
		when "0100010110010111" => data_out <= rom_array(17815);
		when "0100010110011000" => data_out <= rom_array(17816);
		when "0100010110011001" => data_out <= rom_array(17817);
		when "0100010110011010" => data_out <= rom_array(17818);
		when "0100010110011011" => data_out <= rom_array(17819);
		when "0100010110011100" => data_out <= rom_array(17820);
		when "0100010110011101" => data_out <= rom_array(17821);
		when "0100010110011110" => data_out <= rom_array(17822);
		when "0100010110011111" => data_out <= rom_array(17823);
		when "0100010110100000" => data_out <= rom_array(17824);
		when "0100010110100001" => data_out <= rom_array(17825);
		when "0100010110100010" => data_out <= rom_array(17826);
		when "0100010110100011" => data_out <= rom_array(17827);
		when "0100010110100100" => data_out <= rom_array(17828);
		when "0100010110100101" => data_out <= rom_array(17829);
		when "0100010110100110" => data_out <= rom_array(17830);
		when "0100010110100111" => data_out <= rom_array(17831);
		when "0100010110101000" => data_out <= rom_array(17832);
		when "0100010110101001" => data_out <= rom_array(17833);
		when "0100010110101010" => data_out <= rom_array(17834);
		when "0100010110101011" => data_out <= rom_array(17835);
		when "0100010110101100" => data_out <= rom_array(17836);
		when "0100010110101101" => data_out <= rom_array(17837);
		when "0100010110101110" => data_out <= rom_array(17838);
		when "0100010110101111" => data_out <= rom_array(17839);
		when "0100010110110000" => data_out <= rom_array(17840);
		when "0100010110110001" => data_out <= rom_array(17841);
		when "0100010110110010" => data_out <= rom_array(17842);
		when "0100010110110011" => data_out <= rom_array(17843);
		when "0100010110110100" => data_out <= rom_array(17844);
		when "0100010110110101" => data_out <= rom_array(17845);
		when "0100010110110110" => data_out <= rom_array(17846);
		when "0100010110110111" => data_out <= rom_array(17847);
		when "0100010110111000" => data_out <= rom_array(17848);
		when "0100010110111001" => data_out <= rom_array(17849);
		when "0100010110111010" => data_out <= rom_array(17850);
		when "0100010110111011" => data_out <= rom_array(17851);
		when "0100010110111100" => data_out <= rom_array(17852);
		when "0100010110111101" => data_out <= rom_array(17853);
		when "0100010110111110" => data_out <= rom_array(17854);
		when "0100010110111111" => data_out <= rom_array(17855);
		when "0100010111000000" => data_out <= rom_array(17856);
		when "0100010111000001" => data_out <= rom_array(17857);
		when "0100010111000010" => data_out <= rom_array(17858);
		when "0100010111000011" => data_out <= rom_array(17859);
		when "0100010111000100" => data_out <= rom_array(17860);
		when "0100010111000101" => data_out <= rom_array(17861);
		when "0100010111000110" => data_out <= rom_array(17862);
		when "0100010111000111" => data_out <= rom_array(17863);
		when "0100010111001000" => data_out <= rom_array(17864);
		when "0100010111001001" => data_out <= rom_array(17865);
		when "0100010111001010" => data_out <= rom_array(17866);
		when "0100010111001011" => data_out <= rom_array(17867);
		when "0100010111001100" => data_out <= rom_array(17868);
		when "0100010111001101" => data_out <= rom_array(17869);
		when "0100010111001110" => data_out <= rom_array(17870);
		when "0100010111001111" => data_out <= rom_array(17871);
		when "0100010111010000" => data_out <= rom_array(17872);
		when "0100010111010001" => data_out <= rom_array(17873);
		when "0100010111010010" => data_out <= rom_array(17874);
		when "0100010111010011" => data_out <= rom_array(17875);
		when "0100010111010100" => data_out <= rom_array(17876);
		when "0100010111010101" => data_out <= rom_array(17877);
		when "0100010111010110" => data_out <= rom_array(17878);
		when "0100010111010111" => data_out <= rom_array(17879);
		when "0100010111011000" => data_out <= rom_array(17880);
		when "0100010111011001" => data_out <= rom_array(17881);
		when "0100010111011010" => data_out <= rom_array(17882);
		when "0100010111011011" => data_out <= rom_array(17883);
		when "0100010111011100" => data_out <= rom_array(17884);
		when "0100010111011101" => data_out <= rom_array(17885);
		when "0100010111011110" => data_out <= rom_array(17886);
		when "0100010111011111" => data_out <= rom_array(17887);
		when "0100010111100000" => data_out <= rom_array(17888);
		when "0100010111100001" => data_out <= rom_array(17889);
		when "0100010111100010" => data_out <= rom_array(17890);
		when "0100010111100011" => data_out <= rom_array(17891);
		when "0100010111100100" => data_out <= rom_array(17892);
		when "0100010111100101" => data_out <= rom_array(17893);
		when "0100010111100110" => data_out <= rom_array(17894);
		when "0100010111100111" => data_out <= rom_array(17895);
		when "0100010111101000" => data_out <= rom_array(17896);
		when "0100010111101001" => data_out <= rom_array(17897);
		when "0100010111101010" => data_out <= rom_array(17898);
		when "0100010111101011" => data_out <= rom_array(17899);
		when "0100010111101100" => data_out <= rom_array(17900);
		when "0100010111101101" => data_out <= rom_array(17901);
		when "0100010111101110" => data_out <= rom_array(17902);
		when "0100010111101111" => data_out <= rom_array(17903);
		when "0100010111110000" => data_out <= rom_array(17904);
		when "0100010111110001" => data_out <= rom_array(17905);
		when "0100010111110010" => data_out <= rom_array(17906);
		when "0100010111110011" => data_out <= rom_array(17907);
		when "0100010111110100" => data_out <= rom_array(17908);
		when "0100010111110101" => data_out <= rom_array(17909);
		when "0100010111110110" => data_out <= rom_array(17910);
		when "0100010111110111" => data_out <= rom_array(17911);
		when "0100010111111000" => data_out <= rom_array(17912);
		when "0100010111111001" => data_out <= rom_array(17913);
		when "0100010111111010" => data_out <= rom_array(17914);
		when "0100010111111011" => data_out <= rom_array(17915);
		when "0100010111111100" => data_out <= rom_array(17916);
		when "0100010111111101" => data_out <= rom_array(17917);
		when "0100010111111110" => data_out <= rom_array(17918);
		when "0100010111111111" => data_out <= rom_array(17919);
		when "0100011000000000" => data_out <= rom_array(17920);
		when "0100011000000001" => data_out <= rom_array(17921);
		when "0100011000000010" => data_out <= rom_array(17922);
		when "0100011000000011" => data_out <= rom_array(17923);
		when "0100011000000100" => data_out <= rom_array(17924);
		when "0100011000000101" => data_out <= rom_array(17925);
		when "0100011000000110" => data_out <= rom_array(17926);
		when "0100011000000111" => data_out <= rom_array(17927);
		when "0100011000001000" => data_out <= rom_array(17928);
		when "0100011000001001" => data_out <= rom_array(17929);
		when "0100011000001010" => data_out <= rom_array(17930);
		when "0100011000001011" => data_out <= rom_array(17931);
		when "0100011000001100" => data_out <= rom_array(17932);
		when "0100011000001101" => data_out <= rom_array(17933);
		when "0100011000001110" => data_out <= rom_array(17934);
		when "0100011000001111" => data_out <= rom_array(17935);
		when "0100011000010000" => data_out <= rom_array(17936);
		when "0100011000010001" => data_out <= rom_array(17937);
		when "0100011000010010" => data_out <= rom_array(17938);
		when "0100011000010011" => data_out <= rom_array(17939);
		when "0100011000010100" => data_out <= rom_array(17940);
		when "0100011000010101" => data_out <= rom_array(17941);
		when "0100011000010110" => data_out <= rom_array(17942);
		when "0100011000010111" => data_out <= rom_array(17943);
		when "0100011000011000" => data_out <= rom_array(17944);
		when "0100011000011001" => data_out <= rom_array(17945);
		when "0100011000011010" => data_out <= rom_array(17946);
		when "0100011000011011" => data_out <= rom_array(17947);
		when "0100011000011100" => data_out <= rom_array(17948);
		when "0100011000011101" => data_out <= rom_array(17949);
		when "0100011000011110" => data_out <= rom_array(17950);
		when "0100011000011111" => data_out <= rom_array(17951);
		when "0100011000100000" => data_out <= rom_array(17952);
		when "0100011000100001" => data_out <= rom_array(17953);
		when "0100011000100010" => data_out <= rom_array(17954);
		when "0100011000100011" => data_out <= rom_array(17955);
		when "0100011000100100" => data_out <= rom_array(17956);
		when "0100011000100101" => data_out <= rom_array(17957);
		when "0100011000100110" => data_out <= rom_array(17958);
		when "0100011000100111" => data_out <= rom_array(17959);
		when "0100011000101000" => data_out <= rom_array(17960);
		when "0100011000101001" => data_out <= rom_array(17961);
		when "0100011000101010" => data_out <= rom_array(17962);
		when "0100011000101011" => data_out <= rom_array(17963);
		when "0100011000101100" => data_out <= rom_array(17964);
		when "0100011000101101" => data_out <= rom_array(17965);
		when "0100011000101110" => data_out <= rom_array(17966);
		when "0100011000101111" => data_out <= rom_array(17967);
		when "0100011000110000" => data_out <= rom_array(17968);
		when "0100011000110001" => data_out <= rom_array(17969);
		when "0100011000110010" => data_out <= rom_array(17970);
		when "0100011000110011" => data_out <= rom_array(17971);
		when "0100011000110100" => data_out <= rom_array(17972);
		when "0100011000110101" => data_out <= rom_array(17973);
		when "0100011000110110" => data_out <= rom_array(17974);
		when "0100011000110111" => data_out <= rom_array(17975);
		when "0100011000111000" => data_out <= rom_array(17976);
		when "0100011000111001" => data_out <= rom_array(17977);
		when "0100011000111010" => data_out <= rom_array(17978);
		when "0100011000111011" => data_out <= rom_array(17979);
		when "0100011000111100" => data_out <= rom_array(17980);
		when "0100011000111101" => data_out <= rom_array(17981);
		when "0100011000111110" => data_out <= rom_array(17982);
		when "0100011000111111" => data_out <= rom_array(17983);
		when "0100011001000000" => data_out <= rom_array(17984);
		when "0100011001000001" => data_out <= rom_array(17985);
		when "0100011001000010" => data_out <= rom_array(17986);
		when "0100011001000011" => data_out <= rom_array(17987);
		when "0100011001000100" => data_out <= rom_array(17988);
		when "0100011001000101" => data_out <= rom_array(17989);
		when "0100011001000110" => data_out <= rom_array(17990);
		when "0100011001000111" => data_out <= rom_array(17991);
		when "0100011001001000" => data_out <= rom_array(17992);
		when "0100011001001001" => data_out <= rom_array(17993);
		when "0100011001001010" => data_out <= rom_array(17994);
		when "0100011001001011" => data_out <= rom_array(17995);
		when "0100011001001100" => data_out <= rom_array(17996);
		when "0100011001001101" => data_out <= rom_array(17997);
		when "0100011001001110" => data_out <= rom_array(17998);
		when "0100011001001111" => data_out <= rom_array(17999);
		when "0100011001010000" => data_out <= rom_array(18000);
		when "0100011001010001" => data_out <= rom_array(18001);
		when "0100011001010010" => data_out <= rom_array(18002);
		when "0100011001010011" => data_out <= rom_array(18003);
		when "0100011001010100" => data_out <= rom_array(18004);
		when "0100011001010101" => data_out <= rom_array(18005);
		when "0100011001010110" => data_out <= rom_array(18006);
		when "0100011001010111" => data_out <= rom_array(18007);
		when "0100011001011000" => data_out <= rom_array(18008);
		when "0100011001011001" => data_out <= rom_array(18009);
		when "0100011001011010" => data_out <= rom_array(18010);
		when "0100011001011011" => data_out <= rom_array(18011);
		when "0100011001011100" => data_out <= rom_array(18012);
		when "0100011001011101" => data_out <= rom_array(18013);
		when "0100011001011110" => data_out <= rom_array(18014);
		when "0100011001011111" => data_out <= rom_array(18015);
		when "0100011001100000" => data_out <= rom_array(18016);
		when "0100011001100001" => data_out <= rom_array(18017);
		when "0100011001100010" => data_out <= rom_array(18018);
		when "0100011001100011" => data_out <= rom_array(18019);
		when "0100011001100100" => data_out <= rom_array(18020);
		when "0100011001100101" => data_out <= rom_array(18021);
		when "0100011001100110" => data_out <= rom_array(18022);
		when "0100011001100111" => data_out <= rom_array(18023);
		when "0100011001101000" => data_out <= rom_array(18024);
		when "0100011001101001" => data_out <= rom_array(18025);
		when "0100011001101010" => data_out <= rom_array(18026);
		when "0100011001101011" => data_out <= rom_array(18027);
		when "0100011001101100" => data_out <= rom_array(18028);
		when "0100011001101101" => data_out <= rom_array(18029);
		when "0100011001101110" => data_out <= rom_array(18030);
		when "0100011001101111" => data_out <= rom_array(18031);
		when "0100011001110000" => data_out <= rom_array(18032);
		when "0100011001110001" => data_out <= rom_array(18033);
		when "0100011001110010" => data_out <= rom_array(18034);
		when "0100011001110011" => data_out <= rom_array(18035);
		when "0100011001110100" => data_out <= rom_array(18036);
		when "0100011001110101" => data_out <= rom_array(18037);
		when "0100011001110110" => data_out <= rom_array(18038);
		when "0100011001110111" => data_out <= rom_array(18039);
		when "0100011001111000" => data_out <= rom_array(18040);
		when "0100011001111001" => data_out <= rom_array(18041);
		when "0100011001111010" => data_out <= rom_array(18042);
		when "0100011001111011" => data_out <= rom_array(18043);
		when "0100011001111100" => data_out <= rom_array(18044);
		when "0100011001111101" => data_out <= rom_array(18045);
		when "0100011001111110" => data_out <= rom_array(18046);
		when "0100011001111111" => data_out <= rom_array(18047);
		when "0100011010000000" => data_out <= rom_array(18048);
		when "0100011010000001" => data_out <= rom_array(18049);
		when "0100011010000010" => data_out <= rom_array(18050);
		when "0100011010000011" => data_out <= rom_array(18051);
		when "0100011010000100" => data_out <= rom_array(18052);
		when "0100011010000101" => data_out <= rom_array(18053);
		when "0100011010000110" => data_out <= rom_array(18054);
		when "0100011010000111" => data_out <= rom_array(18055);
		when "0100011010001000" => data_out <= rom_array(18056);
		when "0100011010001001" => data_out <= rom_array(18057);
		when "0100011010001010" => data_out <= rom_array(18058);
		when "0100011010001011" => data_out <= rom_array(18059);
		when "0100011010001100" => data_out <= rom_array(18060);
		when "0100011010001101" => data_out <= rom_array(18061);
		when "0100011010001110" => data_out <= rom_array(18062);
		when "0100011010001111" => data_out <= rom_array(18063);
		when "0100011010010000" => data_out <= rom_array(18064);
		when "0100011010010001" => data_out <= rom_array(18065);
		when "0100011010010010" => data_out <= rom_array(18066);
		when "0100011010010011" => data_out <= rom_array(18067);
		when "0100011010010100" => data_out <= rom_array(18068);
		when "0100011010010101" => data_out <= rom_array(18069);
		when "0100011010010110" => data_out <= rom_array(18070);
		when "0100011010010111" => data_out <= rom_array(18071);
		when "0100011010011000" => data_out <= rom_array(18072);
		when "0100011010011001" => data_out <= rom_array(18073);
		when "0100011010011010" => data_out <= rom_array(18074);
		when "0100011010011011" => data_out <= rom_array(18075);
		when "0100011010011100" => data_out <= rom_array(18076);
		when "0100011010011101" => data_out <= rom_array(18077);
		when "0100011010011110" => data_out <= rom_array(18078);
		when "0100011010011111" => data_out <= rom_array(18079);
		when "0100011010100000" => data_out <= rom_array(18080);
		when "0100011010100001" => data_out <= rom_array(18081);
		when "0100011010100010" => data_out <= rom_array(18082);
		when "0100011010100011" => data_out <= rom_array(18083);
		when "0100011010100100" => data_out <= rom_array(18084);
		when "0100011010100101" => data_out <= rom_array(18085);
		when "0100011010100110" => data_out <= rom_array(18086);
		when "0100011010100111" => data_out <= rom_array(18087);
		when "0100011010101000" => data_out <= rom_array(18088);
		when "0100011010101001" => data_out <= rom_array(18089);
		when "0100011010101010" => data_out <= rom_array(18090);
		when "0100011010101011" => data_out <= rom_array(18091);
		when "0100011010101100" => data_out <= rom_array(18092);
		when "0100011010101101" => data_out <= rom_array(18093);
		when "0100011010101110" => data_out <= rom_array(18094);
		when "0100011010101111" => data_out <= rom_array(18095);
		when "0100011010110000" => data_out <= rom_array(18096);
		when "0100011010110001" => data_out <= rom_array(18097);
		when "0100011010110010" => data_out <= rom_array(18098);
		when "0100011010110011" => data_out <= rom_array(18099);
		when "0100011010110100" => data_out <= rom_array(18100);
		when "0100011010110101" => data_out <= rom_array(18101);
		when "0100011010110110" => data_out <= rom_array(18102);
		when "0100011010110111" => data_out <= rom_array(18103);
		when "0100011010111000" => data_out <= rom_array(18104);
		when "0100011010111001" => data_out <= rom_array(18105);
		when "0100011010111010" => data_out <= rom_array(18106);
		when "0100011010111011" => data_out <= rom_array(18107);
		when "0100011010111100" => data_out <= rom_array(18108);
		when "0100011010111101" => data_out <= rom_array(18109);
		when "0100011010111110" => data_out <= rom_array(18110);
		when "0100011010111111" => data_out <= rom_array(18111);
		when "0100011011000000" => data_out <= rom_array(18112);
		when "0100011011000001" => data_out <= rom_array(18113);
		when "0100011011000010" => data_out <= rom_array(18114);
		when "0100011011000011" => data_out <= rom_array(18115);
		when "0100011011000100" => data_out <= rom_array(18116);
		when "0100011011000101" => data_out <= rom_array(18117);
		when "0100011011000110" => data_out <= rom_array(18118);
		when "0100011011000111" => data_out <= rom_array(18119);
		when "0100011011001000" => data_out <= rom_array(18120);
		when "0100011011001001" => data_out <= rom_array(18121);
		when "0100011011001010" => data_out <= rom_array(18122);
		when "0100011011001011" => data_out <= rom_array(18123);
		when "0100011011001100" => data_out <= rom_array(18124);
		when "0100011011001101" => data_out <= rom_array(18125);
		when "0100011011001110" => data_out <= rom_array(18126);
		when "0100011011001111" => data_out <= rom_array(18127);
		when "0100011011010000" => data_out <= rom_array(18128);
		when "0100011011010001" => data_out <= rom_array(18129);
		when "0100011011010010" => data_out <= rom_array(18130);
		when "0100011011010011" => data_out <= rom_array(18131);
		when "0100011011010100" => data_out <= rom_array(18132);
		when "0100011011010101" => data_out <= rom_array(18133);
		when "0100011011010110" => data_out <= rom_array(18134);
		when "0100011011010111" => data_out <= rom_array(18135);
		when "0100011011011000" => data_out <= rom_array(18136);
		when "0100011011011001" => data_out <= rom_array(18137);
		when "0100011011011010" => data_out <= rom_array(18138);
		when "0100011011011011" => data_out <= rom_array(18139);
		when "0100011011011100" => data_out <= rom_array(18140);
		when "0100011011011101" => data_out <= rom_array(18141);
		when "0100011011011110" => data_out <= rom_array(18142);
		when "0100011011011111" => data_out <= rom_array(18143);
		when "0100011011100000" => data_out <= rom_array(18144);
		when "0100011011100001" => data_out <= rom_array(18145);
		when "0100011011100010" => data_out <= rom_array(18146);
		when "0100011011100011" => data_out <= rom_array(18147);
		when "0100011011100100" => data_out <= rom_array(18148);
		when "0100011011100101" => data_out <= rom_array(18149);
		when "0100011011100110" => data_out <= rom_array(18150);
		when "0100011011100111" => data_out <= rom_array(18151);
		when "0100011011101000" => data_out <= rom_array(18152);
		when "0100011011101001" => data_out <= rom_array(18153);
		when "0100011011101010" => data_out <= rom_array(18154);
		when "0100011011101011" => data_out <= rom_array(18155);
		when "0100011011101100" => data_out <= rom_array(18156);
		when "0100011011101101" => data_out <= rom_array(18157);
		when "0100011011101110" => data_out <= rom_array(18158);
		when "0100011011101111" => data_out <= rom_array(18159);
		when "0100011011110000" => data_out <= rom_array(18160);
		when "0100011011110001" => data_out <= rom_array(18161);
		when "0100011011110010" => data_out <= rom_array(18162);
		when "0100011011110011" => data_out <= rom_array(18163);
		when "0100011011110100" => data_out <= rom_array(18164);
		when "0100011011110101" => data_out <= rom_array(18165);
		when "0100011011110110" => data_out <= rom_array(18166);
		when "0100011011110111" => data_out <= rom_array(18167);
		when "0100011011111000" => data_out <= rom_array(18168);
		when "0100011011111001" => data_out <= rom_array(18169);
		when "0100011011111010" => data_out <= rom_array(18170);
		when "0100011011111011" => data_out <= rom_array(18171);
		when "0100011011111100" => data_out <= rom_array(18172);
		when "0100011011111101" => data_out <= rom_array(18173);
		when "0100011011111110" => data_out <= rom_array(18174);
		when "0100011011111111" => data_out <= rom_array(18175);
		when "0100011100000000" => data_out <= rom_array(18176);
		when "0100011100000001" => data_out <= rom_array(18177);
		when "0100011100000010" => data_out <= rom_array(18178);
		when "0100011100000011" => data_out <= rom_array(18179);
		when "0100011100000100" => data_out <= rom_array(18180);
		when "0100011100000101" => data_out <= rom_array(18181);
		when "0100011100000110" => data_out <= rom_array(18182);
		when "0100011100000111" => data_out <= rom_array(18183);
		when "0100011100001000" => data_out <= rom_array(18184);
		when "0100011100001001" => data_out <= rom_array(18185);
		when "0100011100001010" => data_out <= rom_array(18186);
		when "0100011100001011" => data_out <= rom_array(18187);
		when "0100011100001100" => data_out <= rom_array(18188);
		when "0100011100001101" => data_out <= rom_array(18189);
		when "0100011100001110" => data_out <= rom_array(18190);
		when "0100011100001111" => data_out <= rom_array(18191);
		when "0100011100010000" => data_out <= rom_array(18192);
		when "0100011100010001" => data_out <= rom_array(18193);
		when "0100011100010010" => data_out <= rom_array(18194);
		when "0100011100010011" => data_out <= rom_array(18195);
		when "0100011100010100" => data_out <= rom_array(18196);
		when "0100011100010101" => data_out <= rom_array(18197);
		when "0100011100010110" => data_out <= rom_array(18198);
		when "0100011100010111" => data_out <= rom_array(18199);
		when "0100011100011000" => data_out <= rom_array(18200);
		when "0100011100011001" => data_out <= rom_array(18201);
		when "0100011100011010" => data_out <= rom_array(18202);
		when "0100011100011011" => data_out <= rom_array(18203);
		when "0100011100011100" => data_out <= rom_array(18204);
		when "0100011100011101" => data_out <= rom_array(18205);
		when "0100011100011110" => data_out <= rom_array(18206);
		when "0100011100011111" => data_out <= rom_array(18207);
		when "0100011100100000" => data_out <= rom_array(18208);
		when "0100011100100001" => data_out <= rom_array(18209);
		when "0100011100100010" => data_out <= rom_array(18210);
		when "0100011100100011" => data_out <= rom_array(18211);
		when "0100011100100100" => data_out <= rom_array(18212);
		when "0100011100100101" => data_out <= rom_array(18213);
		when "0100011100100110" => data_out <= rom_array(18214);
		when "0100011100100111" => data_out <= rom_array(18215);
		when "0100011100101000" => data_out <= rom_array(18216);
		when "0100011100101001" => data_out <= rom_array(18217);
		when "0100011100101010" => data_out <= rom_array(18218);
		when "0100011100101011" => data_out <= rom_array(18219);
		when "0100011100101100" => data_out <= rom_array(18220);
		when "0100011100101101" => data_out <= rom_array(18221);
		when "0100011100101110" => data_out <= rom_array(18222);
		when "0100011100101111" => data_out <= rom_array(18223);
		when "0100011100110000" => data_out <= rom_array(18224);
		when "0100011100110001" => data_out <= rom_array(18225);
		when "0100011100110010" => data_out <= rom_array(18226);
		when "0100011100110011" => data_out <= rom_array(18227);
		when "0100011100110100" => data_out <= rom_array(18228);
		when "0100011100110101" => data_out <= rom_array(18229);
		when "0100011100110110" => data_out <= rom_array(18230);
		when "0100011100110111" => data_out <= rom_array(18231);
		when "0100011100111000" => data_out <= rom_array(18232);
		when "0100011100111001" => data_out <= rom_array(18233);
		when "0100011100111010" => data_out <= rom_array(18234);
		when "0100011100111011" => data_out <= rom_array(18235);
		when "0100011100111100" => data_out <= rom_array(18236);
		when "0100011100111101" => data_out <= rom_array(18237);
		when "0100011100111110" => data_out <= rom_array(18238);
		when "0100011100111111" => data_out <= rom_array(18239);
		when "0100011101000000" => data_out <= rom_array(18240);
		when "0100011101000001" => data_out <= rom_array(18241);
		when "0100011101000010" => data_out <= rom_array(18242);
		when "0100011101000011" => data_out <= rom_array(18243);
		when "0100011101000100" => data_out <= rom_array(18244);
		when "0100011101000101" => data_out <= rom_array(18245);
		when "0100011101000110" => data_out <= rom_array(18246);
		when "0100011101000111" => data_out <= rom_array(18247);
		when "0100011101001000" => data_out <= rom_array(18248);
		when "0100011101001001" => data_out <= rom_array(18249);
		when "0100011101001010" => data_out <= rom_array(18250);
		when "0100011101001011" => data_out <= rom_array(18251);
		when "0100011101001100" => data_out <= rom_array(18252);
		when "0100011101001101" => data_out <= rom_array(18253);
		when "0100011101001110" => data_out <= rom_array(18254);
		when "0100011101001111" => data_out <= rom_array(18255);
		when "0100011101010000" => data_out <= rom_array(18256);
		when "0100011101010001" => data_out <= rom_array(18257);
		when "0100011101010010" => data_out <= rom_array(18258);
		when "0100011101010011" => data_out <= rom_array(18259);
		when "0100011101010100" => data_out <= rom_array(18260);
		when "0100011101010101" => data_out <= rom_array(18261);
		when "0100011101010110" => data_out <= rom_array(18262);
		when "0100011101010111" => data_out <= rom_array(18263);
		when "0100011101011000" => data_out <= rom_array(18264);
		when "0100011101011001" => data_out <= rom_array(18265);
		when "0100011101011010" => data_out <= rom_array(18266);
		when "0100011101011011" => data_out <= rom_array(18267);
		when "0100011101011100" => data_out <= rom_array(18268);
		when "0100011101011101" => data_out <= rom_array(18269);
		when "0100011101011110" => data_out <= rom_array(18270);
		when "0100011101011111" => data_out <= rom_array(18271);
		when "0100011101100000" => data_out <= rom_array(18272);
		when "0100011101100001" => data_out <= rom_array(18273);
		when "0100011101100010" => data_out <= rom_array(18274);
		when "0100011101100011" => data_out <= rom_array(18275);
		when "0100011101100100" => data_out <= rom_array(18276);
		when "0100011101100101" => data_out <= rom_array(18277);
		when "0100011101100110" => data_out <= rom_array(18278);
		when "0100011101100111" => data_out <= rom_array(18279);
		when "0100011101101000" => data_out <= rom_array(18280);
		when "0100011101101001" => data_out <= rom_array(18281);
		when "0100011101101010" => data_out <= rom_array(18282);
		when "0100011101101011" => data_out <= rom_array(18283);
		when "0100011101101100" => data_out <= rom_array(18284);
		when "0100011101101101" => data_out <= rom_array(18285);
		when "0100011101101110" => data_out <= rom_array(18286);
		when "0100011101101111" => data_out <= rom_array(18287);
		when "0100011101110000" => data_out <= rom_array(18288);
		when "0100011101110001" => data_out <= rom_array(18289);
		when "0100011101110010" => data_out <= rom_array(18290);
		when "0100011101110011" => data_out <= rom_array(18291);
		when "0100011101110100" => data_out <= rom_array(18292);
		when "0100011101110101" => data_out <= rom_array(18293);
		when "0100011101110110" => data_out <= rom_array(18294);
		when "0100011101110111" => data_out <= rom_array(18295);
		when "0100011101111000" => data_out <= rom_array(18296);
		when "0100011101111001" => data_out <= rom_array(18297);
		when "0100011101111010" => data_out <= rom_array(18298);
		when "0100011101111011" => data_out <= rom_array(18299);
		when "0100011101111100" => data_out <= rom_array(18300);
		when "0100011101111101" => data_out <= rom_array(18301);
		when "0100011101111110" => data_out <= rom_array(18302);
		when "0100011101111111" => data_out <= rom_array(18303);
		when "0100011110000000" => data_out <= rom_array(18304);
		when "0100011110000001" => data_out <= rom_array(18305);
		when "0100011110000010" => data_out <= rom_array(18306);
		when "0100011110000011" => data_out <= rom_array(18307);
		when "0100011110000100" => data_out <= rom_array(18308);
		when "0100011110000101" => data_out <= rom_array(18309);
		when "0100011110000110" => data_out <= rom_array(18310);
		when "0100011110000111" => data_out <= rom_array(18311);
		when "0100011110001000" => data_out <= rom_array(18312);
		when "0100011110001001" => data_out <= rom_array(18313);
		when "0100011110001010" => data_out <= rom_array(18314);
		when "0100011110001011" => data_out <= rom_array(18315);
		when "0100011110001100" => data_out <= rom_array(18316);
		when "0100011110001101" => data_out <= rom_array(18317);
		when "0100011110001110" => data_out <= rom_array(18318);
		when "0100011110001111" => data_out <= rom_array(18319);
		when "0100011110010000" => data_out <= rom_array(18320);
		when "0100011110010001" => data_out <= rom_array(18321);
		when "0100011110010010" => data_out <= rom_array(18322);
		when "0100011110010011" => data_out <= rom_array(18323);
		when "0100011110010100" => data_out <= rom_array(18324);
		when "0100011110010101" => data_out <= rom_array(18325);
		when "0100011110010110" => data_out <= rom_array(18326);
		when "0100011110010111" => data_out <= rom_array(18327);
		when "0100011110011000" => data_out <= rom_array(18328);
		when "0100011110011001" => data_out <= rom_array(18329);
		when "0100011110011010" => data_out <= rom_array(18330);
		when "0100011110011011" => data_out <= rom_array(18331);
		when "0100011110011100" => data_out <= rom_array(18332);
		when "0100011110011101" => data_out <= rom_array(18333);
		when "0100011110011110" => data_out <= rom_array(18334);
		when "0100011110011111" => data_out <= rom_array(18335);
		when "0100011110100000" => data_out <= rom_array(18336);
		when "0100011110100001" => data_out <= rom_array(18337);
		when "0100011110100010" => data_out <= rom_array(18338);
		when "0100011110100011" => data_out <= rom_array(18339);
		when "0100011110100100" => data_out <= rom_array(18340);
		when "0100011110100101" => data_out <= rom_array(18341);
		when "0100011110100110" => data_out <= rom_array(18342);
		when "0100011110100111" => data_out <= rom_array(18343);
		when "0100011110101000" => data_out <= rom_array(18344);
		when "0100011110101001" => data_out <= rom_array(18345);
		when "0100011110101010" => data_out <= rom_array(18346);
		when "0100011110101011" => data_out <= rom_array(18347);
		when "0100011110101100" => data_out <= rom_array(18348);
		when "0100011110101101" => data_out <= rom_array(18349);
		when "0100011110101110" => data_out <= rom_array(18350);
		when "0100011110101111" => data_out <= rom_array(18351);
		when "0100011110110000" => data_out <= rom_array(18352);
		when "0100011110110001" => data_out <= rom_array(18353);
		when "0100011110110010" => data_out <= rom_array(18354);
		when "0100011110110011" => data_out <= rom_array(18355);
		when "0100011110110100" => data_out <= rom_array(18356);
		when "0100011110110101" => data_out <= rom_array(18357);
		when "0100011110110110" => data_out <= rom_array(18358);
		when "0100011110110111" => data_out <= rom_array(18359);
		when "0100011110111000" => data_out <= rom_array(18360);
		when "0100011110111001" => data_out <= rom_array(18361);
		when "0100011110111010" => data_out <= rom_array(18362);
		when "0100011110111011" => data_out <= rom_array(18363);
		when "0100011110111100" => data_out <= rom_array(18364);
		when "0100011110111101" => data_out <= rom_array(18365);
		when "0100011110111110" => data_out <= rom_array(18366);
		when "0100011110111111" => data_out <= rom_array(18367);
		when "0100011111000000" => data_out <= rom_array(18368);
		when "0100011111000001" => data_out <= rom_array(18369);
		when "0100011111000010" => data_out <= rom_array(18370);
		when "0100011111000011" => data_out <= rom_array(18371);
		when "0100011111000100" => data_out <= rom_array(18372);
		when "0100011111000101" => data_out <= rom_array(18373);
		when "0100011111000110" => data_out <= rom_array(18374);
		when "0100011111000111" => data_out <= rom_array(18375);
		when "0100011111001000" => data_out <= rom_array(18376);
		when "0100011111001001" => data_out <= rom_array(18377);
		when "0100011111001010" => data_out <= rom_array(18378);
		when "0100011111001011" => data_out <= rom_array(18379);
		when "0100011111001100" => data_out <= rom_array(18380);
		when "0100011111001101" => data_out <= rom_array(18381);
		when "0100011111001110" => data_out <= rom_array(18382);
		when "0100011111001111" => data_out <= rom_array(18383);
		when "0100011111010000" => data_out <= rom_array(18384);
		when "0100011111010001" => data_out <= rom_array(18385);
		when "0100011111010010" => data_out <= rom_array(18386);
		when "0100011111010011" => data_out <= rom_array(18387);
		when "0100011111010100" => data_out <= rom_array(18388);
		when "0100011111010101" => data_out <= rom_array(18389);
		when "0100011111010110" => data_out <= rom_array(18390);
		when "0100011111010111" => data_out <= rom_array(18391);
		when "0100011111011000" => data_out <= rom_array(18392);
		when "0100011111011001" => data_out <= rom_array(18393);
		when "0100011111011010" => data_out <= rom_array(18394);
		when "0100011111011011" => data_out <= rom_array(18395);
		when "0100011111011100" => data_out <= rom_array(18396);
		when "0100011111011101" => data_out <= rom_array(18397);
		when "0100011111011110" => data_out <= rom_array(18398);
		when "0100011111011111" => data_out <= rom_array(18399);
		when "0100011111100000" => data_out <= rom_array(18400);
		when "0100011111100001" => data_out <= rom_array(18401);
		when "0100011111100010" => data_out <= rom_array(18402);
		when "0100011111100011" => data_out <= rom_array(18403);
		when "0100011111100100" => data_out <= rom_array(18404);
		when "0100011111100101" => data_out <= rom_array(18405);
		when "0100011111100110" => data_out <= rom_array(18406);
		when "0100011111100111" => data_out <= rom_array(18407);
		when "0100011111101000" => data_out <= rom_array(18408);
		when "0100011111101001" => data_out <= rom_array(18409);
		when "0100011111101010" => data_out <= rom_array(18410);
		when "0100011111101011" => data_out <= rom_array(18411);
		when "0100011111101100" => data_out <= rom_array(18412);
		when "0100011111101101" => data_out <= rom_array(18413);
		when "0100011111101110" => data_out <= rom_array(18414);
		when "0100011111101111" => data_out <= rom_array(18415);
		when "0100011111110000" => data_out <= rom_array(18416);
		when "0100011111110001" => data_out <= rom_array(18417);
		when "0100011111110010" => data_out <= rom_array(18418);
		when "0100011111110011" => data_out <= rom_array(18419);
		when "0100011111110100" => data_out <= rom_array(18420);
		when "0100011111110101" => data_out <= rom_array(18421);
		when "0100011111110110" => data_out <= rom_array(18422);
		when "0100011111110111" => data_out <= rom_array(18423);
		when "0100011111111000" => data_out <= rom_array(18424);
		when "0100011111111001" => data_out <= rom_array(18425);
		when "0100011111111010" => data_out <= rom_array(18426);
		when "0100011111111011" => data_out <= rom_array(18427);
		when "0100011111111100" => data_out <= rom_array(18428);
		when "0100011111111101" => data_out <= rom_array(18429);
		when "0100011111111110" => data_out <= rom_array(18430);
		when "0100011111111111" => data_out <= rom_array(18431);
		when "0100100000000000" => data_out <= rom_array(18432);
		when "0100100000000001" => data_out <= rom_array(18433);
		when "0100100000000010" => data_out <= rom_array(18434);
		when "0100100000000011" => data_out <= rom_array(18435);
		when "0100100000000100" => data_out <= rom_array(18436);
		when "0100100000000101" => data_out <= rom_array(18437);
		when "0100100000000110" => data_out <= rom_array(18438);
		when "0100100000000111" => data_out <= rom_array(18439);
		when "0100100000001000" => data_out <= rom_array(18440);
		when "0100100000001001" => data_out <= rom_array(18441);
		when "0100100000001010" => data_out <= rom_array(18442);
		when "0100100000001011" => data_out <= rom_array(18443);
		when "0100100000001100" => data_out <= rom_array(18444);
		when "0100100000001101" => data_out <= rom_array(18445);
		when "0100100000001110" => data_out <= rom_array(18446);
		when "0100100000001111" => data_out <= rom_array(18447);
		when "0100100000010000" => data_out <= rom_array(18448);
		when "0100100000010001" => data_out <= rom_array(18449);
		when "0100100000010010" => data_out <= rom_array(18450);
		when "0100100000010011" => data_out <= rom_array(18451);
		when "0100100000010100" => data_out <= rom_array(18452);
		when "0100100000010101" => data_out <= rom_array(18453);
		when "0100100000010110" => data_out <= rom_array(18454);
		when "0100100000010111" => data_out <= rom_array(18455);
		when "0100100000011000" => data_out <= rom_array(18456);
		when "0100100000011001" => data_out <= rom_array(18457);
		when "0100100000011010" => data_out <= rom_array(18458);
		when "0100100000011011" => data_out <= rom_array(18459);
		when "0100100000011100" => data_out <= rom_array(18460);
		when "0100100000011101" => data_out <= rom_array(18461);
		when "0100100000011110" => data_out <= rom_array(18462);
		when "0100100000011111" => data_out <= rom_array(18463);
		when "0100100000100000" => data_out <= rom_array(18464);
		when "0100100000100001" => data_out <= rom_array(18465);
		when "0100100000100010" => data_out <= rom_array(18466);
		when "0100100000100011" => data_out <= rom_array(18467);
		when "0100100000100100" => data_out <= rom_array(18468);
		when "0100100000100101" => data_out <= rom_array(18469);
		when "0100100000100110" => data_out <= rom_array(18470);
		when "0100100000100111" => data_out <= rom_array(18471);
		when "0100100000101000" => data_out <= rom_array(18472);
		when "0100100000101001" => data_out <= rom_array(18473);
		when "0100100000101010" => data_out <= rom_array(18474);
		when "0100100000101011" => data_out <= rom_array(18475);
		when "0100100000101100" => data_out <= rom_array(18476);
		when "0100100000101101" => data_out <= rom_array(18477);
		when "0100100000101110" => data_out <= rom_array(18478);
		when "0100100000101111" => data_out <= rom_array(18479);
		when "0100100000110000" => data_out <= rom_array(18480);
		when "0100100000110001" => data_out <= rom_array(18481);
		when "0100100000110010" => data_out <= rom_array(18482);
		when "0100100000110011" => data_out <= rom_array(18483);
		when "0100100000110100" => data_out <= rom_array(18484);
		when "0100100000110101" => data_out <= rom_array(18485);
		when "0100100000110110" => data_out <= rom_array(18486);
		when "0100100000110111" => data_out <= rom_array(18487);
		when "0100100000111000" => data_out <= rom_array(18488);
		when "0100100000111001" => data_out <= rom_array(18489);
		when "0100100000111010" => data_out <= rom_array(18490);
		when "0100100000111011" => data_out <= rom_array(18491);
		when "0100100000111100" => data_out <= rom_array(18492);
		when "0100100000111101" => data_out <= rom_array(18493);
		when "0100100000111110" => data_out <= rom_array(18494);
		when "0100100000111111" => data_out <= rom_array(18495);
		when "0100100001000000" => data_out <= rom_array(18496);
		when "0100100001000001" => data_out <= rom_array(18497);
		when "0100100001000010" => data_out <= rom_array(18498);
		when "0100100001000011" => data_out <= rom_array(18499);
		when "0100100001000100" => data_out <= rom_array(18500);
		when "0100100001000101" => data_out <= rom_array(18501);
		when "0100100001000110" => data_out <= rom_array(18502);
		when "0100100001000111" => data_out <= rom_array(18503);
		when "0100100001001000" => data_out <= rom_array(18504);
		when "0100100001001001" => data_out <= rom_array(18505);
		when "0100100001001010" => data_out <= rom_array(18506);
		when "0100100001001011" => data_out <= rom_array(18507);
		when "0100100001001100" => data_out <= rom_array(18508);
		when "0100100001001101" => data_out <= rom_array(18509);
		when "0100100001001110" => data_out <= rom_array(18510);
		when "0100100001001111" => data_out <= rom_array(18511);
		when "0100100001010000" => data_out <= rom_array(18512);
		when "0100100001010001" => data_out <= rom_array(18513);
		when "0100100001010010" => data_out <= rom_array(18514);
		when "0100100001010011" => data_out <= rom_array(18515);
		when "0100100001010100" => data_out <= rom_array(18516);
		when "0100100001010101" => data_out <= rom_array(18517);
		when "0100100001010110" => data_out <= rom_array(18518);
		when "0100100001010111" => data_out <= rom_array(18519);
		when "0100100001011000" => data_out <= rom_array(18520);
		when "0100100001011001" => data_out <= rom_array(18521);
		when "0100100001011010" => data_out <= rom_array(18522);
		when "0100100001011011" => data_out <= rom_array(18523);
		when "0100100001011100" => data_out <= rom_array(18524);
		when "0100100001011101" => data_out <= rom_array(18525);
		when "0100100001011110" => data_out <= rom_array(18526);
		when "0100100001011111" => data_out <= rom_array(18527);
		when "0100100001100000" => data_out <= rom_array(18528);
		when "0100100001100001" => data_out <= rom_array(18529);
		when "0100100001100010" => data_out <= rom_array(18530);
		when "0100100001100011" => data_out <= rom_array(18531);
		when "0100100001100100" => data_out <= rom_array(18532);
		when "0100100001100101" => data_out <= rom_array(18533);
		when "0100100001100110" => data_out <= rom_array(18534);
		when "0100100001100111" => data_out <= rom_array(18535);
		when "0100100001101000" => data_out <= rom_array(18536);
		when "0100100001101001" => data_out <= rom_array(18537);
		when "0100100001101010" => data_out <= rom_array(18538);
		when "0100100001101011" => data_out <= rom_array(18539);
		when "0100100001101100" => data_out <= rom_array(18540);
		when "0100100001101101" => data_out <= rom_array(18541);
		when "0100100001101110" => data_out <= rom_array(18542);
		when "0100100001101111" => data_out <= rom_array(18543);
		when "0100100001110000" => data_out <= rom_array(18544);
		when "0100100001110001" => data_out <= rom_array(18545);
		when "0100100001110010" => data_out <= rom_array(18546);
		when "0100100001110011" => data_out <= rom_array(18547);
		when "0100100001110100" => data_out <= rom_array(18548);
		when "0100100001110101" => data_out <= rom_array(18549);
		when "0100100001110110" => data_out <= rom_array(18550);
		when "0100100001110111" => data_out <= rom_array(18551);
		when "0100100001111000" => data_out <= rom_array(18552);
		when "0100100001111001" => data_out <= rom_array(18553);
		when "0100100001111010" => data_out <= rom_array(18554);
		when "0100100001111011" => data_out <= rom_array(18555);
		when "0100100001111100" => data_out <= rom_array(18556);
		when "0100100001111101" => data_out <= rom_array(18557);
		when "0100100001111110" => data_out <= rom_array(18558);
		when "0100100001111111" => data_out <= rom_array(18559);
		when "0100100010000000" => data_out <= rom_array(18560);
		when "0100100010000001" => data_out <= rom_array(18561);
		when "0100100010000010" => data_out <= rom_array(18562);
		when "0100100010000011" => data_out <= rom_array(18563);
		when "0100100010000100" => data_out <= rom_array(18564);
		when "0100100010000101" => data_out <= rom_array(18565);
		when "0100100010000110" => data_out <= rom_array(18566);
		when "0100100010000111" => data_out <= rom_array(18567);
		when "0100100010001000" => data_out <= rom_array(18568);
		when "0100100010001001" => data_out <= rom_array(18569);
		when "0100100010001010" => data_out <= rom_array(18570);
		when "0100100010001011" => data_out <= rom_array(18571);
		when "0100100010001100" => data_out <= rom_array(18572);
		when "0100100010001101" => data_out <= rom_array(18573);
		when "0100100010001110" => data_out <= rom_array(18574);
		when "0100100010001111" => data_out <= rom_array(18575);
		when "0100100010010000" => data_out <= rom_array(18576);
		when "0100100010010001" => data_out <= rom_array(18577);
		when "0100100010010010" => data_out <= rom_array(18578);
		when "0100100010010011" => data_out <= rom_array(18579);
		when "0100100010010100" => data_out <= rom_array(18580);
		when "0100100010010101" => data_out <= rom_array(18581);
		when "0100100010010110" => data_out <= rom_array(18582);
		when "0100100010010111" => data_out <= rom_array(18583);
		when "0100100010011000" => data_out <= rom_array(18584);
		when "0100100010011001" => data_out <= rom_array(18585);
		when "0100100010011010" => data_out <= rom_array(18586);
		when "0100100010011011" => data_out <= rom_array(18587);
		when "0100100010011100" => data_out <= rom_array(18588);
		when "0100100010011101" => data_out <= rom_array(18589);
		when "0100100010011110" => data_out <= rom_array(18590);
		when "0100100010011111" => data_out <= rom_array(18591);
		when "0100100010100000" => data_out <= rom_array(18592);
		when "0100100010100001" => data_out <= rom_array(18593);
		when "0100100010100010" => data_out <= rom_array(18594);
		when "0100100010100011" => data_out <= rom_array(18595);
		when "0100100010100100" => data_out <= rom_array(18596);
		when "0100100010100101" => data_out <= rom_array(18597);
		when "0100100010100110" => data_out <= rom_array(18598);
		when "0100100010100111" => data_out <= rom_array(18599);
		when "0100100010101000" => data_out <= rom_array(18600);
		when "0100100010101001" => data_out <= rom_array(18601);
		when "0100100010101010" => data_out <= rom_array(18602);
		when "0100100010101011" => data_out <= rom_array(18603);
		when "0100100010101100" => data_out <= rom_array(18604);
		when "0100100010101101" => data_out <= rom_array(18605);
		when "0100100010101110" => data_out <= rom_array(18606);
		when "0100100010101111" => data_out <= rom_array(18607);
		when "0100100010110000" => data_out <= rom_array(18608);
		when "0100100010110001" => data_out <= rom_array(18609);
		when "0100100010110010" => data_out <= rom_array(18610);
		when "0100100010110011" => data_out <= rom_array(18611);
		when "0100100010110100" => data_out <= rom_array(18612);
		when "0100100010110101" => data_out <= rom_array(18613);
		when "0100100010110110" => data_out <= rom_array(18614);
		when "0100100010110111" => data_out <= rom_array(18615);
		when "0100100010111000" => data_out <= rom_array(18616);
		when "0100100010111001" => data_out <= rom_array(18617);
		when "0100100010111010" => data_out <= rom_array(18618);
		when "0100100010111011" => data_out <= rom_array(18619);
		when "0100100010111100" => data_out <= rom_array(18620);
		when "0100100010111101" => data_out <= rom_array(18621);
		when "0100100010111110" => data_out <= rom_array(18622);
		when "0100100010111111" => data_out <= rom_array(18623);
		when "0100100011000000" => data_out <= rom_array(18624);
		when "0100100011000001" => data_out <= rom_array(18625);
		when "0100100011000010" => data_out <= rom_array(18626);
		when "0100100011000011" => data_out <= rom_array(18627);
		when "0100100011000100" => data_out <= rom_array(18628);
		when "0100100011000101" => data_out <= rom_array(18629);
		when "0100100011000110" => data_out <= rom_array(18630);
		when "0100100011000111" => data_out <= rom_array(18631);
		when "0100100011001000" => data_out <= rom_array(18632);
		when "0100100011001001" => data_out <= rom_array(18633);
		when "0100100011001010" => data_out <= rom_array(18634);
		when "0100100011001011" => data_out <= rom_array(18635);
		when "0100100011001100" => data_out <= rom_array(18636);
		when "0100100011001101" => data_out <= rom_array(18637);
		when "0100100011001110" => data_out <= rom_array(18638);
		when "0100100011001111" => data_out <= rom_array(18639);
		when "0100100011010000" => data_out <= rom_array(18640);
		when "0100100011010001" => data_out <= rom_array(18641);
		when "0100100011010010" => data_out <= rom_array(18642);
		when "0100100011010011" => data_out <= rom_array(18643);
		when "0100100011010100" => data_out <= rom_array(18644);
		when "0100100011010101" => data_out <= rom_array(18645);
		when "0100100011010110" => data_out <= rom_array(18646);
		when "0100100011010111" => data_out <= rom_array(18647);
		when "0100100011011000" => data_out <= rom_array(18648);
		when "0100100011011001" => data_out <= rom_array(18649);
		when "0100100011011010" => data_out <= rom_array(18650);
		when "0100100011011011" => data_out <= rom_array(18651);
		when "0100100011011100" => data_out <= rom_array(18652);
		when "0100100011011101" => data_out <= rom_array(18653);
		when "0100100011011110" => data_out <= rom_array(18654);
		when "0100100011011111" => data_out <= rom_array(18655);
		when "0100100011100000" => data_out <= rom_array(18656);
		when "0100100011100001" => data_out <= rom_array(18657);
		when "0100100011100010" => data_out <= rom_array(18658);
		when "0100100011100011" => data_out <= rom_array(18659);
		when "0100100011100100" => data_out <= rom_array(18660);
		when "0100100011100101" => data_out <= rom_array(18661);
		when "0100100011100110" => data_out <= rom_array(18662);
		when "0100100011100111" => data_out <= rom_array(18663);
		when "0100100011101000" => data_out <= rom_array(18664);
		when "0100100011101001" => data_out <= rom_array(18665);
		when "0100100011101010" => data_out <= rom_array(18666);
		when "0100100011101011" => data_out <= rom_array(18667);
		when "0100100011101100" => data_out <= rom_array(18668);
		when "0100100011101101" => data_out <= rom_array(18669);
		when "0100100011101110" => data_out <= rom_array(18670);
		when "0100100011101111" => data_out <= rom_array(18671);
		when "0100100011110000" => data_out <= rom_array(18672);
		when "0100100011110001" => data_out <= rom_array(18673);
		when "0100100011110010" => data_out <= rom_array(18674);
		when "0100100011110011" => data_out <= rom_array(18675);
		when "0100100011110100" => data_out <= rom_array(18676);
		when "0100100011110101" => data_out <= rom_array(18677);
		when "0100100011110110" => data_out <= rom_array(18678);
		when "0100100011110111" => data_out <= rom_array(18679);
		when "0100100011111000" => data_out <= rom_array(18680);
		when "0100100011111001" => data_out <= rom_array(18681);
		when "0100100011111010" => data_out <= rom_array(18682);
		when "0100100011111011" => data_out <= rom_array(18683);
		when "0100100011111100" => data_out <= rom_array(18684);
		when "0100100011111101" => data_out <= rom_array(18685);
		when "0100100011111110" => data_out <= rom_array(18686);
		when "0100100011111111" => data_out <= rom_array(18687);
		when "0100100100000000" => data_out <= rom_array(18688);
		when "0100100100000001" => data_out <= rom_array(18689);
		when "0100100100000010" => data_out <= rom_array(18690);
		when "0100100100000011" => data_out <= rom_array(18691);
		when "0100100100000100" => data_out <= rom_array(18692);
		when "0100100100000101" => data_out <= rom_array(18693);
		when "0100100100000110" => data_out <= rom_array(18694);
		when "0100100100000111" => data_out <= rom_array(18695);
		when "0100100100001000" => data_out <= rom_array(18696);
		when "0100100100001001" => data_out <= rom_array(18697);
		when "0100100100001010" => data_out <= rom_array(18698);
		when "0100100100001011" => data_out <= rom_array(18699);
		when "0100100100001100" => data_out <= rom_array(18700);
		when "0100100100001101" => data_out <= rom_array(18701);
		when "0100100100001110" => data_out <= rom_array(18702);
		when "0100100100001111" => data_out <= rom_array(18703);
		when "0100100100010000" => data_out <= rom_array(18704);
		when "0100100100010001" => data_out <= rom_array(18705);
		when "0100100100010010" => data_out <= rom_array(18706);
		when "0100100100010011" => data_out <= rom_array(18707);
		when "0100100100010100" => data_out <= rom_array(18708);
		when "0100100100010101" => data_out <= rom_array(18709);
		when "0100100100010110" => data_out <= rom_array(18710);
		when "0100100100010111" => data_out <= rom_array(18711);
		when "0100100100011000" => data_out <= rom_array(18712);
		when "0100100100011001" => data_out <= rom_array(18713);
		when "0100100100011010" => data_out <= rom_array(18714);
		when "0100100100011011" => data_out <= rom_array(18715);
		when "0100100100011100" => data_out <= rom_array(18716);
		when "0100100100011101" => data_out <= rom_array(18717);
		when "0100100100011110" => data_out <= rom_array(18718);
		when "0100100100011111" => data_out <= rom_array(18719);
		when "0100100100100000" => data_out <= rom_array(18720);
		when "0100100100100001" => data_out <= rom_array(18721);
		when "0100100100100010" => data_out <= rom_array(18722);
		when "0100100100100011" => data_out <= rom_array(18723);
		when "0100100100100100" => data_out <= rom_array(18724);
		when "0100100100100101" => data_out <= rom_array(18725);
		when "0100100100100110" => data_out <= rom_array(18726);
		when "0100100100100111" => data_out <= rom_array(18727);
		when "0100100100101000" => data_out <= rom_array(18728);
		when "0100100100101001" => data_out <= rom_array(18729);
		when "0100100100101010" => data_out <= rom_array(18730);
		when "0100100100101011" => data_out <= rom_array(18731);
		when "0100100100101100" => data_out <= rom_array(18732);
		when "0100100100101101" => data_out <= rom_array(18733);
		when "0100100100101110" => data_out <= rom_array(18734);
		when "0100100100101111" => data_out <= rom_array(18735);
		when "0100100100110000" => data_out <= rom_array(18736);
		when "0100100100110001" => data_out <= rom_array(18737);
		when "0100100100110010" => data_out <= rom_array(18738);
		when "0100100100110011" => data_out <= rom_array(18739);
		when "0100100100110100" => data_out <= rom_array(18740);
		when "0100100100110101" => data_out <= rom_array(18741);
		when "0100100100110110" => data_out <= rom_array(18742);
		when "0100100100110111" => data_out <= rom_array(18743);
		when "0100100100111000" => data_out <= rom_array(18744);
		when "0100100100111001" => data_out <= rom_array(18745);
		when "0100100100111010" => data_out <= rom_array(18746);
		when "0100100100111011" => data_out <= rom_array(18747);
		when "0100100100111100" => data_out <= rom_array(18748);
		when "0100100100111101" => data_out <= rom_array(18749);
		when "0100100100111110" => data_out <= rom_array(18750);
		when "0100100100111111" => data_out <= rom_array(18751);
		when "0100100101000000" => data_out <= rom_array(18752);
		when "0100100101000001" => data_out <= rom_array(18753);
		when "0100100101000010" => data_out <= rom_array(18754);
		when "0100100101000011" => data_out <= rom_array(18755);
		when "0100100101000100" => data_out <= rom_array(18756);
		when "0100100101000101" => data_out <= rom_array(18757);
		when "0100100101000110" => data_out <= rom_array(18758);
		when "0100100101000111" => data_out <= rom_array(18759);
		when "0100100101001000" => data_out <= rom_array(18760);
		when "0100100101001001" => data_out <= rom_array(18761);
		when "0100100101001010" => data_out <= rom_array(18762);
		when "0100100101001011" => data_out <= rom_array(18763);
		when "0100100101001100" => data_out <= rom_array(18764);
		when "0100100101001101" => data_out <= rom_array(18765);
		when "0100100101001110" => data_out <= rom_array(18766);
		when "0100100101001111" => data_out <= rom_array(18767);
		when "0100100101010000" => data_out <= rom_array(18768);
		when "0100100101010001" => data_out <= rom_array(18769);
		when "0100100101010010" => data_out <= rom_array(18770);
		when "0100100101010011" => data_out <= rom_array(18771);
		when "0100100101010100" => data_out <= rom_array(18772);
		when "0100100101010101" => data_out <= rom_array(18773);
		when "0100100101010110" => data_out <= rom_array(18774);
		when "0100100101010111" => data_out <= rom_array(18775);
		when "0100100101011000" => data_out <= rom_array(18776);
		when "0100100101011001" => data_out <= rom_array(18777);
		when "0100100101011010" => data_out <= rom_array(18778);
		when "0100100101011011" => data_out <= rom_array(18779);
		when "0100100101011100" => data_out <= rom_array(18780);
		when "0100100101011101" => data_out <= rom_array(18781);
		when "0100100101011110" => data_out <= rom_array(18782);
		when "0100100101011111" => data_out <= rom_array(18783);
		when "0100100101100000" => data_out <= rom_array(18784);
		when "0100100101100001" => data_out <= rom_array(18785);
		when "0100100101100010" => data_out <= rom_array(18786);
		when "0100100101100011" => data_out <= rom_array(18787);
		when "0100100101100100" => data_out <= rom_array(18788);
		when "0100100101100101" => data_out <= rom_array(18789);
		when "0100100101100110" => data_out <= rom_array(18790);
		when "0100100101100111" => data_out <= rom_array(18791);
		when "0100100101101000" => data_out <= rom_array(18792);
		when "0100100101101001" => data_out <= rom_array(18793);
		when "0100100101101010" => data_out <= rom_array(18794);
		when "0100100101101011" => data_out <= rom_array(18795);
		when "0100100101101100" => data_out <= rom_array(18796);
		when "0100100101101101" => data_out <= rom_array(18797);
		when "0100100101101110" => data_out <= rom_array(18798);
		when "0100100101101111" => data_out <= rom_array(18799);
		when "0100100101110000" => data_out <= rom_array(18800);
		when "0100100101110001" => data_out <= rom_array(18801);
		when "0100100101110010" => data_out <= rom_array(18802);
		when "0100100101110011" => data_out <= rom_array(18803);
		when "0100100101110100" => data_out <= rom_array(18804);
		when "0100100101110101" => data_out <= rom_array(18805);
		when "0100100101110110" => data_out <= rom_array(18806);
		when "0100100101110111" => data_out <= rom_array(18807);
		when "0100100101111000" => data_out <= rom_array(18808);
		when "0100100101111001" => data_out <= rom_array(18809);
		when "0100100101111010" => data_out <= rom_array(18810);
		when "0100100101111011" => data_out <= rom_array(18811);
		when "0100100101111100" => data_out <= rom_array(18812);
		when "0100100101111101" => data_out <= rom_array(18813);
		when "0100100101111110" => data_out <= rom_array(18814);
		when "0100100101111111" => data_out <= rom_array(18815);
		when "0100100110000000" => data_out <= rom_array(18816);
		when "0100100110000001" => data_out <= rom_array(18817);
		when "0100100110000010" => data_out <= rom_array(18818);
		when "0100100110000011" => data_out <= rom_array(18819);
		when "0100100110000100" => data_out <= rom_array(18820);
		when "0100100110000101" => data_out <= rom_array(18821);
		when "0100100110000110" => data_out <= rom_array(18822);
		when "0100100110000111" => data_out <= rom_array(18823);
		when "0100100110001000" => data_out <= rom_array(18824);
		when "0100100110001001" => data_out <= rom_array(18825);
		when "0100100110001010" => data_out <= rom_array(18826);
		when "0100100110001011" => data_out <= rom_array(18827);
		when "0100100110001100" => data_out <= rom_array(18828);
		when "0100100110001101" => data_out <= rom_array(18829);
		when "0100100110001110" => data_out <= rom_array(18830);
		when "0100100110001111" => data_out <= rom_array(18831);
		when "0100100110010000" => data_out <= rom_array(18832);
		when "0100100110010001" => data_out <= rom_array(18833);
		when "0100100110010010" => data_out <= rom_array(18834);
		when "0100100110010011" => data_out <= rom_array(18835);
		when "0100100110010100" => data_out <= rom_array(18836);
		when "0100100110010101" => data_out <= rom_array(18837);
		when "0100100110010110" => data_out <= rom_array(18838);
		when "0100100110010111" => data_out <= rom_array(18839);
		when "0100100110011000" => data_out <= rom_array(18840);
		when "0100100110011001" => data_out <= rom_array(18841);
		when "0100100110011010" => data_out <= rom_array(18842);
		when "0100100110011011" => data_out <= rom_array(18843);
		when "0100100110011100" => data_out <= rom_array(18844);
		when "0100100110011101" => data_out <= rom_array(18845);
		when "0100100110011110" => data_out <= rom_array(18846);
		when "0100100110011111" => data_out <= rom_array(18847);
		when "0100100110100000" => data_out <= rom_array(18848);
		when "0100100110100001" => data_out <= rom_array(18849);
		when "0100100110100010" => data_out <= rom_array(18850);
		when "0100100110100011" => data_out <= rom_array(18851);
		when "0100100110100100" => data_out <= rom_array(18852);
		when "0100100110100101" => data_out <= rom_array(18853);
		when "0100100110100110" => data_out <= rom_array(18854);
		when "0100100110100111" => data_out <= rom_array(18855);
		when "0100100110101000" => data_out <= rom_array(18856);
		when "0100100110101001" => data_out <= rom_array(18857);
		when "0100100110101010" => data_out <= rom_array(18858);
		when "0100100110101011" => data_out <= rom_array(18859);
		when "0100100110101100" => data_out <= rom_array(18860);
		when "0100100110101101" => data_out <= rom_array(18861);
		when "0100100110101110" => data_out <= rom_array(18862);
		when "0100100110101111" => data_out <= rom_array(18863);
		when "0100100110110000" => data_out <= rom_array(18864);
		when "0100100110110001" => data_out <= rom_array(18865);
		when "0100100110110010" => data_out <= rom_array(18866);
		when "0100100110110011" => data_out <= rom_array(18867);
		when "0100100110110100" => data_out <= rom_array(18868);
		when "0100100110110101" => data_out <= rom_array(18869);
		when "0100100110110110" => data_out <= rom_array(18870);
		when "0100100110110111" => data_out <= rom_array(18871);
		when "0100100110111000" => data_out <= rom_array(18872);
		when "0100100110111001" => data_out <= rom_array(18873);
		when "0100100110111010" => data_out <= rom_array(18874);
		when "0100100110111011" => data_out <= rom_array(18875);
		when "0100100110111100" => data_out <= rom_array(18876);
		when "0100100110111101" => data_out <= rom_array(18877);
		when "0100100110111110" => data_out <= rom_array(18878);
		when "0100100110111111" => data_out <= rom_array(18879);
		when "0100100111000000" => data_out <= rom_array(18880);
		when "0100100111000001" => data_out <= rom_array(18881);
		when "0100100111000010" => data_out <= rom_array(18882);
		when "0100100111000011" => data_out <= rom_array(18883);
		when "0100100111000100" => data_out <= rom_array(18884);
		when "0100100111000101" => data_out <= rom_array(18885);
		when "0100100111000110" => data_out <= rom_array(18886);
		when "0100100111000111" => data_out <= rom_array(18887);
		when "0100100111001000" => data_out <= rom_array(18888);
		when "0100100111001001" => data_out <= rom_array(18889);
		when "0100100111001010" => data_out <= rom_array(18890);
		when "0100100111001011" => data_out <= rom_array(18891);
		when "0100100111001100" => data_out <= rom_array(18892);
		when "0100100111001101" => data_out <= rom_array(18893);
		when "0100100111001110" => data_out <= rom_array(18894);
		when "0100100111001111" => data_out <= rom_array(18895);
		when "0100100111010000" => data_out <= rom_array(18896);
		when "0100100111010001" => data_out <= rom_array(18897);
		when "0100100111010010" => data_out <= rom_array(18898);
		when "0100100111010011" => data_out <= rom_array(18899);
		when "0100100111010100" => data_out <= rom_array(18900);
		when "0100100111010101" => data_out <= rom_array(18901);
		when "0100100111010110" => data_out <= rom_array(18902);
		when "0100100111010111" => data_out <= rom_array(18903);
		when "0100100111011000" => data_out <= rom_array(18904);
		when "0100100111011001" => data_out <= rom_array(18905);
		when "0100100111011010" => data_out <= rom_array(18906);
		when "0100100111011011" => data_out <= rom_array(18907);
		when "0100100111011100" => data_out <= rom_array(18908);
		when "0100100111011101" => data_out <= rom_array(18909);
		when "0100100111011110" => data_out <= rom_array(18910);
		when "0100100111011111" => data_out <= rom_array(18911);
		when "0100100111100000" => data_out <= rom_array(18912);
		when "0100100111100001" => data_out <= rom_array(18913);
		when "0100100111100010" => data_out <= rom_array(18914);
		when "0100100111100011" => data_out <= rom_array(18915);
		when "0100100111100100" => data_out <= rom_array(18916);
		when "0100100111100101" => data_out <= rom_array(18917);
		when "0100100111100110" => data_out <= rom_array(18918);
		when "0100100111100111" => data_out <= rom_array(18919);
		when "0100100111101000" => data_out <= rom_array(18920);
		when "0100100111101001" => data_out <= rom_array(18921);
		when "0100100111101010" => data_out <= rom_array(18922);
		when "0100100111101011" => data_out <= rom_array(18923);
		when "0100100111101100" => data_out <= rom_array(18924);
		when "0100100111101101" => data_out <= rom_array(18925);
		when "0100100111101110" => data_out <= rom_array(18926);
		when "0100100111101111" => data_out <= rom_array(18927);
		when "0100100111110000" => data_out <= rom_array(18928);
		when "0100100111110001" => data_out <= rom_array(18929);
		when "0100100111110010" => data_out <= rom_array(18930);
		when "0100100111110011" => data_out <= rom_array(18931);
		when "0100100111110100" => data_out <= rom_array(18932);
		when "0100100111110101" => data_out <= rom_array(18933);
		when "0100100111110110" => data_out <= rom_array(18934);
		when "0100100111110111" => data_out <= rom_array(18935);
		when "0100100111111000" => data_out <= rom_array(18936);
		when "0100100111111001" => data_out <= rom_array(18937);
		when "0100100111111010" => data_out <= rom_array(18938);
		when "0100100111111011" => data_out <= rom_array(18939);
		when "0100100111111100" => data_out <= rom_array(18940);
		when "0100100111111101" => data_out <= rom_array(18941);
		when "0100100111111110" => data_out <= rom_array(18942);
		when "0100100111111111" => data_out <= rom_array(18943);
		when "0100101000000000" => data_out <= rom_array(18944);
		when "0100101000000001" => data_out <= rom_array(18945);
		when "0100101000000010" => data_out <= rom_array(18946);
		when "0100101000000011" => data_out <= rom_array(18947);
		when "0100101000000100" => data_out <= rom_array(18948);
		when "0100101000000101" => data_out <= rom_array(18949);
		when "0100101000000110" => data_out <= rom_array(18950);
		when "0100101000000111" => data_out <= rom_array(18951);
		when "0100101000001000" => data_out <= rom_array(18952);
		when "0100101000001001" => data_out <= rom_array(18953);
		when "0100101000001010" => data_out <= rom_array(18954);
		when "0100101000001011" => data_out <= rom_array(18955);
		when "0100101000001100" => data_out <= rom_array(18956);
		when "0100101000001101" => data_out <= rom_array(18957);
		when "0100101000001110" => data_out <= rom_array(18958);
		when "0100101000001111" => data_out <= rom_array(18959);
		when "0100101000010000" => data_out <= rom_array(18960);
		when "0100101000010001" => data_out <= rom_array(18961);
		when "0100101000010010" => data_out <= rom_array(18962);
		when "0100101000010011" => data_out <= rom_array(18963);
		when "0100101000010100" => data_out <= rom_array(18964);
		when "0100101000010101" => data_out <= rom_array(18965);
		when "0100101000010110" => data_out <= rom_array(18966);
		when "0100101000010111" => data_out <= rom_array(18967);
		when "0100101000011000" => data_out <= rom_array(18968);
		when "0100101000011001" => data_out <= rom_array(18969);
		when "0100101000011010" => data_out <= rom_array(18970);
		when "0100101000011011" => data_out <= rom_array(18971);
		when "0100101000011100" => data_out <= rom_array(18972);
		when "0100101000011101" => data_out <= rom_array(18973);
		when "0100101000011110" => data_out <= rom_array(18974);
		when "0100101000011111" => data_out <= rom_array(18975);
		when "0100101000100000" => data_out <= rom_array(18976);
		when "0100101000100001" => data_out <= rom_array(18977);
		when "0100101000100010" => data_out <= rom_array(18978);
		when "0100101000100011" => data_out <= rom_array(18979);
		when "0100101000100100" => data_out <= rom_array(18980);
		when "0100101000100101" => data_out <= rom_array(18981);
		when "0100101000100110" => data_out <= rom_array(18982);
		when "0100101000100111" => data_out <= rom_array(18983);
		when "0100101000101000" => data_out <= rom_array(18984);
		when "0100101000101001" => data_out <= rom_array(18985);
		when "0100101000101010" => data_out <= rom_array(18986);
		when "0100101000101011" => data_out <= rom_array(18987);
		when "0100101000101100" => data_out <= rom_array(18988);
		when "0100101000101101" => data_out <= rom_array(18989);
		when "0100101000101110" => data_out <= rom_array(18990);
		when "0100101000101111" => data_out <= rom_array(18991);
		when "0100101000110000" => data_out <= rom_array(18992);
		when "0100101000110001" => data_out <= rom_array(18993);
		when "0100101000110010" => data_out <= rom_array(18994);
		when "0100101000110011" => data_out <= rom_array(18995);
		when "0100101000110100" => data_out <= rom_array(18996);
		when "0100101000110101" => data_out <= rom_array(18997);
		when "0100101000110110" => data_out <= rom_array(18998);
		when "0100101000110111" => data_out <= rom_array(18999);
		when "0100101000111000" => data_out <= rom_array(19000);
		when "0100101000111001" => data_out <= rom_array(19001);
		when "0100101000111010" => data_out <= rom_array(19002);
		when "0100101000111011" => data_out <= rom_array(19003);
		when "0100101000111100" => data_out <= rom_array(19004);
		when "0100101000111101" => data_out <= rom_array(19005);
		when "0100101000111110" => data_out <= rom_array(19006);
		when "0100101000111111" => data_out <= rom_array(19007);
		when "0100101001000000" => data_out <= rom_array(19008);
		when "0100101001000001" => data_out <= rom_array(19009);
		when "0100101001000010" => data_out <= rom_array(19010);
		when "0100101001000011" => data_out <= rom_array(19011);
		when "0100101001000100" => data_out <= rom_array(19012);
		when "0100101001000101" => data_out <= rom_array(19013);
		when "0100101001000110" => data_out <= rom_array(19014);
		when "0100101001000111" => data_out <= rom_array(19015);
		when "0100101001001000" => data_out <= rom_array(19016);
		when "0100101001001001" => data_out <= rom_array(19017);
		when "0100101001001010" => data_out <= rom_array(19018);
		when "0100101001001011" => data_out <= rom_array(19019);
		when "0100101001001100" => data_out <= rom_array(19020);
		when "0100101001001101" => data_out <= rom_array(19021);
		when "0100101001001110" => data_out <= rom_array(19022);
		when "0100101001001111" => data_out <= rom_array(19023);
		when "0100101001010000" => data_out <= rom_array(19024);
		when "0100101001010001" => data_out <= rom_array(19025);
		when "0100101001010010" => data_out <= rom_array(19026);
		when "0100101001010011" => data_out <= rom_array(19027);
		when "0100101001010100" => data_out <= rom_array(19028);
		when "0100101001010101" => data_out <= rom_array(19029);
		when "0100101001010110" => data_out <= rom_array(19030);
		when "0100101001010111" => data_out <= rom_array(19031);
		when "0100101001011000" => data_out <= rom_array(19032);
		when "0100101001011001" => data_out <= rom_array(19033);
		when "0100101001011010" => data_out <= rom_array(19034);
		when "0100101001011011" => data_out <= rom_array(19035);
		when "0100101001011100" => data_out <= rom_array(19036);
		when "0100101001011101" => data_out <= rom_array(19037);
		when "0100101001011110" => data_out <= rom_array(19038);
		when "0100101001011111" => data_out <= rom_array(19039);
		when "0100101001100000" => data_out <= rom_array(19040);
		when "0100101001100001" => data_out <= rom_array(19041);
		when "0100101001100010" => data_out <= rom_array(19042);
		when "0100101001100011" => data_out <= rom_array(19043);
		when "0100101001100100" => data_out <= rom_array(19044);
		when "0100101001100101" => data_out <= rom_array(19045);
		when "0100101001100110" => data_out <= rom_array(19046);
		when "0100101001100111" => data_out <= rom_array(19047);
		when "0100101001101000" => data_out <= rom_array(19048);
		when "0100101001101001" => data_out <= rom_array(19049);
		when "0100101001101010" => data_out <= rom_array(19050);
		when "0100101001101011" => data_out <= rom_array(19051);
		when "0100101001101100" => data_out <= rom_array(19052);
		when "0100101001101101" => data_out <= rom_array(19053);
		when "0100101001101110" => data_out <= rom_array(19054);
		when "0100101001101111" => data_out <= rom_array(19055);
		when "0100101001110000" => data_out <= rom_array(19056);
		when "0100101001110001" => data_out <= rom_array(19057);
		when "0100101001110010" => data_out <= rom_array(19058);
		when "0100101001110011" => data_out <= rom_array(19059);
		when "0100101001110100" => data_out <= rom_array(19060);
		when "0100101001110101" => data_out <= rom_array(19061);
		when "0100101001110110" => data_out <= rom_array(19062);
		when "0100101001110111" => data_out <= rom_array(19063);
		when "0100101001111000" => data_out <= rom_array(19064);
		when "0100101001111001" => data_out <= rom_array(19065);
		when "0100101001111010" => data_out <= rom_array(19066);
		when "0100101001111011" => data_out <= rom_array(19067);
		when "0100101001111100" => data_out <= rom_array(19068);
		when "0100101001111101" => data_out <= rom_array(19069);
		when "0100101001111110" => data_out <= rom_array(19070);
		when "0100101001111111" => data_out <= rom_array(19071);
		when "0100101010000000" => data_out <= rom_array(19072);
		when "0100101010000001" => data_out <= rom_array(19073);
		when "0100101010000010" => data_out <= rom_array(19074);
		when "0100101010000011" => data_out <= rom_array(19075);
		when "0100101010000100" => data_out <= rom_array(19076);
		when "0100101010000101" => data_out <= rom_array(19077);
		when "0100101010000110" => data_out <= rom_array(19078);
		when "0100101010000111" => data_out <= rom_array(19079);
		when "0100101010001000" => data_out <= rom_array(19080);
		when "0100101010001001" => data_out <= rom_array(19081);
		when "0100101010001010" => data_out <= rom_array(19082);
		when "0100101010001011" => data_out <= rom_array(19083);
		when "0100101010001100" => data_out <= rom_array(19084);
		when "0100101010001101" => data_out <= rom_array(19085);
		when "0100101010001110" => data_out <= rom_array(19086);
		when "0100101010001111" => data_out <= rom_array(19087);
		when "0100101010010000" => data_out <= rom_array(19088);
		when "0100101010010001" => data_out <= rom_array(19089);
		when "0100101010010010" => data_out <= rom_array(19090);
		when "0100101010010011" => data_out <= rom_array(19091);
		when "0100101010010100" => data_out <= rom_array(19092);
		when "0100101010010101" => data_out <= rom_array(19093);
		when "0100101010010110" => data_out <= rom_array(19094);
		when "0100101010010111" => data_out <= rom_array(19095);
		when "0100101010011000" => data_out <= rom_array(19096);
		when "0100101010011001" => data_out <= rom_array(19097);
		when "0100101010011010" => data_out <= rom_array(19098);
		when "0100101010011011" => data_out <= rom_array(19099);
		when "0100101010011100" => data_out <= rom_array(19100);
		when "0100101010011101" => data_out <= rom_array(19101);
		when "0100101010011110" => data_out <= rom_array(19102);
		when "0100101010011111" => data_out <= rom_array(19103);
		when "0100101010100000" => data_out <= rom_array(19104);
		when "0100101010100001" => data_out <= rom_array(19105);
		when "0100101010100010" => data_out <= rom_array(19106);
		when "0100101010100011" => data_out <= rom_array(19107);
		when "0100101010100100" => data_out <= rom_array(19108);
		when "0100101010100101" => data_out <= rom_array(19109);
		when "0100101010100110" => data_out <= rom_array(19110);
		when "0100101010100111" => data_out <= rom_array(19111);
		when "0100101010101000" => data_out <= rom_array(19112);
		when "0100101010101001" => data_out <= rom_array(19113);
		when "0100101010101010" => data_out <= rom_array(19114);
		when "0100101010101011" => data_out <= rom_array(19115);
		when "0100101010101100" => data_out <= rom_array(19116);
		when "0100101010101101" => data_out <= rom_array(19117);
		when "0100101010101110" => data_out <= rom_array(19118);
		when "0100101010101111" => data_out <= rom_array(19119);
		when "0100101010110000" => data_out <= rom_array(19120);
		when "0100101010110001" => data_out <= rom_array(19121);
		when "0100101010110010" => data_out <= rom_array(19122);
		when "0100101010110011" => data_out <= rom_array(19123);
		when "0100101010110100" => data_out <= rom_array(19124);
		when "0100101010110101" => data_out <= rom_array(19125);
		when "0100101010110110" => data_out <= rom_array(19126);
		when "0100101010110111" => data_out <= rom_array(19127);
		when "0100101010111000" => data_out <= rom_array(19128);
		when "0100101010111001" => data_out <= rom_array(19129);
		when "0100101010111010" => data_out <= rom_array(19130);
		when "0100101010111011" => data_out <= rom_array(19131);
		when "0100101010111100" => data_out <= rom_array(19132);
		when "0100101010111101" => data_out <= rom_array(19133);
		when "0100101010111110" => data_out <= rom_array(19134);
		when "0100101010111111" => data_out <= rom_array(19135);
		when "0100101011000000" => data_out <= rom_array(19136);
		when "0100101011000001" => data_out <= rom_array(19137);
		when "0100101011000010" => data_out <= rom_array(19138);
		when "0100101011000011" => data_out <= rom_array(19139);
		when "0100101011000100" => data_out <= rom_array(19140);
		when "0100101011000101" => data_out <= rom_array(19141);
		when "0100101011000110" => data_out <= rom_array(19142);
		when "0100101011000111" => data_out <= rom_array(19143);
		when "0100101011001000" => data_out <= rom_array(19144);
		when "0100101011001001" => data_out <= rom_array(19145);
		when "0100101011001010" => data_out <= rom_array(19146);
		when "0100101011001011" => data_out <= rom_array(19147);
		when "0100101011001100" => data_out <= rom_array(19148);
		when "0100101011001101" => data_out <= rom_array(19149);
		when "0100101011001110" => data_out <= rom_array(19150);
		when "0100101011001111" => data_out <= rom_array(19151);
		when "0100101011010000" => data_out <= rom_array(19152);
		when "0100101011010001" => data_out <= rom_array(19153);
		when "0100101011010010" => data_out <= rom_array(19154);
		when "0100101011010011" => data_out <= rom_array(19155);
		when "0100101011010100" => data_out <= rom_array(19156);
		when "0100101011010101" => data_out <= rom_array(19157);
		when "0100101011010110" => data_out <= rom_array(19158);
		when "0100101011010111" => data_out <= rom_array(19159);
		when "0100101011011000" => data_out <= rom_array(19160);
		when "0100101011011001" => data_out <= rom_array(19161);
		when "0100101011011010" => data_out <= rom_array(19162);
		when "0100101011011011" => data_out <= rom_array(19163);
		when "0100101011011100" => data_out <= rom_array(19164);
		when "0100101011011101" => data_out <= rom_array(19165);
		when "0100101011011110" => data_out <= rom_array(19166);
		when "0100101011011111" => data_out <= rom_array(19167);
		when "0100101011100000" => data_out <= rom_array(19168);
		when "0100101011100001" => data_out <= rom_array(19169);
		when "0100101011100010" => data_out <= rom_array(19170);
		when "0100101011100011" => data_out <= rom_array(19171);
		when "0100101011100100" => data_out <= rom_array(19172);
		when "0100101011100101" => data_out <= rom_array(19173);
		when "0100101011100110" => data_out <= rom_array(19174);
		when "0100101011100111" => data_out <= rom_array(19175);
		when "0100101011101000" => data_out <= rom_array(19176);
		when "0100101011101001" => data_out <= rom_array(19177);
		when "0100101011101010" => data_out <= rom_array(19178);
		when "0100101011101011" => data_out <= rom_array(19179);
		when "0100101011101100" => data_out <= rom_array(19180);
		when "0100101011101101" => data_out <= rom_array(19181);
		when "0100101011101110" => data_out <= rom_array(19182);
		when "0100101011101111" => data_out <= rom_array(19183);
		when "0100101011110000" => data_out <= rom_array(19184);
		when "0100101011110001" => data_out <= rom_array(19185);
		when "0100101011110010" => data_out <= rom_array(19186);
		when "0100101011110011" => data_out <= rom_array(19187);
		when "0100101011110100" => data_out <= rom_array(19188);
		when "0100101011110101" => data_out <= rom_array(19189);
		when "0100101011110110" => data_out <= rom_array(19190);
		when "0100101011110111" => data_out <= rom_array(19191);
		when "0100101011111000" => data_out <= rom_array(19192);
		when "0100101011111001" => data_out <= rom_array(19193);
		when "0100101011111010" => data_out <= rom_array(19194);
		when "0100101011111011" => data_out <= rom_array(19195);
		when "0100101011111100" => data_out <= rom_array(19196);
		when "0100101011111101" => data_out <= rom_array(19197);
		when "0100101011111110" => data_out <= rom_array(19198);
		when "0100101011111111" => data_out <= rom_array(19199);
		when "0100101100000000" => data_out <= rom_array(19200);
		when "0100101100000001" => data_out <= rom_array(19201);
		when "0100101100000010" => data_out <= rom_array(19202);
		when "0100101100000011" => data_out <= rom_array(19203);
		when "0100101100000100" => data_out <= rom_array(19204);
		when "0100101100000101" => data_out <= rom_array(19205);
		when "0100101100000110" => data_out <= rom_array(19206);
		when "0100101100000111" => data_out <= rom_array(19207);
		when "0100101100001000" => data_out <= rom_array(19208);
		when "0100101100001001" => data_out <= rom_array(19209);
		when "0100101100001010" => data_out <= rom_array(19210);
		when "0100101100001011" => data_out <= rom_array(19211);
		when "0100101100001100" => data_out <= rom_array(19212);
		when "0100101100001101" => data_out <= rom_array(19213);
		when "0100101100001110" => data_out <= rom_array(19214);
		when "0100101100001111" => data_out <= rom_array(19215);
		when "0100101100010000" => data_out <= rom_array(19216);
		when "0100101100010001" => data_out <= rom_array(19217);
		when "0100101100010010" => data_out <= rom_array(19218);
		when "0100101100010011" => data_out <= rom_array(19219);
		when "0100101100010100" => data_out <= rom_array(19220);
		when "0100101100010101" => data_out <= rom_array(19221);
		when "0100101100010110" => data_out <= rom_array(19222);
		when "0100101100010111" => data_out <= rom_array(19223);
		when "0100101100011000" => data_out <= rom_array(19224);
		when "0100101100011001" => data_out <= rom_array(19225);
		when "0100101100011010" => data_out <= rom_array(19226);
		when "0100101100011011" => data_out <= rom_array(19227);
		when "0100101100011100" => data_out <= rom_array(19228);
		when "0100101100011101" => data_out <= rom_array(19229);
		when "0100101100011110" => data_out <= rom_array(19230);
		when "0100101100011111" => data_out <= rom_array(19231);
		when "0100101100100000" => data_out <= rom_array(19232);
		when "0100101100100001" => data_out <= rom_array(19233);
		when "0100101100100010" => data_out <= rom_array(19234);
		when "0100101100100011" => data_out <= rom_array(19235);
		when "0100101100100100" => data_out <= rom_array(19236);
		when "0100101100100101" => data_out <= rom_array(19237);
		when "0100101100100110" => data_out <= rom_array(19238);
		when "0100101100100111" => data_out <= rom_array(19239);
		when "0100101100101000" => data_out <= rom_array(19240);
		when "0100101100101001" => data_out <= rom_array(19241);
		when "0100101100101010" => data_out <= rom_array(19242);
		when "0100101100101011" => data_out <= rom_array(19243);
		when "0100101100101100" => data_out <= rom_array(19244);
		when "0100101100101101" => data_out <= rom_array(19245);
		when "0100101100101110" => data_out <= rom_array(19246);
		when "0100101100101111" => data_out <= rom_array(19247);
		when "0100101100110000" => data_out <= rom_array(19248);
		when "0100101100110001" => data_out <= rom_array(19249);
		when "0100101100110010" => data_out <= rom_array(19250);
		when "0100101100110011" => data_out <= rom_array(19251);
		when "0100101100110100" => data_out <= rom_array(19252);
		when "0100101100110101" => data_out <= rom_array(19253);
		when "0100101100110110" => data_out <= rom_array(19254);
		when "0100101100110111" => data_out <= rom_array(19255);
		when "0100101100111000" => data_out <= rom_array(19256);
		when "0100101100111001" => data_out <= rom_array(19257);
		when "0100101100111010" => data_out <= rom_array(19258);
		when "0100101100111011" => data_out <= rom_array(19259);
		when "0100101100111100" => data_out <= rom_array(19260);
		when "0100101100111101" => data_out <= rom_array(19261);
		when "0100101100111110" => data_out <= rom_array(19262);
		when "0100101100111111" => data_out <= rom_array(19263);
		when "0100101101000000" => data_out <= rom_array(19264);
		when "0100101101000001" => data_out <= rom_array(19265);
		when "0100101101000010" => data_out <= rom_array(19266);
		when "0100101101000011" => data_out <= rom_array(19267);
		when "0100101101000100" => data_out <= rom_array(19268);
		when "0100101101000101" => data_out <= rom_array(19269);
		when "0100101101000110" => data_out <= rom_array(19270);
		when "0100101101000111" => data_out <= rom_array(19271);
		when "0100101101001000" => data_out <= rom_array(19272);
		when "0100101101001001" => data_out <= rom_array(19273);
		when "0100101101001010" => data_out <= rom_array(19274);
		when "0100101101001011" => data_out <= rom_array(19275);
		when "0100101101001100" => data_out <= rom_array(19276);
		when "0100101101001101" => data_out <= rom_array(19277);
		when "0100101101001110" => data_out <= rom_array(19278);
		when "0100101101001111" => data_out <= rom_array(19279);
		when "0100101101010000" => data_out <= rom_array(19280);
		when "0100101101010001" => data_out <= rom_array(19281);
		when "0100101101010010" => data_out <= rom_array(19282);
		when "0100101101010011" => data_out <= rom_array(19283);
		when "0100101101010100" => data_out <= rom_array(19284);
		when "0100101101010101" => data_out <= rom_array(19285);
		when "0100101101010110" => data_out <= rom_array(19286);
		when "0100101101010111" => data_out <= rom_array(19287);
		when "0100101101011000" => data_out <= rom_array(19288);
		when "0100101101011001" => data_out <= rom_array(19289);
		when "0100101101011010" => data_out <= rom_array(19290);
		when "0100101101011011" => data_out <= rom_array(19291);
		when "0100101101011100" => data_out <= rom_array(19292);
		when "0100101101011101" => data_out <= rom_array(19293);
		when "0100101101011110" => data_out <= rom_array(19294);
		when "0100101101011111" => data_out <= rom_array(19295);
		when "0100101101100000" => data_out <= rom_array(19296);
		when "0100101101100001" => data_out <= rom_array(19297);
		when "0100101101100010" => data_out <= rom_array(19298);
		when "0100101101100011" => data_out <= rom_array(19299);
		when "0100101101100100" => data_out <= rom_array(19300);
		when "0100101101100101" => data_out <= rom_array(19301);
		when "0100101101100110" => data_out <= rom_array(19302);
		when "0100101101100111" => data_out <= rom_array(19303);
		when "0100101101101000" => data_out <= rom_array(19304);
		when "0100101101101001" => data_out <= rom_array(19305);
		when "0100101101101010" => data_out <= rom_array(19306);
		when "0100101101101011" => data_out <= rom_array(19307);
		when "0100101101101100" => data_out <= rom_array(19308);
		when "0100101101101101" => data_out <= rom_array(19309);
		when "0100101101101110" => data_out <= rom_array(19310);
		when "0100101101101111" => data_out <= rom_array(19311);
		when "0100101101110000" => data_out <= rom_array(19312);
		when "0100101101110001" => data_out <= rom_array(19313);
		when "0100101101110010" => data_out <= rom_array(19314);
		when "0100101101110011" => data_out <= rom_array(19315);
		when "0100101101110100" => data_out <= rom_array(19316);
		when "0100101101110101" => data_out <= rom_array(19317);
		when "0100101101110110" => data_out <= rom_array(19318);
		when "0100101101110111" => data_out <= rom_array(19319);
		when "0100101101111000" => data_out <= rom_array(19320);
		when "0100101101111001" => data_out <= rom_array(19321);
		when "0100101101111010" => data_out <= rom_array(19322);
		when "0100101101111011" => data_out <= rom_array(19323);
		when "0100101101111100" => data_out <= rom_array(19324);
		when "0100101101111101" => data_out <= rom_array(19325);
		when "0100101101111110" => data_out <= rom_array(19326);
		when "0100101101111111" => data_out <= rom_array(19327);
		when "0100101110000000" => data_out <= rom_array(19328);
		when "0100101110000001" => data_out <= rom_array(19329);
		when "0100101110000010" => data_out <= rom_array(19330);
		when "0100101110000011" => data_out <= rom_array(19331);
		when "0100101110000100" => data_out <= rom_array(19332);
		when "0100101110000101" => data_out <= rom_array(19333);
		when "0100101110000110" => data_out <= rom_array(19334);
		when "0100101110000111" => data_out <= rom_array(19335);
		when "0100101110001000" => data_out <= rom_array(19336);
		when "0100101110001001" => data_out <= rom_array(19337);
		when "0100101110001010" => data_out <= rom_array(19338);
		when "0100101110001011" => data_out <= rom_array(19339);
		when "0100101110001100" => data_out <= rom_array(19340);
		when "0100101110001101" => data_out <= rom_array(19341);
		when "0100101110001110" => data_out <= rom_array(19342);
		when "0100101110001111" => data_out <= rom_array(19343);
		when "0100101110010000" => data_out <= rom_array(19344);
		when "0100101110010001" => data_out <= rom_array(19345);
		when "0100101110010010" => data_out <= rom_array(19346);
		when "0100101110010011" => data_out <= rom_array(19347);
		when "0100101110010100" => data_out <= rom_array(19348);
		when "0100101110010101" => data_out <= rom_array(19349);
		when "0100101110010110" => data_out <= rom_array(19350);
		when "0100101110010111" => data_out <= rom_array(19351);
		when "0100101110011000" => data_out <= rom_array(19352);
		when "0100101110011001" => data_out <= rom_array(19353);
		when "0100101110011010" => data_out <= rom_array(19354);
		when "0100101110011011" => data_out <= rom_array(19355);
		when "0100101110011100" => data_out <= rom_array(19356);
		when "0100101110011101" => data_out <= rom_array(19357);
		when "0100101110011110" => data_out <= rom_array(19358);
		when "0100101110011111" => data_out <= rom_array(19359);
		when "0100101110100000" => data_out <= rom_array(19360);
		when "0100101110100001" => data_out <= rom_array(19361);
		when "0100101110100010" => data_out <= rom_array(19362);
		when "0100101110100011" => data_out <= rom_array(19363);
		when "0100101110100100" => data_out <= rom_array(19364);
		when "0100101110100101" => data_out <= rom_array(19365);
		when "0100101110100110" => data_out <= rom_array(19366);
		when "0100101110100111" => data_out <= rom_array(19367);
		when "0100101110101000" => data_out <= rom_array(19368);
		when "0100101110101001" => data_out <= rom_array(19369);
		when "0100101110101010" => data_out <= rom_array(19370);
		when "0100101110101011" => data_out <= rom_array(19371);
		when "0100101110101100" => data_out <= rom_array(19372);
		when "0100101110101101" => data_out <= rom_array(19373);
		when "0100101110101110" => data_out <= rom_array(19374);
		when "0100101110101111" => data_out <= rom_array(19375);
		when "0100101110110000" => data_out <= rom_array(19376);
		when "0100101110110001" => data_out <= rom_array(19377);
		when "0100101110110010" => data_out <= rom_array(19378);
		when "0100101110110011" => data_out <= rom_array(19379);
		when "0100101110110100" => data_out <= rom_array(19380);
		when "0100101110110101" => data_out <= rom_array(19381);
		when "0100101110110110" => data_out <= rom_array(19382);
		when "0100101110110111" => data_out <= rom_array(19383);
		when "0100101110111000" => data_out <= rom_array(19384);
		when "0100101110111001" => data_out <= rom_array(19385);
		when "0100101110111010" => data_out <= rom_array(19386);
		when "0100101110111011" => data_out <= rom_array(19387);
		when "0100101110111100" => data_out <= rom_array(19388);
		when "0100101110111101" => data_out <= rom_array(19389);
		when "0100101110111110" => data_out <= rom_array(19390);
		when "0100101110111111" => data_out <= rom_array(19391);
		when "0100101111000000" => data_out <= rom_array(19392);
		when "0100101111000001" => data_out <= rom_array(19393);
		when "0100101111000010" => data_out <= rom_array(19394);
		when "0100101111000011" => data_out <= rom_array(19395);
		when "0100101111000100" => data_out <= rom_array(19396);
		when "0100101111000101" => data_out <= rom_array(19397);
		when "0100101111000110" => data_out <= rom_array(19398);
		when "0100101111000111" => data_out <= rom_array(19399);
		when "0100101111001000" => data_out <= rom_array(19400);
		when "0100101111001001" => data_out <= rom_array(19401);
		when "0100101111001010" => data_out <= rom_array(19402);
		when "0100101111001011" => data_out <= rom_array(19403);
		when "0100101111001100" => data_out <= rom_array(19404);
		when "0100101111001101" => data_out <= rom_array(19405);
		when "0100101111001110" => data_out <= rom_array(19406);
		when "0100101111001111" => data_out <= rom_array(19407);
		when "0100101111010000" => data_out <= rom_array(19408);
		when "0100101111010001" => data_out <= rom_array(19409);
		when "0100101111010010" => data_out <= rom_array(19410);
		when "0100101111010011" => data_out <= rom_array(19411);
		when "0100101111010100" => data_out <= rom_array(19412);
		when "0100101111010101" => data_out <= rom_array(19413);
		when "0100101111010110" => data_out <= rom_array(19414);
		when "0100101111010111" => data_out <= rom_array(19415);
		when "0100101111011000" => data_out <= rom_array(19416);
		when "0100101111011001" => data_out <= rom_array(19417);
		when "0100101111011010" => data_out <= rom_array(19418);
		when "0100101111011011" => data_out <= rom_array(19419);
		when "0100101111011100" => data_out <= rom_array(19420);
		when "0100101111011101" => data_out <= rom_array(19421);
		when "0100101111011110" => data_out <= rom_array(19422);
		when "0100101111011111" => data_out <= rom_array(19423);
		when "0100101111100000" => data_out <= rom_array(19424);
		when "0100101111100001" => data_out <= rom_array(19425);
		when "0100101111100010" => data_out <= rom_array(19426);
		when "0100101111100011" => data_out <= rom_array(19427);
		when "0100101111100100" => data_out <= rom_array(19428);
		when "0100101111100101" => data_out <= rom_array(19429);
		when "0100101111100110" => data_out <= rom_array(19430);
		when "0100101111100111" => data_out <= rom_array(19431);
		when "0100101111101000" => data_out <= rom_array(19432);
		when "0100101111101001" => data_out <= rom_array(19433);
		when "0100101111101010" => data_out <= rom_array(19434);
		when "0100101111101011" => data_out <= rom_array(19435);
		when "0100101111101100" => data_out <= rom_array(19436);
		when "0100101111101101" => data_out <= rom_array(19437);
		when "0100101111101110" => data_out <= rom_array(19438);
		when "0100101111101111" => data_out <= rom_array(19439);
		when "0100101111110000" => data_out <= rom_array(19440);
		when "0100101111110001" => data_out <= rom_array(19441);
		when "0100101111110010" => data_out <= rom_array(19442);
		when "0100101111110011" => data_out <= rom_array(19443);
		when "0100101111110100" => data_out <= rom_array(19444);
		when "0100101111110101" => data_out <= rom_array(19445);
		when "0100101111110110" => data_out <= rom_array(19446);
		when "0100101111110111" => data_out <= rom_array(19447);
		when "0100101111111000" => data_out <= rom_array(19448);
		when "0100101111111001" => data_out <= rom_array(19449);
		when "0100101111111010" => data_out <= rom_array(19450);
		when "0100101111111011" => data_out <= rom_array(19451);
		when "0100101111111100" => data_out <= rom_array(19452);
		when "0100101111111101" => data_out <= rom_array(19453);
		when "0100101111111110" => data_out <= rom_array(19454);
		when "0100101111111111" => data_out <= rom_array(19455);
		when "0100110000000000" => data_out <= rom_array(19456);
		when "0100110000000001" => data_out <= rom_array(19457);
		when "0100110000000010" => data_out <= rom_array(19458);
		when "0100110000000011" => data_out <= rom_array(19459);
		when "0100110000000100" => data_out <= rom_array(19460);
		when "0100110000000101" => data_out <= rom_array(19461);
		when "0100110000000110" => data_out <= rom_array(19462);
		when "0100110000000111" => data_out <= rom_array(19463);
		when "0100110000001000" => data_out <= rom_array(19464);
		when "0100110000001001" => data_out <= rom_array(19465);
		when "0100110000001010" => data_out <= rom_array(19466);
		when "0100110000001011" => data_out <= rom_array(19467);
		when "0100110000001100" => data_out <= rom_array(19468);
		when "0100110000001101" => data_out <= rom_array(19469);
		when "0100110000001110" => data_out <= rom_array(19470);
		when "0100110000001111" => data_out <= rom_array(19471);
		when "0100110000010000" => data_out <= rom_array(19472);
		when "0100110000010001" => data_out <= rom_array(19473);
		when "0100110000010010" => data_out <= rom_array(19474);
		when "0100110000010011" => data_out <= rom_array(19475);
		when "0100110000010100" => data_out <= rom_array(19476);
		when "0100110000010101" => data_out <= rom_array(19477);
		when "0100110000010110" => data_out <= rom_array(19478);
		when "0100110000010111" => data_out <= rom_array(19479);
		when "0100110000011000" => data_out <= rom_array(19480);
		when "0100110000011001" => data_out <= rom_array(19481);
		when "0100110000011010" => data_out <= rom_array(19482);
		when "0100110000011011" => data_out <= rom_array(19483);
		when "0100110000011100" => data_out <= rom_array(19484);
		when "0100110000011101" => data_out <= rom_array(19485);
		when "0100110000011110" => data_out <= rom_array(19486);
		when "0100110000011111" => data_out <= rom_array(19487);
		when "0100110000100000" => data_out <= rom_array(19488);
		when "0100110000100001" => data_out <= rom_array(19489);
		when "0100110000100010" => data_out <= rom_array(19490);
		when "0100110000100011" => data_out <= rom_array(19491);
		when "0100110000100100" => data_out <= rom_array(19492);
		when "0100110000100101" => data_out <= rom_array(19493);
		when "0100110000100110" => data_out <= rom_array(19494);
		when "0100110000100111" => data_out <= rom_array(19495);
		when "0100110000101000" => data_out <= rom_array(19496);
		when "0100110000101001" => data_out <= rom_array(19497);
		when "0100110000101010" => data_out <= rom_array(19498);
		when "0100110000101011" => data_out <= rom_array(19499);
		when "0100110000101100" => data_out <= rom_array(19500);
		when "0100110000101101" => data_out <= rom_array(19501);
		when "0100110000101110" => data_out <= rom_array(19502);
		when "0100110000101111" => data_out <= rom_array(19503);
		when "0100110000110000" => data_out <= rom_array(19504);
		when "0100110000110001" => data_out <= rom_array(19505);
		when "0100110000110010" => data_out <= rom_array(19506);
		when "0100110000110011" => data_out <= rom_array(19507);
		when "0100110000110100" => data_out <= rom_array(19508);
		when "0100110000110101" => data_out <= rom_array(19509);
		when "0100110000110110" => data_out <= rom_array(19510);
		when "0100110000110111" => data_out <= rom_array(19511);
		when "0100110000111000" => data_out <= rom_array(19512);
		when "0100110000111001" => data_out <= rom_array(19513);
		when "0100110000111010" => data_out <= rom_array(19514);
		when "0100110000111011" => data_out <= rom_array(19515);
		when "0100110000111100" => data_out <= rom_array(19516);
		when "0100110000111101" => data_out <= rom_array(19517);
		when "0100110000111110" => data_out <= rom_array(19518);
		when "0100110000111111" => data_out <= rom_array(19519);
		when "0100110001000000" => data_out <= rom_array(19520);
		when "0100110001000001" => data_out <= rom_array(19521);
		when "0100110001000010" => data_out <= rom_array(19522);
		when "0100110001000011" => data_out <= rom_array(19523);
		when "0100110001000100" => data_out <= rom_array(19524);
		when "0100110001000101" => data_out <= rom_array(19525);
		when "0100110001000110" => data_out <= rom_array(19526);
		when "0100110001000111" => data_out <= rom_array(19527);
		when "0100110001001000" => data_out <= rom_array(19528);
		when "0100110001001001" => data_out <= rom_array(19529);
		when "0100110001001010" => data_out <= rom_array(19530);
		when "0100110001001011" => data_out <= rom_array(19531);
		when "0100110001001100" => data_out <= rom_array(19532);
		when "0100110001001101" => data_out <= rom_array(19533);
		when "0100110001001110" => data_out <= rom_array(19534);
		when "0100110001001111" => data_out <= rom_array(19535);
		when "0100110001010000" => data_out <= rom_array(19536);
		when "0100110001010001" => data_out <= rom_array(19537);
		when "0100110001010010" => data_out <= rom_array(19538);
		when "0100110001010011" => data_out <= rom_array(19539);
		when "0100110001010100" => data_out <= rom_array(19540);
		when "0100110001010101" => data_out <= rom_array(19541);
		when "0100110001010110" => data_out <= rom_array(19542);
		when "0100110001010111" => data_out <= rom_array(19543);
		when "0100110001011000" => data_out <= rom_array(19544);
		when "0100110001011001" => data_out <= rom_array(19545);
		when "0100110001011010" => data_out <= rom_array(19546);
		when "0100110001011011" => data_out <= rom_array(19547);
		when "0100110001011100" => data_out <= rom_array(19548);
		when "0100110001011101" => data_out <= rom_array(19549);
		when "0100110001011110" => data_out <= rom_array(19550);
		when "0100110001011111" => data_out <= rom_array(19551);
		when "0100110001100000" => data_out <= rom_array(19552);
		when "0100110001100001" => data_out <= rom_array(19553);
		when "0100110001100010" => data_out <= rom_array(19554);
		when "0100110001100011" => data_out <= rom_array(19555);
		when "0100110001100100" => data_out <= rom_array(19556);
		when "0100110001100101" => data_out <= rom_array(19557);
		when "0100110001100110" => data_out <= rom_array(19558);
		when "0100110001100111" => data_out <= rom_array(19559);
		when "0100110001101000" => data_out <= rom_array(19560);
		when "0100110001101001" => data_out <= rom_array(19561);
		when "0100110001101010" => data_out <= rom_array(19562);
		when "0100110001101011" => data_out <= rom_array(19563);
		when "0100110001101100" => data_out <= rom_array(19564);
		when "0100110001101101" => data_out <= rom_array(19565);
		when "0100110001101110" => data_out <= rom_array(19566);
		when "0100110001101111" => data_out <= rom_array(19567);
		when "0100110001110000" => data_out <= rom_array(19568);
		when "0100110001110001" => data_out <= rom_array(19569);
		when "0100110001110010" => data_out <= rom_array(19570);
		when "0100110001110011" => data_out <= rom_array(19571);
		when "0100110001110100" => data_out <= rom_array(19572);
		when "0100110001110101" => data_out <= rom_array(19573);
		when "0100110001110110" => data_out <= rom_array(19574);
		when "0100110001110111" => data_out <= rom_array(19575);
		when "0100110001111000" => data_out <= rom_array(19576);
		when "0100110001111001" => data_out <= rom_array(19577);
		when "0100110001111010" => data_out <= rom_array(19578);
		when "0100110001111011" => data_out <= rom_array(19579);
		when "0100110001111100" => data_out <= rom_array(19580);
		when "0100110001111101" => data_out <= rom_array(19581);
		when "0100110001111110" => data_out <= rom_array(19582);
		when "0100110001111111" => data_out <= rom_array(19583);
		when "0100110010000000" => data_out <= rom_array(19584);
		when "0100110010000001" => data_out <= rom_array(19585);
		when "0100110010000010" => data_out <= rom_array(19586);
		when "0100110010000011" => data_out <= rom_array(19587);
		when "0100110010000100" => data_out <= rom_array(19588);
		when "0100110010000101" => data_out <= rom_array(19589);
		when "0100110010000110" => data_out <= rom_array(19590);
		when "0100110010000111" => data_out <= rom_array(19591);
		when "0100110010001000" => data_out <= rom_array(19592);
		when "0100110010001001" => data_out <= rom_array(19593);
		when "0100110010001010" => data_out <= rom_array(19594);
		when "0100110010001011" => data_out <= rom_array(19595);
		when "0100110010001100" => data_out <= rom_array(19596);
		when "0100110010001101" => data_out <= rom_array(19597);
		when "0100110010001110" => data_out <= rom_array(19598);
		when "0100110010001111" => data_out <= rom_array(19599);
		when "0100110010010000" => data_out <= rom_array(19600);
		when "0100110010010001" => data_out <= rom_array(19601);
		when "0100110010010010" => data_out <= rom_array(19602);
		when "0100110010010011" => data_out <= rom_array(19603);
		when "0100110010010100" => data_out <= rom_array(19604);
		when "0100110010010101" => data_out <= rom_array(19605);
		when "0100110010010110" => data_out <= rom_array(19606);
		when "0100110010010111" => data_out <= rom_array(19607);
		when "0100110010011000" => data_out <= rom_array(19608);
		when "0100110010011001" => data_out <= rom_array(19609);
		when "0100110010011010" => data_out <= rom_array(19610);
		when "0100110010011011" => data_out <= rom_array(19611);
		when "0100110010011100" => data_out <= rom_array(19612);
		when "0100110010011101" => data_out <= rom_array(19613);
		when "0100110010011110" => data_out <= rom_array(19614);
		when "0100110010011111" => data_out <= rom_array(19615);
		when "0100110010100000" => data_out <= rom_array(19616);
		when "0100110010100001" => data_out <= rom_array(19617);
		when "0100110010100010" => data_out <= rom_array(19618);
		when "0100110010100011" => data_out <= rom_array(19619);
		when "0100110010100100" => data_out <= rom_array(19620);
		when "0100110010100101" => data_out <= rom_array(19621);
		when "0100110010100110" => data_out <= rom_array(19622);
		when "0100110010100111" => data_out <= rom_array(19623);
		when "0100110010101000" => data_out <= rom_array(19624);
		when "0100110010101001" => data_out <= rom_array(19625);
		when "0100110010101010" => data_out <= rom_array(19626);
		when "0100110010101011" => data_out <= rom_array(19627);
		when "0100110010101100" => data_out <= rom_array(19628);
		when "0100110010101101" => data_out <= rom_array(19629);
		when "0100110010101110" => data_out <= rom_array(19630);
		when "0100110010101111" => data_out <= rom_array(19631);
		when "0100110010110000" => data_out <= rom_array(19632);
		when "0100110010110001" => data_out <= rom_array(19633);
		when "0100110010110010" => data_out <= rom_array(19634);
		when "0100110010110011" => data_out <= rom_array(19635);
		when "0100110010110100" => data_out <= rom_array(19636);
		when "0100110010110101" => data_out <= rom_array(19637);
		when "0100110010110110" => data_out <= rom_array(19638);
		when "0100110010110111" => data_out <= rom_array(19639);
		when "0100110010111000" => data_out <= rom_array(19640);
		when "0100110010111001" => data_out <= rom_array(19641);
		when "0100110010111010" => data_out <= rom_array(19642);
		when "0100110010111011" => data_out <= rom_array(19643);
		when "0100110010111100" => data_out <= rom_array(19644);
		when "0100110010111101" => data_out <= rom_array(19645);
		when "0100110010111110" => data_out <= rom_array(19646);
		when "0100110010111111" => data_out <= rom_array(19647);
		when "0100110011000000" => data_out <= rom_array(19648);
		when "0100110011000001" => data_out <= rom_array(19649);
		when "0100110011000010" => data_out <= rom_array(19650);
		when "0100110011000011" => data_out <= rom_array(19651);
		when "0100110011000100" => data_out <= rom_array(19652);
		when "0100110011000101" => data_out <= rom_array(19653);
		when "0100110011000110" => data_out <= rom_array(19654);
		when "0100110011000111" => data_out <= rom_array(19655);
		when "0100110011001000" => data_out <= rom_array(19656);
		when "0100110011001001" => data_out <= rom_array(19657);
		when "0100110011001010" => data_out <= rom_array(19658);
		when "0100110011001011" => data_out <= rom_array(19659);
		when "0100110011001100" => data_out <= rom_array(19660);
		when "0100110011001101" => data_out <= rom_array(19661);
		when "0100110011001110" => data_out <= rom_array(19662);
		when "0100110011001111" => data_out <= rom_array(19663);
		when "0100110011010000" => data_out <= rom_array(19664);
		when "0100110011010001" => data_out <= rom_array(19665);
		when "0100110011010010" => data_out <= rom_array(19666);
		when "0100110011010011" => data_out <= rom_array(19667);
		when "0100110011010100" => data_out <= rom_array(19668);
		when "0100110011010101" => data_out <= rom_array(19669);
		when "0100110011010110" => data_out <= rom_array(19670);
		when "0100110011010111" => data_out <= rom_array(19671);
		when "0100110011011000" => data_out <= rom_array(19672);
		when "0100110011011001" => data_out <= rom_array(19673);
		when "0100110011011010" => data_out <= rom_array(19674);
		when "0100110011011011" => data_out <= rom_array(19675);
		when "0100110011011100" => data_out <= rom_array(19676);
		when "0100110011011101" => data_out <= rom_array(19677);
		when "0100110011011110" => data_out <= rom_array(19678);
		when "0100110011011111" => data_out <= rom_array(19679);
		when "0100110011100000" => data_out <= rom_array(19680);
		when "0100110011100001" => data_out <= rom_array(19681);
		when "0100110011100010" => data_out <= rom_array(19682);
		when "0100110011100011" => data_out <= rom_array(19683);
		when "0100110011100100" => data_out <= rom_array(19684);
		when "0100110011100101" => data_out <= rom_array(19685);
		when "0100110011100110" => data_out <= rom_array(19686);
		when "0100110011100111" => data_out <= rom_array(19687);
		when "0100110011101000" => data_out <= rom_array(19688);
		when "0100110011101001" => data_out <= rom_array(19689);
		when "0100110011101010" => data_out <= rom_array(19690);
		when "0100110011101011" => data_out <= rom_array(19691);
		when "0100110011101100" => data_out <= rom_array(19692);
		when "0100110011101101" => data_out <= rom_array(19693);
		when "0100110011101110" => data_out <= rom_array(19694);
		when "0100110011101111" => data_out <= rom_array(19695);
		when "0100110011110000" => data_out <= rom_array(19696);
		when "0100110011110001" => data_out <= rom_array(19697);
		when "0100110011110010" => data_out <= rom_array(19698);
		when "0100110011110011" => data_out <= rom_array(19699);
		when "0100110011110100" => data_out <= rom_array(19700);
		when "0100110011110101" => data_out <= rom_array(19701);
		when "0100110011110110" => data_out <= rom_array(19702);
		when "0100110011110111" => data_out <= rom_array(19703);
		when "0100110011111000" => data_out <= rom_array(19704);
		when "0100110011111001" => data_out <= rom_array(19705);
		when "0100110011111010" => data_out <= rom_array(19706);
		when "0100110011111011" => data_out <= rom_array(19707);
		when "0100110011111100" => data_out <= rom_array(19708);
		when "0100110011111101" => data_out <= rom_array(19709);
		when "0100110011111110" => data_out <= rom_array(19710);
		when "0100110011111111" => data_out <= rom_array(19711);
		when "0100110100000000" => data_out <= rom_array(19712);
		when "0100110100000001" => data_out <= rom_array(19713);
		when "0100110100000010" => data_out <= rom_array(19714);
		when "0100110100000011" => data_out <= rom_array(19715);
		when "0100110100000100" => data_out <= rom_array(19716);
		when "0100110100000101" => data_out <= rom_array(19717);
		when "0100110100000110" => data_out <= rom_array(19718);
		when "0100110100000111" => data_out <= rom_array(19719);
		when "0100110100001000" => data_out <= rom_array(19720);
		when "0100110100001001" => data_out <= rom_array(19721);
		when "0100110100001010" => data_out <= rom_array(19722);
		when "0100110100001011" => data_out <= rom_array(19723);
		when "0100110100001100" => data_out <= rom_array(19724);
		when "0100110100001101" => data_out <= rom_array(19725);
		when "0100110100001110" => data_out <= rom_array(19726);
		when "0100110100001111" => data_out <= rom_array(19727);
		when "0100110100010000" => data_out <= rom_array(19728);
		when "0100110100010001" => data_out <= rom_array(19729);
		when "0100110100010010" => data_out <= rom_array(19730);
		when "0100110100010011" => data_out <= rom_array(19731);
		when "0100110100010100" => data_out <= rom_array(19732);
		when "0100110100010101" => data_out <= rom_array(19733);
		when "0100110100010110" => data_out <= rom_array(19734);
		when "0100110100010111" => data_out <= rom_array(19735);
		when "0100110100011000" => data_out <= rom_array(19736);
		when "0100110100011001" => data_out <= rom_array(19737);
		when "0100110100011010" => data_out <= rom_array(19738);
		when "0100110100011011" => data_out <= rom_array(19739);
		when "0100110100011100" => data_out <= rom_array(19740);
		when "0100110100011101" => data_out <= rom_array(19741);
		when "0100110100011110" => data_out <= rom_array(19742);
		when "0100110100011111" => data_out <= rom_array(19743);
		when "0100110100100000" => data_out <= rom_array(19744);
		when "0100110100100001" => data_out <= rom_array(19745);
		when "0100110100100010" => data_out <= rom_array(19746);
		when "0100110100100011" => data_out <= rom_array(19747);
		when "0100110100100100" => data_out <= rom_array(19748);
		when "0100110100100101" => data_out <= rom_array(19749);
		when "0100110100100110" => data_out <= rom_array(19750);
		when "0100110100100111" => data_out <= rom_array(19751);
		when "0100110100101000" => data_out <= rom_array(19752);
		when "0100110100101001" => data_out <= rom_array(19753);
		when "0100110100101010" => data_out <= rom_array(19754);
		when "0100110100101011" => data_out <= rom_array(19755);
		when "0100110100101100" => data_out <= rom_array(19756);
		when "0100110100101101" => data_out <= rom_array(19757);
		when "0100110100101110" => data_out <= rom_array(19758);
		when "0100110100101111" => data_out <= rom_array(19759);
		when "0100110100110000" => data_out <= rom_array(19760);
		when "0100110100110001" => data_out <= rom_array(19761);
		when "0100110100110010" => data_out <= rom_array(19762);
		when "0100110100110011" => data_out <= rom_array(19763);
		when "0100110100110100" => data_out <= rom_array(19764);
		when "0100110100110101" => data_out <= rom_array(19765);
		when "0100110100110110" => data_out <= rom_array(19766);
		when "0100110100110111" => data_out <= rom_array(19767);
		when "0100110100111000" => data_out <= rom_array(19768);
		when "0100110100111001" => data_out <= rom_array(19769);
		when "0100110100111010" => data_out <= rom_array(19770);
		when "0100110100111011" => data_out <= rom_array(19771);
		when "0100110100111100" => data_out <= rom_array(19772);
		when "0100110100111101" => data_out <= rom_array(19773);
		when "0100110100111110" => data_out <= rom_array(19774);
		when "0100110100111111" => data_out <= rom_array(19775);
		when "0100110101000000" => data_out <= rom_array(19776);
		when "0100110101000001" => data_out <= rom_array(19777);
		when "0100110101000010" => data_out <= rom_array(19778);
		when "0100110101000011" => data_out <= rom_array(19779);
		when "0100110101000100" => data_out <= rom_array(19780);
		when "0100110101000101" => data_out <= rom_array(19781);
		when "0100110101000110" => data_out <= rom_array(19782);
		when "0100110101000111" => data_out <= rom_array(19783);
		when "0100110101001000" => data_out <= rom_array(19784);
		when "0100110101001001" => data_out <= rom_array(19785);
		when "0100110101001010" => data_out <= rom_array(19786);
		when "0100110101001011" => data_out <= rom_array(19787);
		when "0100110101001100" => data_out <= rom_array(19788);
		when "0100110101001101" => data_out <= rom_array(19789);
		when "0100110101001110" => data_out <= rom_array(19790);
		when "0100110101001111" => data_out <= rom_array(19791);
		when "0100110101010000" => data_out <= rom_array(19792);
		when "0100110101010001" => data_out <= rom_array(19793);
		when "0100110101010010" => data_out <= rom_array(19794);
		when "0100110101010011" => data_out <= rom_array(19795);
		when "0100110101010100" => data_out <= rom_array(19796);
		when "0100110101010101" => data_out <= rom_array(19797);
		when "0100110101010110" => data_out <= rom_array(19798);
		when "0100110101010111" => data_out <= rom_array(19799);
		when "0100110101011000" => data_out <= rom_array(19800);
		when "0100110101011001" => data_out <= rom_array(19801);
		when "0100110101011010" => data_out <= rom_array(19802);
		when "0100110101011011" => data_out <= rom_array(19803);
		when "0100110101011100" => data_out <= rom_array(19804);
		when "0100110101011101" => data_out <= rom_array(19805);
		when "0100110101011110" => data_out <= rom_array(19806);
		when "0100110101011111" => data_out <= rom_array(19807);
		when "0100110101100000" => data_out <= rom_array(19808);
		when "0100110101100001" => data_out <= rom_array(19809);
		when "0100110101100010" => data_out <= rom_array(19810);
		when "0100110101100011" => data_out <= rom_array(19811);
		when "0100110101100100" => data_out <= rom_array(19812);
		when "0100110101100101" => data_out <= rom_array(19813);
		when "0100110101100110" => data_out <= rom_array(19814);
		when "0100110101100111" => data_out <= rom_array(19815);
		when "0100110101101000" => data_out <= rom_array(19816);
		when "0100110101101001" => data_out <= rom_array(19817);
		when "0100110101101010" => data_out <= rom_array(19818);
		when "0100110101101011" => data_out <= rom_array(19819);
		when "0100110101101100" => data_out <= rom_array(19820);
		when "0100110101101101" => data_out <= rom_array(19821);
		when "0100110101101110" => data_out <= rom_array(19822);
		when "0100110101101111" => data_out <= rom_array(19823);
		when "0100110101110000" => data_out <= rom_array(19824);
		when "0100110101110001" => data_out <= rom_array(19825);
		when "0100110101110010" => data_out <= rom_array(19826);
		when "0100110101110011" => data_out <= rom_array(19827);
		when "0100110101110100" => data_out <= rom_array(19828);
		when "0100110101110101" => data_out <= rom_array(19829);
		when "0100110101110110" => data_out <= rom_array(19830);
		when "0100110101110111" => data_out <= rom_array(19831);
		when "0100110101111000" => data_out <= rom_array(19832);
		when "0100110101111001" => data_out <= rom_array(19833);
		when "0100110101111010" => data_out <= rom_array(19834);
		when "0100110101111011" => data_out <= rom_array(19835);
		when "0100110101111100" => data_out <= rom_array(19836);
		when "0100110101111101" => data_out <= rom_array(19837);
		when "0100110101111110" => data_out <= rom_array(19838);
		when "0100110101111111" => data_out <= rom_array(19839);
		when "0100110110000000" => data_out <= rom_array(19840);
		when "0100110110000001" => data_out <= rom_array(19841);
		when "0100110110000010" => data_out <= rom_array(19842);
		when "0100110110000011" => data_out <= rom_array(19843);
		when "0100110110000100" => data_out <= rom_array(19844);
		when "0100110110000101" => data_out <= rom_array(19845);
		when "0100110110000110" => data_out <= rom_array(19846);
		when "0100110110000111" => data_out <= rom_array(19847);
		when "0100110110001000" => data_out <= rom_array(19848);
		when "0100110110001001" => data_out <= rom_array(19849);
		when "0100110110001010" => data_out <= rom_array(19850);
		when "0100110110001011" => data_out <= rom_array(19851);
		when "0100110110001100" => data_out <= rom_array(19852);
		when "0100110110001101" => data_out <= rom_array(19853);
		when "0100110110001110" => data_out <= rom_array(19854);
		when "0100110110001111" => data_out <= rom_array(19855);
		when "0100110110010000" => data_out <= rom_array(19856);
		when "0100110110010001" => data_out <= rom_array(19857);
		when "0100110110010010" => data_out <= rom_array(19858);
		when "0100110110010011" => data_out <= rom_array(19859);
		when "0100110110010100" => data_out <= rom_array(19860);
		when "0100110110010101" => data_out <= rom_array(19861);
		when "0100110110010110" => data_out <= rom_array(19862);
		when "0100110110010111" => data_out <= rom_array(19863);
		when "0100110110011000" => data_out <= rom_array(19864);
		when "0100110110011001" => data_out <= rom_array(19865);
		when "0100110110011010" => data_out <= rom_array(19866);
		when "0100110110011011" => data_out <= rom_array(19867);
		when "0100110110011100" => data_out <= rom_array(19868);
		when "0100110110011101" => data_out <= rom_array(19869);
		when "0100110110011110" => data_out <= rom_array(19870);
		when "0100110110011111" => data_out <= rom_array(19871);
		when "0100110110100000" => data_out <= rom_array(19872);
		when "0100110110100001" => data_out <= rom_array(19873);
		when "0100110110100010" => data_out <= rom_array(19874);
		when "0100110110100011" => data_out <= rom_array(19875);
		when "0100110110100100" => data_out <= rom_array(19876);
		when "0100110110100101" => data_out <= rom_array(19877);
		when "0100110110100110" => data_out <= rom_array(19878);
		when "0100110110100111" => data_out <= rom_array(19879);
		when "0100110110101000" => data_out <= rom_array(19880);
		when "0100110110101001" => data_out <= rom_array(19881);
		when "0100110110101010" => data_out <= rom_array(19882);
		when "0100110110101011" => data_out <= rom_array(19883);
		when "0100110110101100" => data_out <= rom_array(19884);
		when "0100110110101101" => data_out <= rom_array(19885);
		when "0100110110101110" => data_out <= rom_array(19886);
		when "0100110110101111" => data_out <= rom_array(19887);
		when "0100110110110000" => data_out <= rom_array(19888);
		when "0100110110110001" => data_out <= rom_array(19889);
		when "0100110110110010" => data_out <= rom_array(19890);
		when "0100110110110011" => data_out <= rom_array(19891);
		when "0100110110110100" => data_out <= rom_array(19892);
		when "0100110110110101" => data_out <= rom_array(19893);
		when "0100110110110110" => data_out <= rom_array(19894);
		when "0100110110110111" => data_out <= rom_array(19895);
		when "0100110110111000" => data_out <= rom_array(19896);
		when "0100110110111001" => data_out <= rom_array(19897);
		when "0100110110111010" => data_out <= rom_array(19898);
		when "0100110110111011" => data_out <= rom_array(19899);
		when "0100110110111100" => data_out <= rom_array(19900);
		when "0100110110111101" => data_out <= rom_array(19901);
		when "0100110110111110" => data_out <= rom_array(19902);
		when "0100110110111111" => data_out <= rom_array(19903);
		when "0100110111000000" => data_out <= rom_array(19904);
		when "0100110111000001" => data_out <= rom_array(19905);
		when "0100110111000010" => data_out <= rom_array(19906);
		when "0100110111000011" => data_out <= rom_array(19907);
		when "0100110111000100" => data_out <= rom_array(19908);
		when "0100110111000101" => data_out <= rom_array(19909);
		when "0100110111000110" => data_out <= rom_array(19910);
		when "0100110111000111" => data_out <= rom_array(19911);
		when "0100110111001000" => data_out <= rom_array(19912);
		when "0100110111001001" => data_out <= rom_array(19913);
		when "0100110111001010" => data_out <= rom_array(19914);
		when "0100110111001011" => data_out <= rom_array(19915);
		when "0100110111001100" => data_out <= rom_array(19916);
		when "0100110111001101" => data_out <= rom_array(19917);
		when "0100110111001110" => data_out <= rom_array(19918);
		when "0100110111001111" => data_out <= rom_array(19919);
		when "0100110111010000" => data_out <= rom_array(19920);
		when "0100110111010001" => data_out <= rom_array(19921);
		when "0100110111010010" => data_out <= rom_array(19922);
		when "0100110111010011" => data_out <= rom_array(19923);
		when "0100110111010100" => data_out <= rom_array(19924);
		when "0100110111010101" => data_out <= rom_array(19925);
		when "0100110111010110" => data_out <= rom_array(19926);
		when "0100110111010111" => data_out <= rom_array(19927);
		when "0100110111011000" => data_out <= rom_array(19928);
		when "0100110111011001" => data_out <= rom_array(19929);
		when "0100110111011010" => data_out <= rom_array(19930);
		when "0100110111011011" => data_out <= rom_array(19931);
		when "0100110111011100" => data_out <= rom_array(19932);
		when "0100110111011101" => data_out <= rom_array(19933);
		when "0100110111011110" => data_out <= rom_array(19934);
		when "0100110111011111" => data_out <= rom_array(19935);
		when "0100110111100000" => data_out <= rom_array(19936);
		when "0100110111100001" => data_out <= rom_array(19937);
		when "0100110111100010" => data_out <= rom_array(19938);
		when "0100110111100011" => data_out <= rom_array(19939);
		when "0100110111100100" => data_out <= rom_array(19940);
		when "0100110111100101" => data_out <= rom_array(19941);
		when "0100110111100110" => data_out <= rom_array(19942);
		when "0100110111100111" => data_out <= rom_array(19943);
		when "0100110111101000" => data_out <= rom_array(19944);
		when "0100110111101001" => data_out <= rom_array(19945);
		when "0100110111101010" => data_out <= rom_array(19946);
		when "0100110111101011" => data_out <= rom_array(19947);
		when "0100110111101100" => data_out <= rom_array(19948);
		when "0100110111101101" => data_out <= rom_array(19949);
		when "0100110111101110" => data_out <= rom_array(19950);
		when "0100110111101111" => data_out <= rom_array(19951);
		when "0100110111110000" => data_out <= rom_array(19952);
		when "0100110111110001" => data_out <= rom_array(19953);
		when "0100110111110010" => data_out <= rom_array(19954);
		when "0100110111110011" => data_out <= rom_array(19955);
		when "0100110111110100" => data_out <= rom_array(19956);
		when "0100110111110101" => data_out <= rom_array(19957);
		when "0100110111110110" => data_out <= rom_array(19958);
		when "0100110111110111" => data_out <= rom_array(19959);
		when "0100110111111000" => data_out <= rom_array(19960);
		when "0100110111111001" => data_out <= rom_array(19961);
		when "0100110111111010" => data_out <= rom_array(19962);
		when "0100110111111011" => data_out <= rom_array(19963);
		when "0100110111111100" => data_out <= rom_array(19964);
		when "0100110111111101" => data_out <= rom_array(19965);
		when "0100110111111110" => data_out <= rom_array(19966);
		when "0100110111111111" => data_out <= rom_array(19967);
		when "0100111000000000" => data_out <= rom_array(19968);
		when "0100111000000001" => data_out <= rom_array(19969);
		when "0100111000000010" => data_out <= rom_array(19970);
		when "0100111000000011" => data_out <= rom_array(19971);
		when "0100111000000100" => data_out <= rom_array(19972);
		when "0100111000000101" => data_out <= rom_array(19973);
		when "0100111000000110" => data_out <= rom_array(19974);
		when "0100111000000111" => data_out <= rom_array(19975);
		when "0100111000001000" => data_out <= rom_array(19976);
		when "0100111000001001" => data_out <= rom_array(19977);
		when "0100111000001010" => data_out <= rom_array(19978);
		when "0100111000001011" => data_out <= rom_array(19979);
		when "0100111000001100" => data_out <= rom_array(19980);
		when "0100111000001101" => data_out <= rom_array(19981);
		when "0100111000001110" => data_out <= rom_array(19982);
		when "0100111000001111" => data_out <= rom_array(19983);
		when "0100111000010000" => data_out <= rom_array(19984);
		when "0100111000010001" => data_out <= rom_array(19985);
		when "0100111000010010" => data_out <= rom_array(19986);
		when "0100111000010011" => data_out <= rom_array(19987);
		when "0100111000010100" => data_out <= rom_array(19988);
		when "0100111000010101" => data_out <= rom_array(19989);
		when "0100111000010110" => data_out <= rom_array(19990);
		when "0100111000010111" => data_out <= rom_array(19991);
		when "0100111000011000" => data_out <= rom_array(19992);
		when "0100111000011001" => data_out <= rom_array(19993);
		when "0100111000011010" => data_out <= rom_array(19994);
		when "0100111000011011" => data_out <= rom_array(19995);
		when "0100111000011100" => data_out <= rom_array(19996);
		when "0100111000011101" => data_out <= rom_array(19997);
		when "0100111000011110" => data_out <= rom_array(19998);
		when "0100111000011111" => data_out <= rom_array(19999);
		when "0100111000100000" => data_out <= rom_array(20000);
		when "0100111000100001" => data_out <= rom_array(20001);
		when "0100111000100010" => data_out <= rom_array(20002);
		when "0100111000100011" => data_out <= rom_array(20003);
		when "0100111000100100" => data_out <= rom_array(20004);
		when "0100111000100101" => data_out <= rom_array(20005);
		when "0100111000100110" => data_out <= rom_array(20006);
		when "0100111000100111" => data_out <= rom_array(20007);
		when "0100111000101000" => data_out <= rom_array(20008);
		when "0100111000101001" => data_out <= rom_array(20009);
		when "0100111000101010" => data_out <= rom_array(20010);
		when "0100111000101011" => data_out <= rom_array(20011);
		when "0100111000101100" => data_out <= rom_array(20012);
		when "0100111000101101" => data_out <= rom_array(20013);
		when "0100111000101110" => data_out <= rom_array(20014);
		when "0100111000101111" => data_out <= rom_array(20015);
		when "0100111000110000" => data_out <= rom_array(20016);
		when "0100111000110001" => data_out <= rom_array(20017);
		when "0100111000110010" => data_out <= rom_array(20018);
		when "0100111000110011" => data_out <= rom_array(20019);
		when "0100111000110100" => data_out <= rom_array(20020);
		when "0100111000110101" => data_out <= rom_array(20021);
		when "0100111000110110" => data_out <= rom_array(20022);
		when "0100111000110111" => data_out <= rom_array(20023);
		when "0100111000111000" => data_out <= rom_array(20024);
		when "0100111000111001" => data_out <= rom_array(20025);
		when "0100111000111010" => data_out <= rom_array(20026);
		when "0100111000111011" => data_out <= rom_array(20027);
		when "0100111000111100" => data_out <= rom_array(20028);
		when "0100111000111101" => data_out <= rom_array(20029);
		when "0100111000111110" => data_out <= rom_array(20030);
		when "0100111000111111" => data_out <= rom_array(20031);
		when "0100111001000000" => data_out <= rom_array(20032);
		when "0100111001000001" => data_out <= rom_array(20033);
		when "0100111001000010" => data_out <= rom_array(20034);
		when "0100111001000011" => data_out <= rom_array(20035);
		when "0100111001000100" => data_out <= rom_array(20036);
		when "0100111001000101" => data_out <= rom_array(20037);
		when "0100111001000110" => data_out <= rom_array(20038);
		when "0100111001000111" => data_out <= rom_array(20039);
		when "0100111001001000" => data_out <= rom_array(20040);
		when "0100111001001001" => data_out <= rom_array(20041);
		when "0100111001001010" => data_out <= rom_array(20042);
		when "0100111001001011" => data_out <= rom_array(20043);
		when "0100111001001100" => data_out <= rom_array(20044);
		when "0100111001001101" => data_out <= rom_array(20045);
		when "0100111001001110" => data_out <= rom_array(20046);
		when "0100111001001111" => data_out <= rom_array(20047);
		when "0100111001010000" => data_out <= rom_array(20048);
		when "0100111001010001" => data_out <= rom_array(20049);
		when "0100111001010010" => data_out <= rom_array(20050);
		when "0100111001010011" => data_out <= rom_array(20051);
		when "0100111001010100" => data_out <= rom_array(20052);
		when "0100111001010101" => data_out <= rom_array(20053);
		when "0100111001010110" => data_out <= rom_array(20054);
		when "0100111001010111" => data_out <= rom_array(20055);
		when "0100111001011000" => data_out <= rom_array(20056);
		when "0100111001011001" => data_out <= rom_array(20057);
		when "0100111001011010" => data_out <= rom_array(20058);
		when "0100111001011011" => data_out <= rom_array(20059);
		when "0100111001011100" => data_out <= rom_array(20060);
		when "0100111001011101" => data_out <= rom_array(20061);
		when "0100111001011110" => data_out <= rom_array(20062);
		when "0100111001011111" => data_out <= rom_array(20063);
		when "0100111001100000" => data_out <= rom_array(20064);
		when "0100111001100001" => data_out <= rom_array(20065);
		when "0100111001100010" => data_out <= rom_array(20066);
		when "0100111001100011" => data_out <= rom_array(20067);
		when "0100111001100100" => data_out <= rom_array(20068);
		when "0100111001100101" => data_out <= rom_array(20069);
		when "0100111001100110" => data_out <= rom_array(20070);
		when "0100111001100111" => data_out <= rom_array(20071);
		when "0100111001101000" => data_out <= rom_array(20072);
		when "0100111001101001" => data_out <= rom_array(20073);
		when "0100111001101010" => data_out <= rom_array(20074);
		when "0100111001101011" => data_out <= rom_array(20075);
		when "0100111001101100" => data_out <= rom_array(20076);
		when "0100111001101101" => data_out <= rom_array(20077);
		when "0100111001101110" => data_out <= rom_array(20078);
		when "0100111001101111" => data_out <= rom_array(20079);
		when "0100111001110000" => data_out <= rom_array(20080);
		when "0100111001110001" => data_out <= rom_array(20081);
		when "0100111001110010" => data_out <= rom_array(20082);
		when "0100111001110011" => data_out <= rom_array(20083);
		when "0100111001110100" => data_out <= rom_array(20084);
		when "0100111001110101" => data_out <= rom_array(20085);
		when "0100111001110110" => data_out <= rom_array(20086);
		when "0100111001110111" => data_out <= rom_array(20087);
		when "0100111001111000" => data_out <= rom_array(20088);
		when "0100111001111001" => data_out <= rom_array(20089);
		when "0100111001111010" => data_out <= rom_array(20090);
		when "0100111001111011" => data_out <= rom_array(20091);
		when "0100111001111100" => data_out <= rom_array(20092);
		when "0100111001111101" => data_out <= rom_array(20093);
		when "0100111001111110" => data_out <= rom_array(20094);
		when "0100111001111111" => data_out <= rom_array(20095);
		when "0100111010000000" => data_out <= rom_array(20096);
		when "0100111010000001" => data_out <= rom_array(20097);
		when "0100111010000010" => data_out <= rom_array(20098);
		when "0100111010000011" => data_out <= rom_array(20099);
		when "0100111010000100" => data_out <= rom_array(20100);
		when "0100111010000101" => data_out <= rom_array(20101);
		when "0100111010000110" => data_out <= rom_array(20102);
		when "0100111010000111" => data_out <= rom_array(20103);
		when "0100111010001000" => data_out <= rom_array(20104);
		when "0100111010001001" => data_out <= rom_array(20105);
		when "0100111010001010" => data_out <= rom_array(20106);
		when "0100111010001011" => data_out <= rom_array(20107);
		when "0100111010001100" => data_out <= rom_array(20108);
		when "0100111010001101" => data_out <= rom_array(20109);
		when "0100111010001110" => data_out <= rom_array(20110);
		when "0100111010001111" => data_out <= rom_array(20111);
		when "0100111010010000" => data_out <= rom_array(20112);
		when "0100111010010001" => data_out <= rom_array(20113);
		when "0100111010010010" => data_out <= rom_array(20114);
		when "0100111010010011" => data_out <= rom_array(20115);
		when "0100111010010100" => data_out <= rom_array(20116);
		when "0100111010010101" => data_out <= rom_array(20117);
		when "0100111010010110" => data_out <= rom_array(20118);
		when "0100111010010111" => data_out <= rom_array(20119);
		when "0100111010011000" => data_out <= rom_array(20120);
		when "0100111010011001" => data_out <= rom_array(20121);
		when "0100111010011010" => data_out <= rom_array(20122);
		when "0100111010011011" => data_out <= rom_array(20123);
		when "0100111010011100" => data_out <= rom_array(20124);
		when "0100111010011101" => data_out <= rom_array(20125);
		when "0100111010011110" => data_out <= rom_array(20126);
		when "0100111010011111" => data_out <= rom_array(20127);
		when "0100111010100000" => data_out <= rom_array(20128);
		when "0100111010100001" => data_out <= rom_array(20129);
		when "0100111010100010" => data_out <= rom_array(20130);
		when "0100111010100011" => data_out <= rom_array(20131);
		when "0100111010100100" => data_out <= rom_array(20132);
		when "0100111010100101" => data_out <= rom_array(20133);
		when "0100111010100110" => data_out <= rom_array(20134);
		when "0100111010100111" => data_out <= rom_array(20135);
		when "0100111010101000" => data_out <= rom_array(20136);
		when "0100111010101001" => data_out <= rom_array(20137);
		when "0100111010101010" => data_out <= rom_array(20138);
		when "0100111010101011" => data_out <= rom_array(20139);
		when "0100111010101100" => data_out <= rom_array(20140);
		when "0100111010101101" => data_out <= rom_array(20141);
		when "0100111010101110" => data_out <= rom_array(20142);
		when "0100111010101111" => data_out <= rom_array(20143);
		when "0100111010110000" => data_out <= rom_array(20144);
		when "0100111010110001" => data_out <= rom_array(20145);
		when "0100111010110010" => data_out <= rom_array(20146);
		when "0100111010110011" => data_out <= rom_array(20147);
		when "0100111010110100" => data_out <= rom_array(20148);
		when "0100111010110101" => data_out <= rom_array(20149);
		when "0100111010110110" => data_out <= rom_array(20150);
		when "0100111010110111" => data_out <= rom_array(20151);
		when "0100111010111000" => data_out <= rom_array(20152);
		when "0100111010111001" => data_out <= rom_array(20153);
		when "0100111010111010" => data_out <= rom_array(20154);
		when "0100111010111011" => data_out <= rom_array(20155);
		when "0100111010111100" => data_out <= rom_array(20156);
		when "0100111010111101" => data_out <= rom_array(20157);
		when "0100111010111110" => data_out <= rom_array(20158);
		when "0100111010111111" => data_out <= rom_array(20159);
		when "0100111011000000" => data_out <= rom_array(20160);
		when "0100111011000001" => data_out <= rom_array(20161);
		when "0100111011000010" => data_out <= rom_array(20162);
		when "0100111011000011" => data_out <= rom_array(20163);
		when "0100111011000100" => data_out <= rom_array(20164);
		when "0100111011000101" => data_out <= rom_array(20165);
		when "0100111011000110" => data_out <= rom_array(20166);
		when "0100111011000111" => data_out <= rom_array(20167);
		when "0100111011001000" => data_out <= rom_array(20168);
		when "0100111011001001" => data_out <= rom_array(20169);
		when "0100111011001010" => data_out <= rom_array(20170);
		when "0100111011001011" => data_out <= rom_array(20171);
		when "0100111011001100" => data_out <= rom_array(20172);
		when "0100111011001101" => data_out <= rom_array(20173);
		when "0100111011001110" => data_out <= rom_array(20174);
		when "0100111011001111" => data_out <= rom_array(20175);
		when "0100111011010000" => data_out <= rom_array(20176);
		when "0100111011010001" => data_out <= rom_array(20177);
		when "0100111011010010" => data_out <= rom_array(20178);
		when "0100111011010011" => data_out <= rom_array(20179);
		when "0100111011010100" => data_out <= rom_array(20180);
		when "0100111011010101" => data_out <= rom_array(20181);
		when "0100111011010110" => data_out <= rom_array(20182);
		when "0100111011010111" => data_out <= rom_array(20183);
		when "0100111011011000" => data_out <= rom_array(20184);
		when "0100111011011001" => data_out <= rom_array(20185);
		when "0100111011011010" => data_out <= rom_array(20186);
		when "0100111011011011" => data_out <= rom_array(20187);
		when "0100111011011100" => data_out <= rom_array(20188);
		when "0100111011011101" => data_out <= rom_array(20189);
		when "0100111011011110" => data_out <= rom_array(20190);
		when "0100111011011111" => data_out <= rom_array(20191);
		when "0100111011100000" => data_out <= rom_array(20192);
		when "0100111011100001" => data_out <= rom_array(20193);
		when "0100111011100010" => data_out <= rom_array(20194);
		when "0100111011100011" => data_out <= rom_array(20195);
		when "0100111011100100" => data_out <= rom_array(20196);
		when "0100111011100101" => data_out <= rom_array(20197);
		when "0100111011100110" => data_out <= rom_array(20198);
		when "0100111011100111" => data_out <= rom_array(20199);
		when "0100111011101000" => data_out <= rom_array(20200);
		when "0100111011101001" => data_out <= rom_array(20201);
		when "0100111011101010" => data_out <= rom_array(20202);
		when "0100111011101011" => data_out <= rom_array(20203);
		when "0100111011101100" => data_out <= rom_array(20204);
		when "0100111011101101" => data_out <= rom_array(20205);
		when "0100111011101110" => data_out <= rom_array(20206);
		when "0100111011101111" => data_out <= rom_array(20207);
		when "0100111011110000" => data_out <= rom_array(20208);
		when "0100111011110001" => data_out <= rom_array(20209);
		when "0100111011110010" => data_out <= rom_array(20210);
		when "0100111011110011" => data_out <= rom_array(20211);
		when "0100111011110100" => data_out <= rom_array(20212);
		when "0100111011110101" => data_out <= rom_array(20213);
		when "0100111011110110" => data_out <= rom_array(20214);
		when "0100111011110111" => data_out <= rom_array(20215);
		when "0100111011111000" => data_out <= rom_array(20216);
		when "0100111011111001" => data_out <= rom_array(20217);
		when "0100111011111010" => data_out <= rom_array(20218);
		when "0100111011111011" => data_out <= rom_array(20219);
		when "0100111011111100" => data_out <= rom_array(20220);
		when "0100111011111101" => data_out <= rom_array(20221);
		when "0100111011111110" => data_out <= rom_array(20222);
		when "0100111011111111" => data_out <= rom_array(20223);
		when "0100111100000000" => data_out <= rom_array(20224);
		when "0100111100000001" => data_out <= rom_array(20225);
		when "0100111100000010" => data_out <= rom_array(20226);
		when "0100111100000011" => data_out <= rom_array(20227);
		when "0100111100000100" => data_out <= rom_array(20228);
		when "0100111100000101" => data_out <= rom_array(20229);
		when "0100111100000110" => data_out <= rom_array(20230);
		when "0100111100000111" => data_out <= rom_array(20231);
		when "0100111100001000" => data_out <= rom_array(20232);
		when "0100111100001001" => data_out <= rom_array(20233);
		when "0100111100001010" => data_out <= rom_array(20234);
		when "0100111100001011" => data_out <= rom_array(20235);
		when "0100111100001100" => data_out <= rom_array(20236);
		when "0100111100001101" => data_out <= rom_array(20237);
		when "0100111100001110" => data_out <= rom_array(20238);
		when "0100111100001111" => data_out <= rom_array(20239);
		when "0100111100010000" => data_out <= rom_array(20240);
		when "0100111100010001" => data_out <= rom_array(20241);
		when "0100111100010010" => data_out <= rom_array(20242);
		when "0100111100010011" => data_out <= rom_array(20243);
		when "0100111100010100" => data_out <= rom_array(20244);
		when "0100111100010101" => data_out <= rom_array(20245);
		when "0100111100010110" => data_out <= rom_array(20246);
		when "0100111100010111" => data_out <= rom_array(20247);
		when "0100111100011000" => data_out <= rom_array(20248);
		when "0100111100011001" => data_out <= rom_array(20249);
		when "0100111100011010" => data_out <= rom_array(20250);
		when "0100111100011011" => data_out <= rom_array(20251);
		when "0100111100011100" => data_out <= rom_array(20252);
		when "0100111100011101" => data_out <= rom_array(20253);
		when "0100111100011110" => data_out <= rom_array(20254);
		when "0100111100011111" => data_out <= rom_array(20255);
		when "0100111100100000" => data_out <= rom_array(20256);
		when "0100111100100001" => data_out <= rom_array(20257);
		when "0100111100100010" => data_out <= rom_array(20258);
		when "0100111100100011" => data_out <= rom_array(20259);
		when "0100111100100100" => data_out <= rom_array(20260);
		when "0100111100100101" => data_out <= rom_array(20261);
		when "0100111100100110" => data_out <= rom_array(20262);
		when "0100111100100111" => data_out <= rom_array(20263);
		when "0100111100101000" => data_out <= rom_array(20264);
		when "0100111100101001" => data_out <= rom_array(20265);
		when "0100111100101010" => data_out <= rom_array(20266);
		when "0100111100101011" => data_out <= rom_array(20267);
		when "0100111100101100" => data_out <= rom_array(20268);
		when "0100111100101101" => data_out <= rom_array(20269);
		when "0100111100101110" => data_out <= rom_array(20270);
		when "0100111100101111" => data_out <= rom_array(20271);
		when "0100111100110000" => data_out <= rom_array(20272);
		when "0100111100110001" => data_out <= rom_array(20273);
		when "0100111100110010" => data_out <= rom_array(20274);
		when "0100111100110011" => data_out <= rom_array(20275);
		when "0100111100110100" => data_out <= rom_array(20276);
		when "0100111100110101" => data_out <= rom_array(20277);
		when "0100111100110110" => data_out <= rom_array(20278);
		when "0100111100110111" => data_out <= rom_array(20279);
		when "0100111100111000" => data_out <= rom_array(20280);
		when "0100111100111001" => data_out <= rom_array(20281);
		when "0100111100111010" => data_out <= rom_array(20282);
		when "0100111100111011" => data_out <= rom_array(20283);
		when "0100111100111100" => data_out <= rom_array(20284);
		when "0100111100111101" => data_out <= rom_array(20285);
		when "0100111100111110" => data_out <= rom_array(20286);
		when "0100111100111111" => data_out <= rom_array(20287);
		when "0100111101000000" => data_out <= rom_array(20288);
		when "0100111101000001" => data_out <= rom_array(20289);
		when "0100111101000010" => data_out <= rom_array(20290);
		when "0100111101000011" => data_out <= rom_array(20291);
		when "0100111101000100" => data_out <= rom_array(20292);
		when "0100111101000101" => data_out <= rom_array(20293);
		when "0100111101000110" => data_out <= rom_array(20294);
		when "0100111101000111" => data_out <= rom_array(20295);
		when "0100111101001000" => data_out <= rom_array(20296);
		when "0100111101001001" => data_out <= rom_array(20297);
		when "0100111101001010" => data_out <= rom_array(20298);
		when "0100111101001011" => data_out <= rom_array(20299);
		when "0100111101001100" => data_out <= rom_array(20300);
		when "0100111101001101" => data_out <= rom_array(20301);
		when "0100111101001110" => data_out <= rom_array(20302);
		when "0100111101001111" => data_out <= rom_array(20303);
		when "0100111101010000" => data_out <= rom_array(20304);
		when "0100111101010001" => data_out <= rom_array(20305);
		when "0100111101010010" => data_out <= rom_array(20306);
		when "0100111101010011" => data_out <= rom_array(20307);
		when "0100111101010100" => data_out <= rom_array(20308);
		when "0100111101010101" => data_out <= rom_array(20309);
		when "0100111101010110" => data_out <= rom_array(20310);
		when "0100111101010111" => data_out <= rom_array(20311);
		when "0100111101011000" => data_out <= rom_array(20312);
		when "0100111101011001" => data_out <= rom_array(20313);
		when "0100111101011010" => data_out <= rom_array(20314);
		when "0100111101011011" => data_out <= rom_array(20315);
		when "0100111101011100" => data_out <= rom_array(20316);
		when "0100111101011101" => data_out <= rom_array(20317);
		when "0100111101011110" => data_out <= rom_array(20318);
		when "0100111101011111" => data_out <= rom_array(20319);
		when "0100111101100000" => data_out <= rom_array(20320);
		when "0100111101100001" => data_out <= rom_array(20321);
		when "0100111101100010" => data_out <= rom_array(20322);
		when "0100111101100011" => data_out <= rom_array(20323);
		when "0100111101100100" => data_out <= rom_array(20324);
		when "0100111101100101" => data_out <= rom_array(20325);
		when "0100111101100110" => data_out <= rom_array(20326);
		when "0100111101100111" => data_out <= rom_array(20327);
		when "0100111101101000" => data_out <= rom_array(20328);
		when "0100111101101001" => data_out <= rom_array(20329);
		when "0100111101101010" => data_out <= rom_array(20330);
		when "0100111101101011" => data_out <= rom_array(20331);
		when "0100111101101100" => data_out <= rom_array(20332);
		when "0100111101101101" => data_out <= rom_array(20333);
		when "0100111101101110" => data_out <= rom_array(20334);
		when "0100111101101111" => data_out <= rom_array(20335);
		when "0100111101110000" => data_out <= rom_array(20336);
		when "0100111101110001" => data_out <= rom_array(20337);
		when "0100111101110010" => data_out <= rom_array(20338);
		when "0100111101110011" => data_out <= rom_array(20339);
		when "0100111101110100" => data_out <= rom_array(20340);
		when "0100111101110101" => data_out <= rom_array(20341);
		when "0100111101110110" => data_out <= rom_array(20342);
		when "0100111101110111" => data_out <= rom_array(20343);
		when "0100111101111000" => data_out <= rom_array(20344);
		when "0100111101111001" => data_out <= rom_array(20345);
		when "0100111101111010" => data_out <= rom_array(20346);
		when "0100111101111011" => data_out <= rom_array(20347);
		when "0100111101111100" => data_out <= rom_array(20348);
		when "0100111101111101" => data_out <= rom_array(20349);
		when "0100111101111110" => data_out <= rom_array(20350);
		when "0100111101111111" => data_out <= rom_array(20351);
		when "0100111110000000" => data_out <= rom_array(20352);
		when "0100111110000001" => data_out <= rom_array(20353);
		when "0100111110000010" => data_out <= rom_array(20354);
		when "0100111110000011" => data_out <= rom_array(20355);
		when "0100111110000100" => data_out <= rom_array(20356);
		when "0100111110000101" => data_out <= rom_array(20357);
		when "0100111110000110" => data_out <= rom_array(20358);
		when "0100111110000111" => data_out <= rom_array(20359);
		when "0100111110001000" => data_out <= rom_array(20360);
		when "0100111110001001" => data_out <= rom_array(20361);
		when "0100111110001010" => data_out <= rom_array(20362);
		when "0100111110001011" => data_out <= rom_array(20363);
		when "0100111110001100" => data_out <= rom_array(20364);
		when "0100111110001101" => data_out <= rom_array(20365);
		when "0100111110001110" => data_out <= rom_array(20366);
		when "0100111110001111" => data_out <= rom_array(20367);
		when "0100111110010000" => data_out <= rom_array(20368);
		when "0100111110010001" => data_out <= rom_array(20369);
		when "0100111110010010" => data_out <= rom_array(20370);
		when "0100111110010011" => data_out <= rom_array(20371);
		when "0100111110010100" => data_out <= rom_array(20372);
		when "0100111110010101" => data_out <= rom_array(20373);
		when "0100111110010110" => data_out <= rom_array(20374);
		when "0100111110010111" => data_out <= rom_array(20375);
		when "0100111110011000" => data_out <= rom_array(20376);
		when "0100111110011001" => data_out <= rom_array(20377);
		when "0100111110011010" => data_out <= rom_array(20378);
		when "0100111110011011" => data_out <= rom_array(20379);
		when "0100111110011100" => data_out <= rom_array(20380);
		when "0100111110011101" => data_out <= rom_array(20381);
		when "0100111110011110" => data_out <= rom_array(20382);
		when "0100111110011111" => data_out <= rom_array(20383);
		when "0100111110100000" => data_out <= rom_array(20384);
		when "0100111110100001" => data_out <= rom_array(20385);
		when "0100111110100010" => data_out <= rom_array(20386);
		when "0100111110100011" => data_out <= rom_array(20387);
		when "0100111110100100" => data_out <= rom_array(20388);
		when "0100111110100101" => data_out <= rom_array(20389);
		when "0100111110100110" => data_out <= rom_array(20390);
		when "0100111110100111" => data_out <= rom_array(20391);
		when "0100111110101000" => data_out <= rom_array(20392);
		when "0100111110101001" => data_out <= rom_array(20393);
		when "0100111110101010" => data_out <= rom_array(20394);
		when "0100111110101011" => data_out <= rom_array(20395);
		when "0100111110101100" => data_out <= rom_array(20396);
		when "0100111110101101" => data_out <= rom_array(20397);
		when "0100111110101110" => data_out <= rom_array(20398);
		when "0100111110101111" => data_out <= rom_array(20399);
		when "0100111110110000" => data_out <= rom_array(20400);
		when "0100111110110001" => data_out <= rom_array(20401);
		when "0100111110110010" => data_out <= rom_array(20402);
		when "0100111110110011" => data_out <= rom_array(20403);
		when "0100111110110100" => data_out <= rom_array(20404);
		when "0100111110110101" => data_out <= rom_array(20405);
		when "0100111110110110" => data_out <= rom_array(20406);
		when "0100111110110111" => data_out <= rom_array(20407);
		when "0100111110111000" => data_out <= rom_array(20408);
		when "0100111110111001" => data_out <= rom_array(20409);
		when "0100111110111010" => data_out <= rom_array(20410);
		when "0100111110111011" => data_out <= rom_array(20411);
		when "0100111110111100" => data_out <= rom_array(20412);
		when "0100111110111101" => data_out <= rom_array(20413);
		when "0100111110111110" => data_out <= rom_array(20414);
		when "0100111110111111" => data_out <= rom_array(20415);
		when "0100111111000000" => data_out <= rom_array(20416);
		when "0100111111000001" => data_out <= rom_array(20417);
		when "0100111111000010" => data_out <= rom_array(20418);
		when "0100111111000011" => data_out <= rom_array(20419);
		when "0100111111000100" => data_out <= rom_array(20420);
		when "0100111111000101" => data_out <= rom_array(20421);
		when "0100111111000110" => data_out <= rom_array(20422);
		when "0100111111000111" => data_out <= rom_array(20423);
		when "0100111111001000" => data_out <= rom_array(20424);
		when "0100111111001001" => data_out <= rom_array(20425);
		when "0100111111001010" => data_out <= rom_array(20426);
		when "0100111111001011" => data_out <= rom_array(20427);
		when "0100111111001100" => data_out <= rom_array(20428);
		when "0100111111001101" => data_out <= rom_array(20429);
		when "0100111111001110" => data_out <= rom_array(20430);
		when "0100111111001111" => data_out <= rom_array(20431);
		when "0100111111010000" => data_out <= rom_array(20432);
		when "0100111111010001" => data_out <= rom_array(20433);
		when "0100111111010010" => data_out <= rom_array(20434);
		when "0100111111010011" => data_out <= rom_array(20435);
		when "0100111111010100" => data_out <= rom_array(20436);
		when "0100111111010101" => data_out <= rom_array(20437);
		when "0100111111010110" => data_out <= rom_array(20438);
		when "0100111111010111" => data_out <= rom_array(20439);
		when "0100111111011000" => data_out <= rom_array(20440);
		when "0100111111011001" => data_out <= rom_array(20441);
		when "0100111111011010" => data_out <= rom_array(20442);
		when "0100111111011011" => data_out <= rom_array(20443);
		when "0100111111011100" => data_out <= rom_array(20444);
		when "0100111111011101" => data_out <= rom_array(20445);
		when "0100111111011110" => data_out <= rom_array(20446);
		when "0100111111011111" => data_out <= rom_array(20447);
		when "0100111111100000" => data_out <= rom_array(20448);
		when "0100111111100001" => data_out <= rom_array(20449);
		when "0100111111100010" => data_out <= rom_array(20450);
		when "0100111111100011" => data_out <= rom_array(20451);
		when "0100111111100100" => data_out <= rom_array(20452);
		when "0100111111100101" => data_out <= rom_array(20453);
		when "0100111111100110" => data_out <= rom_array(20454);
		when "0100111111100111" => data_out <= rom_array(20455);
		when "0100111111101000" => data_out <= rom_array(20456);
		when "0100111111101001" => data_out <= rom_array(20457);
		when "0100111111101010" => data_out <= rom_array(20458);
		when "0100111111101011" => data_out <= rom_array(20459);
		when "0100111111101100" => data_out <= rom_array(20460);
		when "0100111111101101" => data_out <= rom_array(20461);
		when "0100111111101110" => data_out <= rom_array(20462);
		when "0100111111101111" => data_out <= rom_array(20463);
		when "0100111111110000" => data_out <= rom_array(20464);
		when "0100111111110001" => data_out <= rom_array(20465);
		when "0100111111110010" => data_out <= rom_array(20466);
		when "0100111111110011" => data_out <= rom_array(20467);
		when "0100111111110100" => data_out <= rom_array(20468);
		when "0100111111110101" => data_out <= rom_array(20469);
		when "0100111111110110" => data_out <= rom_array(20470);
		when "0100111111110111" => data_out <= rom_array(20471);
		when "0100111111111000" => data_out <= rom_array(20472);
		when "0100111111111001" => data_out <= rom_array(20473);
		when "0100111111111010" => data_out <= rom_array(20474);
		when "0100111111111011" => data_out <= rom_array(20475);
		when "0100111111111100" => data_out <= rom_array(20476);
		when "0100111111111101" => data_out <= rom_array(20477);
		when "0100111111111110" => data_out <= rom_array(20478);
		when "0100111111111111" => data_out <= rom_array(20479);
		when "0101000000000000" => data_out <= rom_array(20480);
		when "0101000000000001" => data_out <= rom_array(20481);
		when "0101000000000010" => data_out <= rom_array(20482);
		when "0101000000000011" => data_out <= rom_array(20483);
		when "0101000000000100" => data_out <= rom_array(20484);
		when "0101000000000101" => data_out <= rom_array(20485);
		when "0101000000000110" => data_out <= rom_array(20486);
		when "0101000000000111" => data_out <= rom_array(20487);
		when "0101000000001000" => data_out <= rom_array(20488);
		when "0101000000001001" => data_out <= rom_array(20489);
		when "0101000000001010" => data_out <= rom_array(20490);
		when "0101000000001011" => data_out <= rom_array(20491);
		when "0101000000001100" => data_out <= rom_array(20492);
		when "0101000000001101" => data_out <= rom_array(20493);
		when "0101000000001110" => data_out <= rom_array(20494);
		when "0101000000001111" => data_out <= rom_array(20495);
		when "0101000000010000" => data_out <= rom_array(20496);
		when "0101000000010001" => data_out <= rom_array(20497);
		when "0101000000010010" => data_out <= rom_array(20498);
		when "0101000000010011" => data_out <= rom_array(20499);
		when "0101000000010100" => data_out <= rom_array(20500);
		when "0101000000010101" => data_out <= rom_array(20501);
		when "0101000000010110" => data_out <= rom_array(20502);
		when "0101000000010111" => data_out <= rom_array(20503);
		when "0101000000011000" => data_out <= rom_array(20504);
		when "0101000000011001" => data_out <= rom_array(20505);
		when "0101000000011010" => data_out <= rom_array(20506);
		when "0101000000011011" => data_out <= rom_array(20507);
		when "0101000000011100" => data_out <= rom_array(20508);
		when "0101000000011101" => data_out <= rom_array(20509);
		when "0101000000011110" => data_out <= rom_array(20510);
		when "0101000000011111" => data_out <= rom_array(20511);
		when "0101000000100000" => data_out <= rom_array(20512);
		when "0101000000100001" => data_out <= rom_array(20513);
		when "0101000000100010" => data_out <= rom_array(20514);
		when "0101000000100011" => data_out <= rom_array(20515);
		when "0101000000100100" => data_out <= rom_array(20516);
		when "0101000000100101" => data_out <= rom_array(20517);
		when "0101000000100110" => data_out <= rom_array(20518);
		when "0101000000100111" => data_out <= rom_array(20519);
		when "0101000000101000" => data_out <= rom_array(20520);
		when "0101000000101001" => data_out <= rom_array(20521);
		when "0101000000101010" => data_out <= rom_array(20522);
		when "0101000000101011" => data_out <= rom_array(20523);
		when "0101000000101100" => data_out <= rom_array(20524);
		when "0101000000101101" => data_out <= rom_array(20525);
		when "0101000000101110" => data_out <= rom_array(20526);
		when "0101000000101111" => data_out <= rom_array(20527);
		when "0101000000110000" => data_out <= rom_array(20528);
		when "0101000000110001" => data_out <= rom_array(20529);
		when "0101000000110010" => data_out <= rom_array(20530);
		when "0101000000110011" => data_out <= rom_array(20531);
		when "0101000000110100" => data_out <= rom_array(20532);
		when "0101000000110101" => data_out <= rom_array(20533);
		when "0101000000110110" => data_out <= rom_array(20534);
		when "0101000000110111" => data_out <= rom_array(20535);
		when "0101000000111000" => data_out <= rom_array(20536);
		when "0101000000111001" => data_out <= rom_array(20537);
		when "0101000000111010" => data_out <= rom_array(20538);
		when "0101000000111011" => data_out <= rom_array(20539);
		when "0101000000111100" => data_out <= rom_array(20540);
		when "0101000000111101" => data_out <= rom_array(20541);
		when "0101000000111110" => data_out <= rom_array(20542);
		when "0101000000111111" => data_out <= rom_array(20543);
		when "0101000001000000" => data_out <= rom_array(20544);
		when "0101000001000001" => data_out <= rom_array(20545);
		when "0101000001000010" => data_out <= rom_array(20546);
		when "0101000001000011" => data_out <= rom_array(20547);
		when "0101000001000100" => data_out <= rom_array(20548);
		when "0101000001000101" => data_out <= rom_array(20549);
		when "0101000001000110" => data_out <= rom_array(20550);
		when "0101000001000111" => data_out <= rom_array(20551);
		when "0101000001001000" => data_out <= rom_array(20552);
		when "0101000001001001" => data_out <= rom_array(20553);
		when "0101000001001010" => data_out <= rom_array(20554);
		when "0101000001001011" => data_out <= rom_array(20555);
		when "0101000001001100" => data_out <= rom_array(20556);
		when "0101000001001101" => data_out <= rom_array(20557);
		when "0101000001001110" => data_out <= rom_array(20558);
		when "0101000001001111" => data_out <= rom_array(20559);
		when "0101000001010000" => data_out <= rom_array(20560);
		when "0101000001010001" => data_out <= rom_array(20561);
		when "0101000001010010" => data_out <= rom_array(20562);
		when "0101000001010011" => data_out <= rom_array(20563);
		when "0101000001010100" => data_out <= rom_array(20564);
		when "0101000001010101" => data_out <= rom_array(20565);
		when "0101000001010110" => data_out <= rom_array(20566);
		when "0101000001010111" => data_out <= rom_array(20567);
		when "0101000001011000" => data_out <= rom_array(20568);
		when "0101000001011001" => data_out <= rom_array(20569);
		when "0101000001011010" => data_out <= rom_array(20570);
		when "0101000001011011" => data_out <= rom_array(20571);
		when "0101000001011100" => data_out <= rom_array(20572);
		when "0101000001011101" => data_out <= rom_array(20573);
		when "0101000001011110" => data_out <= rom_array(20574);
		when "0101000001011111" => data_out <= rom_array(20575);
		when "0101000001100000" => data_out <= rom_array(20576);
		when "0101000001100001" => data_out <= rom_array(20577);
		when "0101000001100010" => data_out <= rom_array(20578);
		when "0101000001100011" => data_out <= rom_array(20579);
		when "0101000001100100" => data_out <= rom_array(20580);
		when "0101000001100101" => data_out <= rom_array(20581);
		when "0101000001100110" => data_out <= rom_array(20582);
		when "0101000001100111" => data_out <= rom_array(20583);
		when "0101000001101000" => data_out <= rom_array(20584);
		when "0101000001101001" => data_out <= rom_array(20585);
		when "0101000001101010" => data_out <= rom_array(20586);
		when "0101000001101011" => data_out <= rom_array(20587);
		when "0101000001101100" => data_out <= rom_array(20588);
		when "0101000001101101" => data_out <= rom_array(20589);
		when "0101000001101110" => data_out <= rom_array(20590);
		when "0101000001101111" => data_out <= rom_array(20591);
		when "0101000001110000" => data_out <= rom_array(20592);
		when "0101000001110001" => data_out <= rom_array(20593);
		when "0101000001110010" => data_out <= rom_array(20594);
		when "0101000001110011" => data_out <= rom_array(20595);
		when "0101000001110100" => data_out <= rom_array(20596);
		when "0101000001110101" => data_out <= rom_array(20597);
		when "0101000001110110" => data_out <= rom_array(20598);
		when "0101000001110111" => data_out <= rom_array(20599);
		when "0101000001111000" => data_out <= rom_array(20600);
		when "0101000001111001" => data_out <= rom_array(20601);
		when "0101000001111010" => data_out <= rom_array(20602);
		when "0101000001111011" => data_out <= rom_array(20603);
		when "0101000001111100" => data_out <= rom_array(20604);
		when "0101000001111101" => data_out <= rom_array(20605);
		when "0101000001111110" => data_out <= rom_array(20606);
		when "0101000001111111" => data_out <= rom_array(20607);
		when "0101000010000000" => data_out <= rom_array(20608);
		when "0101000010000001" => data_out <= rom_array(20609);
		when "0101000010000010" => data_out <= rom_array(20610);
		when "0101000010000011" => data_out <= rom_array(20611);
		when "0101000010000100" => data_out <= rom_array(20612);
		when "0101000010000101" => data_out <= rom_array(20613);
		when "0101000010000110" => data_out <= rom_array(20614);
		when "0101000010000111" => data_out <= rom_array(20615);
		when "0101000010001000" => data_out <= rom_array(20616);
		when "0101000010001001" => data_out <= rom_array(20617);
		when "0101000010001010" => data_out <= rom_array(20618);
		when "0101000010001011" => data_out <= rom_array(20619);
		when "0101000010001100" => data_out <= rom_array(20620);
		when "0101000010001101" => data_out <= rom_array(20621);
		when "0101000010001110" => data_out <= rom_array(20622);
		when "0101000010001111" => data_out <= rom_array(20623);
		when "0101000010010000" => data_out <= rom_array(20624);
		when "0101000010010001" => data_out <= rom_array(20625);
		when "0101000010010010" => data_out <= rom_array(20626);
		when "0101000010010011" => data_out <= rom_array(20627);
		when "0101000010010100" => data_out <= rom_array(20628);
		when "0101000010010101" => data_out <= rom_array(20629);
		when "0101000010010110" => data_out <= rom_array(20630);
		when "0101000010010111" => data_out <= rom_array(20631);
		when "0101000010011000" => data_out <= rom_array(20632);
		when "0101000010011001" => data_out <= rom_array(20633);
		when "0101000010011010" => data_out <= rom_array(20634);
		when "0101000010011011" => data_out <= rom_array(20635);
		when "0101000010011100" => data_out <= rom_array(20636);
		when "0101000010011101" => data_out <= rom_array(20637);
		when "0101000010011110" => data_out <= rom_array(20638);
		when "0101000010011111" => data_out <= rom_array(20639);
		when "0101000010100000" => data_out <= rom_array(20640);
		when "0101000010100001" => data_out <= rom_array(20641);
		when "0101000010100010" => data_out <= rom_array(20642);
		when "0101000010100011" => data_out <= rom_array(20643);
		when "0101000010100100" => data_out <= rom_array(20644);
		when "0101000010100101" => data_out <= rom_array(20645);
		when "0101000010100110" => data_out <= rom_array(20646);
		when "0101000010100111" => data_out <= rom_array(20647);
		when "0101000010101000" => data_out <= rom_array(20648);
		when "0101000010101001" => data_out <= rom_array(20649);
		when "0101000010101010" => data_out <= rom_array(20650);
		when "0101000010101011" => data_out <= rom_array(20651);
		when "0101000010101100" => data_out <= rom_array(20652);
		when "0101000010101101" => data_out <= rom_array(20653);
		when "0101000010101110" => data_out <= rom_array(20654);
		when "0101000010101111" => data_out <= rom_array(20655);
		when "0101000010110000" => data_out <= rom_array(20656);
		when "0101000010110001" => data_out <= rom_array(20657);
		when "0101000010110010" => data_out <= rom_array(20658);
		when "0101000010110011" => data_out <= rom_array(20659);
		when "0101000010110100" => data_out <= rom_array(20660);
		when "0101000010110101" => data_out <= rom_array(20661);
		when "0101000010110110" => data_out <= rom_array(20662);
		when "0101000010110111" => data_out <= rom_array(20663);
		when "0101000010111000" => data_out <= rom_array(20664);
		when "0101000010111001" => data_out <= rom_array(20665);
		when "0101000010111010" => data_out <= rom_array(20666);
		when "0101000010111011" => data_out <= rom_array(20667);
		when "0101000010111100" => data_out <= rom_array(20668);
		when "0101000010111101" => data_out <= rom_array(20669);
		when "0101000010111110" => data_out <= rom_array(20670);
		when "0101000010111111" => data_out <= rom_array(20671);
		when "0101000011000000" => data_out <= rom_array(20672);
		when "0101000011000001" => data_out <= rom_array(20673);
		when "0101000011000010" => data_out <= rom_array(20674);
		when "0101000011000011" => data_out <= rom_array(20675);
		when "0101000011000100" => data_out <= rom_array(20676);
		when "0101000011000101" => data_out <= rom_array(20677);
		when "0101000011000110" => data_out <= rom_array(20678);
		when "0101000011000111" => data_out <= rom_array(20679);
		when "0101000011001000" => data_out <= rom_array(20680);
		when "0101000011001001" => data_out <= rom_array(20681);
		when "0101000011001010" => data_out <= rom_array(20682);
		when "0101000011001011" => data_out <= rom_array(20683);
		when "0101000011001100" => data_out <= rom_array(20684);
		when "0101000011001101" => data_out <= rom_array(20685);
		when "0101000011001110" => data_out <= rom_array(20686);
		when "0101000011001111" => data_out <= rom_array(20687);
		when "0101000011010000" => data_out <= rom_array(20688);
		when "0101000011010001" => data_out <= rom_array(20689);
		when "0101000011010010" => data_out <= rom_array(20690);
		when "0101000011010011" => data_out <= rom_array(20691);
		when "0101000011010100" => data_out <= rom_array(20692);
		when "0101000011010101" => data_out <= rom_array(20693);
		when "0101000011010110" => data_out <= rom_array(20694);
		when "0101000011010111" => data_out <= rom_array(20695);
		when "0101000011011000" => data_out <= rom_array(20696);
		when "0101000011011001" => data_out <= rom_array(20697);
		when "0101000011011010" => data_out <= rom_array(20698);
		when "0101000011011011" => data_out <= rom_array(20699);
		when "0101000011011100" => data_out <= rom_array(20700);
		when "0101000011011101" => data_out <= rom_array(20701);
		when "0101000011011110" => data_out <= rom_array(20702);
		when "0101000011011111" => data_out <= rom_array(20703);
		when "0101000011100000" => data_out <= rom_array(20704);
		when "0101000011100001" => data_out <= rom_array(20705);
		when "0101000011100010" => data_out <= rom_array(20706);
		when "0101000011100011" => data_out <= rom_array(20707);
		when "0101000011100100" => data_out <= rom_array(20708);
		when "0101000011100101" => data_out <= rom_array(20709);
		when "0101000011100110" => data_out <= rom_array(20710);
		when "0101000011100111" => data_out <= rom_array(20711);
		when "0101000011101000" => data_out <= rom_array(20712);
		when "0101000011101001" => data_out <= rom_array(20713);
		when "0101000011101010" => data_out <= rom_array(20714);
		when "0101000011101011" => data_out <= rom_array(20715);
		when "0101000011101100" => data_out <= rom_array(20716);
		when "0101000011101101" => data_out <= rom_array(20717);
		when "0101000011101110" => data_out <= rom_array(20718);
		when "0101000011101111" => data_out <= rom_array(20719);
		when "0101000011110000" => data_out <= rom_array(20720);
		when "0101000011110001" => data_out <= rom_array(20721);
		when "0101000011110010" => data_out <= rom_array(20722);
		when "0101000011110011" => data_out <= rom_array(20723);
		when "0101000011110100" => data_out <= rom_array(20724);
		when "0101000011110101" => data_out <= rom_array(20725);
		when "0101000011110110" => data_out <= rom_array(20726);
		when "0101000011110111" => data_out <= rom_array(20727);
		when "0101000011111000" => data_out <= rom_array(20728);
		when "0101000011111001" => data_out <= rom_array(20729);
		when "0101000011111010" => data_out <= rom_array(20730);
		when "0101000011111011" => data_out <= rom_array(20731);
		when "0101000011111100" => data_out <= rom_array(20732);
		when "0101000011111101" => data_out <= rom_array(20733);
		when "0101000011111110" => data_out <= rom_array(20734);
		when "0101000011111111" => data_out <= rom_array(20735);
		when "0101000100000000" => data_out <= rom_array(20736);
		when "0101000100000001" => data_out <= rom_array(20737);
		when "0101000100000010" => data_out <= rom_array(20738);
		when "0101000100000011" => data_out <= rom_array(20739);
		when "0101000100000100" => data_out <= rom_array(20740);
		when "0101000100000101" => data_out <= rom_array(20741);
		when "0101000100000110" => data_out <= rom_array(20742);
		when "0101000100000111" => data_out <= rom_array(20743);
		when "0101000100001000" => data_out <= rom_array(20744);
		when "0101000100001001" => data_out <= rom_array(20745);
		when "0101000100001010" => data_out <= rom_array(20746);
		when "0101000100001011" => data_out <= rom_array(20747);
		when "0101000100001100" => data_out <= rom_array(20748);
		when "0101000100001101" => data_out <= rom_array(20749);
		when "0101000100001110" => data_out <= rom_array(20750);
		when "0101000100001111" => data_out <= rom_array(20751);
		when "0101000100010000" => data_out <= rom_array(20752);
		when "0101000100010001" => data_out <= rom_array(20753);
		when "0101000100010010" => data_out <= rom_array(20754);
		when "0101000100010011" => data_out <= rom_array(20755);
		when "0101000100010100" => data_out <= rom_array(20756);
		when "0101000100010101" => data_out <= rom_array(20757);
		when "0101000100010110" => data_out <= rom_array(20758);
		when "0101000100010111" => data_out <= rom_array(20759);
		when "0101000100011000" => data_out <= rom_array(20760);
		when "0101000100011001" => data_out <= rom_array(20761);
		when "0101000100011010" => data_out <= rom_array(20762);
		when "0101000100011011" => data_out <= rom_array(20763);
		when "0101000100011100" => data_out <= rom_array(20764);
		when "0101000100011101" => data_out <= rom_array(20765);
		when "0101000100011110" => data_out <= rom_array(20766);
		when "0101000100011111" => data_out <= rom_array(20767);
		when "0101000100100000" => data_out <= rom_array(20768);
		when "0101000100100001" => data_out <= rom_array(20769);
		when "0101000100100010" => data_out <= rom_array(20770);
		when "0101000100100011" => data_out <= rom_array(20771);
		when "0101000100100100" => data_out <= rom_array(20772);
		when "0101000100100101" => data_out <= rom_array(20773);
		when "0101000100100110" => data_out <= rom_array(20774);
		when "0101000100100111" => data_out <= rom_array(20775);
		when "0101000100101000" => data_out <= rom_array(20776);
		when "0101000100101001" => data_out <= rom_array(20777);
		when "0101000100101010" => data_out <= rom_array(20778);
		when "0101000100101011" => data_out <= rom_array(20779);
		when "0101000100101100" => data_out <= rom_array(20780);
		when "0101000100101101" => data_out <= rom_array(20781);
		when "0101000100101110" => data_out <= rom_array(20782);
		when "0101000100101111" => data_out <= rom_array(20783);
		when "0101000100110000" => data_out <= rom_array(20784);
		when "0101000100110001" => data_out <= rom_array(20785);
		when "0101000100110010" => data_out <= rom_array(20786);
		when "0101000100110011" => data_out <= rom_array(20787);
		when "0101000100110100" => data_out <= rom_array(20788);
		when "0101000100110101" => data_out <= rom_array(20789);
		when "0101000100110110" => data_out <= rom_array(20790);
		when "0101000100110111" => data_out <= rom_array(20791);
		when "0101000100111000" => data_out <= rom_array(20792);
		when "0101000100111001" => data_out <= rom_array(20793);
		when "0101000100111010" => data_out <= rom_array(20794);
		when "0101000100111011" => data_out <= rom_array(20795);
		when "0101000100111100" => data_out <= rom_array(20796);
		when "0101000100111101" => data_out <= rom_array(20797);
		when "0101000100111110" => data_out <= rom_array(20798);
		when "0101000100111111" => data_out <= rom_array(20799);
		when "0101000101000000" => data_out <= rom_array(20800);
		when "0101000101000001" => data_out <= rom_array(20801);
		when "0101000101000010" => data_out <= rom_array(20802);
		when "0101000101000011" => data_out <= rom_array(20803);
		when "0101000101000100" => data_out <= rom_array(20804);
		when "0101000101000101" => data_out <= rom_array(20805);
		when "0101000101000110" => data_out <= rom_array(20806);
		when "0101000101000111" => data_out <= rom_array(20807);
		when "0101000101001000" => data_out <= rom_array(20808);
		when "0101000101001001" => data_out <= rom_array(20809);
		when "0101000101001010" => data_out <= rom_array(20810);
		when "0101000101001011" => data_out <= rom_array(20811);
		when "0101000101001100" => data_out <= rom_array(20812);
		when "0101000101001101" => data_out <= rom_array(20813);
		when "0101000101001110" => data_out <= rom_array(20814);
		when "0101000101001111" => data_out <= rom_array(20815);
		when "0101000101010000" => data_out <= rom_array(20816);
		when "0101000101010001" => data_out <= rom_array(20817);
		when "0101000101010010" => data_out <= rom_array(20818);
		when "0101000101010011" => data_out <= rom_array(20819);
		when "0101000101010100" => data_out <= rom_array(20820);
		when "0101000101010101" => data_out <= rom_array(20821);
		when "0101000101010110" => data_out <= rom_array(20822);
		when "0101000101010111" => data_out <= rom_array(20823);
		when "0101000101011000" => data_out <= rom_array(20824);
		when "0101000101011001" => data_out <= rom_array(20825);
		when "0101000101011010" => data_out <= rom_array(20826);
		when "0101000101011011" => data_out <= rom_array(20827);
		when "0101000101011100" => data_out <= rom_array(20828);
		when "0101000101011101" => data_out <= rom_array(20829);
		when "0101000101011110" => data_out <= rom_array(20830);
		when "0101000101011111" => data_out <= rom_array(20831);
		when "0101000101100000" => data_out <= rom_array(20832);
		when "0101000101100001" => data_out <= rom_array(20833);
		when "0101000101100010" => data_out <= rom_array(20834);
		when "0101000101100011" => data_out <= rom_array(20835);
		when "0101000101100100" => data_out <= rom_array(20836);
		when "0101000101100101" => data_out <= rom_array(20837);
		when "0101000101100110" => data_out <= rom_array(20838);
		when "0101000101100111" => data_out <= rom_array(20839);
		when "0101000101101000" => data_out <= rom_array(20840);
		when "0101000101101001" => data_out <= rom_array(20841);
		when "0101000101101010" => data_out <= rom_array(20842);
		when "0101000101101011" => data_out <= rom_array(20843);
		when "0101000101101100" => data_out <= rom_array(20844);
		when "0101000101101101" => data_out <= rom_array(20845);
		when "0101000101101110" => data_out <= rom_array(20846);
		when "0101000101101111" => data_out <= rom_array(20847);
		when "0101000101110000" => data_out <= rom_array(20848);
		when "0101000101110001" => data_out <= rom_array(20849);
		when "0101000101110010" => data_out <= rom_array(20850);
		when "0101000101110011" => data_out <= rom_array(20851);
		when "0101000101110100" => data_out <= rom_array(20852);
		when "0101000101110101" => data_out <= rom_array(20853);
		when "0101000101110110" => data_out <= rom_array(20854);
		when "0101000101110111" => data_out <= rom_array(20855);
		when "0101000101111000" => data_out <= rom_array(20856);
		when "0101000101111001" => data_out <= rom_array(20857);
		when "0101000101111010" => data_out <= rom_array(20858);
		when "0101000101111011" => data_out <= rom_array(20859);
		when "0101000101111100" => data_out <= rom_array(20860);
		when "0101000101111101" => data_out <= rom_array(20861);
		when "0101000101111110" => data_out <= rom_array(20862);
		when "0101000101111111" => data_out <= rom_array(20863);
		when "0101000110000000" => data_out <= rom_array(20864);
		when "0101000110000001" => data_out <= rom_array(20865);
		when "0101000110000010" => data_out <= rom_array(20866);
		when "0101000110000011" => data_out <= rom_array(20867);
		when "0101000110000100" => data_out <= rom_array(20868);
		when "0101000110000101" => data_out <= rom_array(20869);
		when "0101000110000110" => data_out <= rom_array(20870);
		when "0101000110000111" => data_out <= rom_array(20871);
		when "0101000110001000" => data_out <= rom_array(20872);
		when "0101000110001001" => data_out <= rom_array(20873);
		when "0101000110001010" => data_out <= rom_array(20874);
		when "0101000110001011" => data_out <= rom_array(20875);
		when "0101000110001100" => data_out <= rom_array(20876);
		when "0101000110001101" => data_out <= rom_array(20877);
		when "0101000110001110" => data_out <= rom_array(20878);
		when "0101000110001111" => data_out <= rom_array(20879);
		when "0101000110010000" => data_out <= rom_array(20880);
		when "0101000110010001" => data_out <= rom_array(20881);
		when "0101000110010010" => data_out <= rom_array(20882);
		when "0101000110010011" => data_out <= rom_array(20883);
		when "0101000110010100" => data_out <= rom_array(20884);
		when "0101000110010101" => data_out <= rom_array(20885);
		when "0101000110010110" => data_out <= rom_array(20886);
		when "0101000110010111" => data_out <= rom_array(20887);
		when "0101000110011000" => data_out <= rom_array(20888);
		when "0101000110011001" => data_out <= rom_array(20889);
		when "0101000110011010" => data_out <= rom_array(20890);
		when "0101000110011011" => data_out <= rom_array(20891);
		when "0101000110011100" => data_out <= rom_array(20892);
		when "0101000110011101" => data_out <= rom_array(20893);
		when "0101000110011110" => data_out <= rom_array(20894);
		when "0101000110011111" => data_out <= rom_array(20895);
		when "0101000110100000" => data_out <= rom_array(20896);
		when "0101000110100001" => data_out <= rom_array(20897);
		when "0101000110100010" => data_out <= rom_array(20898);
		when "0101000110100011" => data_out <= rom_array(20899);
		when "0101000110100100" => data_out <= rom_array(20900);
		when "0101000110100101" => data_out <= rom_array(20901);
		when "0101000110100110" => data_out <= rom_array(20902);
		when "0101000110100111" => data_out <= rom_array(20903);
		when "0101000110101000" => data_out <= rom_array(20904);
		when "0101000110101001" => data_out <= rom_array(20905);
		when "0101000110101010" => data_out <= rom_array(20906);
		when "0101000110101011" => data_out <= rom_array(20907);
		when "0101000110101100" => data_out <= rom_array(20908);
		when "0101000110101101" => data_out <= rom_array(20909);
		when "0101000110101110" => data_out <= rom_array(20910);
		when "0101000110101111" => data_out <= rom_array(20911);
		when "0101000110110000" => data_out <= rom_array(20912);
		when "0101000110110001" => data_out <= rom_array(20913);
		when "0101000110110010" => data_out <= rom_array(20914);
		when "0101000110110011" => data_out <= rom_array(20915);
		when "0101000110110100" => data_out <= rom_array(20916);
		when "0101000110110101" => data_out <= rom_array(20917);
		when "0101000110110110" => data_out <= rom_array(20918);
		when "0101000110110111" => data_out <= rom_array(20919);
		when "0101000110111000" => data_out <= rom_array(20920);
		when "0101000110111001" => data_out <= rom_array(20921);
		when "0101000110111010" => data_out <= rom_array(20922);
		when "0101000110111011" => data_out <= rom_array(20923);
		when "0101000110111100" => data_out <= rom_array(20924);
		when "0101000110111101" => data_out <= rom_array(20925);
		when "0101000110111110" => data_out <= rom_array(20926);
		when "0101000110111111" => data_out <= rom_array(20927);
		when "0101000111000000" => data_out <= rom_array(20928);
		when "0101000111000001" => data_out <= rom_array(20929);
		when "0101000111000010" => data_out <= rom_array(20930);
		when "0101000111000011" => data_out <= rom_array(20931);
		when "0101000111000100" => data_out <= rom_array(20932);
		when "0101000111000101" => data_out <= rom_array(20933);
		when "0101000111000110" => data_out <= rom_array(20934);
		when "0101000111000111" => data_out <= rom_array(20935);
		when "0101000111001000" => data_out <= rom_array(20936);
		when "0101000111001001" => data_out <= rom_array(20937);
		when "0101000111001010" => data_out <= rom_array(20938);
		when "0101000111001011" => data_out <= rom_array(20939);
		when "0101000111001100" => data_out <= rom_array(20940);
		when "0101000111001101" => data_out <= rom_array(20941);
		when "0101000111001110" => data_out <= rom_array(20942);
		when "0101000111001111" => data_out <= rom_array(20943);
		when "0101000111010000" => data_out <= rom_array(20944);
		when "0101000111010001" => data_out <= rom_array(20945);
		when "0101000111010010" => data_out <= rom_array(20946);
		when "0101000111010011" => data_out <= rom_array(20947);
		when "0101000111010100" => data_out <= rom_array(20948);
		when "0101000111010101" => data_out <= rom_array(20949);
		when "0101000111010110" => data_out <= rom_array(20950);
		when "0101000111010111" => data_out <= rom_array(20951);
		when "0101000111011000" => data_out <= rom_array(20952);
		when "0101000111011001" => data_out <= rom_array(20953);
		when "0101000111011010" => data_out <= rom_array(20954);
		when "0101000111011011" => data_out <= rom_array(20955);
		when "0101000111011100" => data_out <= rom_array(20956);
		when "0101000111011101" => data_out <= rom_array(20957);
		when "0101000111011110" => data_out <= rom_array(20958);
		when "0101000111011111" => data_out <= rom_array(20959);
		when "0101000111100000" => data_out <= rom_array(20960);
		when "0101000111100001" => data_out <= rom_array(20961);
		when "0101000111100010" => data_out <= rom_array(20962);
		when "0101000111100011" => data_out <= rom_array(20963);
		when "0101000111100100" => data_out <= rom_array(20964);
		when "0101000111100101" => data_out <= rom_array(20965);
		when "0101000111100110" => data_out <= rom_array(20966);
		when "0101000111100111" => data_out <= rom_array(20967);
		when "0101000111101000" => data_out <= rom_array(20968);
		when "0101000111101001" => data_out <= rom_array(20969);
		when "0101000111101010" => data_out <= rom_array(20970);
		when "0101000111101011" => data_out <= rom_array(20971);
		when "0101000111101100" => data_out <= rom_array(20972);
		when "0101000111101101" => data_out <= rom_array(20973);
		when "0101000111101110" => data_out <= rom_array(20974);
		when "0101000111101111" => data_out <= rom_array(20975);
		when "0101000111110000" => data_out <= rom_array(20976);
		when "0101000111110001" => data_out <= rom_array(20977);
		when "0101000111110010" => data_out <= rom_array(20978);
		when "0101000111110011" => data_out <= rom_array(20979);
		when "0101000111110100" => data_out <= rom_array(20980);
		when "0101000111110101" => data_out <= rom_array(20981);
		when "0101000111110110" => data_out <= rom_array(20982);
		when "0101000111110111" => data_out <= rom_array(20983);
		when "0101000111111000" => data_out <= rom_array(20984);
		when "0101000111111001" => data_out <= rom_array(20985);
		when "0101000111111010" => data_out <= rom_array(20986);
		when "0101000111111011" => data_out <= rom_array(20987);
		when "0101000111111100" => data_out <= rom_array(20988);
		when "0101000111111101" => data_out <= rom_array(20989);
		when "0101000111111110" => data_out <= rom_array(20990);
		when "0101000111111111" => data_out <= rom_array(20991);
		when "0101001000000000" => data_out <= rom_array(20992);
		when "0101001000000001" => data_out <= rom_array(20993);
		when "0101001000000010" => data_out <= rom_array(20994);
		when "0101001000000011" => data_out <= rom_array(20995);
		when "0101001000000100" => data_out <= rom_array(20996);
		when "0101001000000101" => data_out <= rom_array(20997);
		when "0101001000000110" => data_out <= rom_array(20998);
		when "0101001000000111" => data_out <= rom_array(20999);
		when "0101001000001000" => data_out <= rom_array(21000);
		when "0101001000001001" => data_out <= rom_array(21001);
		when "0101001000001010" => data_out <= rom_array(21002);
		when "0101001000001011" => data_out <= rom_array(21003);
		when "0101001000001100" => data_out <= rom_array(21004);
		when "0101001000001101" => data_out <= rom_array(21005);
		when "0101001000001110" => data_out <= rom_array(21006);
		when "0101001000001111" => data_out <= rom_array(21007);
		when "0101001000010000" => data_out <= rom_array(21008);
		when "0101001000010001" => data_out <= rom_array(21009);
		when "0101001000010010" => data_out <= rom_array(21010);
		when "0101001000010011" => data_out <= rom_array(21011);
		when "0101001000010100" => data_out <= rom_array(21012);
		when "0101001000010101" => data_out <= rom_array(21013);
		when "0101001000010110" => data_out <= rom_array(21014);
		when "0101001000010111" => data_out <= rom_array(21015);
		when "0101001000011000" => data_out <= rom_array(21016);
		when "0101001000011001" => data_out <= rom_array(21017);
		when "0101001000011010" => data_out <= rom_array(21018);
		when "0101001000011011" => data_out <= rom_array(21019);
		when "0101001000011100" => data_out <= rom_array(21020);
		when "0101001000011101" => data_out <= rom_array(21021);
		when "0101001000011110" => data_out <= rom_array(21022);
		when "0101001000011111" => data_out <= rom_array(21023);
		when "0101001000100000" => data_out <= rom_array(21024);
		when "0101001000100001" => data_out <= rom_array(21025);
		when "0101001000100010" => data_out <= rom_array(21026);
		when "0101001000100011" => data_out <= rom_array(21027);
		when "0101001000100100" => data_out <= rom_array(21028);
		when "0101001000100101" => data_out <= rom_array(21029);
		when "0101001000100110" => data_out <= rom_array(21030);
		when "0101001000100111" => data_out <= rom_array(21031);
		when "0101001000101000" => data_out <= rom_array(21032);
		when "0101001000101001" => data_out <= rom_array(21033);
		when "0101001000101010" => data_out <= rom_array(21034);
		when "0101001000101011" => data_out <= rom_array(21035);
		when "0101001000101100" => data_out <= rom_array(21036);
		when "0101001000101101" => data_out <= rom_array(21037);
		when "0101001000101110" => data_out <= rom_array(21038);
		when "0101001000101111" => data_out <= rom_array(21039);
		when "0101001000110000" => data_out <= rom_array(21040);
		when "0101001000110001" => data_out <= rom_array(21041);
		when "0101001000110010" => data_out <= rom_array(21042);
		when "0101001000110011" => data_out <= rom_array(21043);
		when "0101001000110100" => data_out <= rom_array(21044);
		when "0101001000110101" => data_out <= rom_array(21045);
		when "0101001000110110" => data_out <= rom_array(21046);
		when "0101001000110111" => data_out <= rom_array(21047);
		when "0101001000111000" => data_out <= rom_array(21048);
		when "0101001000111001" => data_out <= rom_array(21049);
		when "0101001000111010" => data_out <= rom_array(21050);
		when "0101001000111011" => data_out <= rom_array(21051);
		when "0101001000111100" => data_out <= rom_array(21052);
		when "0101001000111101" => data_out <= rom_array(21053);
		when "0101001000111110" => data_out <= rom_array(21054);
		when "0101001000111111" => data_out <= rom_array(21055);
		when "0101001001000000" => data_out <= rom_array(21056);
		when "0101001001000001" => data_out <= rom_array(21057);
		when "0101001001000010" => data_out <= rom_array(21058);
		when "0101001001000011" => data_out <= rom_array(21059);
		when "0101001001000100" => data_out <= rom_array(21060);
		when "0101001001000101" => data_out <= rom_array(21061);
		when "0101001001000110" => data_out <= rom_array(21062);
		when "0101001001000111" => data_out <= rom_array(21063);
		when "0101001001001000" => data_out <= rom_array(21064);
		when "0101001001001001" => data_out <= rom_array(21065);
		when "0101001001001010" => data_out <= rom_array(21066);
		when "0101001001001011" => data_out <= rom_array(21067);
		when "0101001001001100" => data_out <= rom_array(21068);
		when "0101001001001101" => data_out <= rom_array(21069);
		when "0101001001001110" => data_out <= rom_array(21070);
		when "0101001001001111" => data_out <= rom_array(21071);
		when "0101001001010000" => data_out <= rom_array(21072);
		when "0101001001010001" => data_out <= rom_array(21073);
		when "0101001001010010" => data_out <= rom_array(21074);
		when "0101001001010011" => data_out <= rom_array(21075);
		when "0101001001010100" => data_out <= rom_array(21076);
		when "0101001001010101" => data_out <= rom_array(21077);
		when "0101001001010110" => data_out <= rom_array(21078);
		when "0101001001010111" => data_out <= rom_array(21079);
		when "0101001001011000" => data_out <= rom_array(21080);
		when "0101001001011001" => data_out <= rom_array(21081);
		when "0101001001011010" => data_out <= rom_array(21082);
		when "0101001001011011" => data_out <= rom_array(21083);
		when "0101001001011100" => data_out <= rom_array(21084);
		when "0101001001011101" => data_out <= rom_array(21085);
		when "0101001001011110" => data_out <= rom_array(21086);
		when "0101001001011111" => data_out <= rom_array(21087);
		when "0101001001100000" => data_out <= rom_array(21088);
		when "0101001001100001" => data_out <= rom_array(21089);
		when "0101001001100010" => data_out <= rom_array(21090);
		when "0101001001100011" => data_out <= rom_array(21091);
		when "0101001001100100" => data_out <= rom_array(21092);
		when "0101001001100101" => data_out <= rom_array(21093);
		when "0101001001100110" => data_out <= rom_array(21094);
		when "0101001001100111" => data_out <= rom_array(21095);
		when "0101001001101000" => data_out <= rom_array(21096);
		when "0101001001101001" => data_out <= rom_array(21097);
		when "0101001001101010" => data_out <= rom_array(21098);
		when "0101001001101011" => data_out <= rom_array(21099);
		when "0101001001101100" => data_out <= rom_array(21100);
		when "0101001001101101" => data_out <= rom_array(21101);
		when "0101001001101110" => data_out <= rom_array(21102);
		when "0101001001101111" => data_out <= rom_array(21103);
		when "0101001001110000" => data_out <= rom_array(21104);
		when "0101001001110001" => data_out <= rom_array(21105);
		when "0101001001110010" => data_out <= rom_array(21106);
		when "0101001001110011" => data_out <= rom_array(21107);
		when "0101001001110100" => data_out <= rom_array(21108);
		when "0101001001110101" => data_out <= rom_array(21109);
		when "0101001001110110" => data_out <= rom_array(21110);
		when "0101001001110111" => data_out <= rom_array(21111);
		when "0101001001111000" => data_out <= rom_array(21112);
		when "0101001001111001" => data_out <= rom_array(21113);
		when "0101001001111010" => data_out <= rom_array(21114);
		when "0101001001111011" => data_out <= rom_array(21115);
		when "0101001001111100" => data_out <= rom_array(21116);
		when "0101001001111101" => data_out <= rom_array(21117);
		when "0101001001111110" => data_out <= rom_array(21118);
		when "0101001001111111" => data_out <= rom_array(21119);
		when "0101001010000000" => data_out <= rom_array(21120);
		when "0101001010000001" => data_out <= rom_array(21121);
		when "0101001010000010" => data_out <= rom_array(21122);
		when "0101001010000011" => data_out <= rom_array(21123);
		when "0101001010000100" => data_out <= rom_array(21124);
		when "0101001010000101" => data_out <= rom_array(21125);
		when "0101001010000110" => data_out <= rom_array(21126);
		when "0101001010000111" => data_out <= rom_array(21127);
		when "0101001010001000" => data_out <= rom_array(21128);
		when "0101001010001001" => data_out <= rom_array(21129);
		when "0101001010001010" => data_out <= rom_array(21130);
		when "0101001010001011" => data_out <= rom_array(21131);
		when "0101001010001100" => data_out <= rom_array(21132);
		when "0101001010001101" => data_out <= rom_array(21133);
		when "0101001010001110" => data_out <= rom_array(21134);
		when "0101001010001111" => data_out <= rom_array(21135);
		when "0101001010010000" => data_out <= rom_array(21136);
		when "0101001010010001" => data_out <= rom_array(21137);
		when "0101001010010010" => data_out <= rom_array(21138);
		when "0101001010010011" => data_out <= rom_array(21139);
		when "0101001010010100" => data_out <= rom_array(21140);
		when "0101001010010101" => data_out <= rom_array(21141);
		when "0101001010010110" => data_out <= rom_array(21142);
		when "0101001010010111" => data_out <= rom_array(21143);
		when "0101001010011000" => data_out <= rom_array(21144);
		when "0101001010011001" => data_out <= rom_array(21145);
		when "0101001010011010" => data_out <= rom_array(21146);
		when "0101001010011011" => data_out <= rom_array(21147);
		when "0101001010011100" => data_out <= rom_array(21148);
		when "0101001010011101" => data_out <= rom_array(21149);
		when "0101001010011110" => data_out <= rom_array(21150);
		when "0101001010011111" => data_out <= rom_array(21151);
		when "0101001010100000" => data_out <= rom_array(21152);
		when "0101001010100001" => data_out <= rom_array(21153);
		when "0101001010100010" => data_out <= rom_array(21154);
		when "0101001010100011" => data_out <= rom_array(21155);
		when "0101001010100100" => data_out <= rom_array(21156);
		when "0101001010100101" => data_out <= rom_array(21157);
		when "0101001010100110" => data_out <= rom_array(21158);
		when "0101001010100111" => data_out <= rom_array(21159);
		when "0101001010101000" => data_out <= rom_array(21160);
		when "0101001010101001" => data_out <= rom_array(21161);
		when "0101001010101010" => data_out <= rom_array(21162);
		when "0101001010101011" => data_out <= rom_array(21163);
		when "0101001010101100" => data_out <= rom_array(21164);
		when "0101001010101101" => data_out <= rom_array(21165);
		when "0101001010101110" => data_out <= rom_array(21166);
		when "0101001010101111" => data_out <= rom_array(21167);
		when "0101001010110000" => data_out <= rom_array(21168);
		when "0101001010110001" => data_out <= rom_array(21169);
		when "0101001010110010" => data_out <= rom_array(21170);
		when "0101001010110011" => data_out <= rom_array(21171);
		when "0101001010110100" => data_out <= rom_array(21172);
		when "0101001010110101" => data_out <= rom_array(21173);
		when "0101001010110110" => data_out <= rom_array(21174);
		when "0101001010110111" => data_out <= rom_array(21175);
		when "0101001010111000" => data_out <= rom_array(21176);
		when "0101001010111001" => data_out <= rom_array(21177);
		when "0101001010111010" => data_out <= rom_array(21178);
		when "0101001010111011" => data_out <= rom_array(21179);
		when "0101001010111100" => data_out <= rom_array(21180);
		when "0101001010111101" => data_out <= rom_array(21181);
		when "0101001010111110" => data_out <= rom_array(21182);
		when "0101001010111111" => data_out <= rom_array(21183);
		when "0101001011000000" => data_out <= rom_array(21184);
		when "0101001011000001" => data_out <= rom_array(21185);
		when "0101001011000010" => data_out <= rom_array(21186);
		when "0101001011000011" => data_out <= rom_array(21187);
		when "0101001011000100" => data_out <= rom_array(21188);
		when "0101001011000101" => data_out <= rom_array(21189);
		when "0101001011000110" => data_out <= rom_array(21190);
		when "0101001011000111" => data_out <= rom_array(21191);
		when "0101001011001000" => data_out <= rom_array(21192);
		when "0101001011001001" => data_out <= rom_array(21193);
		when "0101001011001010" => data_out <= rom_array(21194);
		when "0101001011001011" => data_out <= rom_array(21195);
		when "0101001011001100" => data_out <= rom_array(21196);
		when "0101001011001101" => data_out <= rom_array(21197);
		when "0101001011001110" => data_out <= rom_array(21198);
		when "0101001011001111" => data_out <= rom_array(21199);
		when "0101001011010000" => data_out <= rom_array(21200);
		when "0101001011010001" => data_out <= rom_array(21201);
		when "0101001011010010" => data_out <= rom_array(21202);
		when "0101001011010011" => data_out <= rom_array(21203);
		when "0101001011010100" => data_out <= rom_array(21204);
		when "0101001011010101" => data_out <= rom_array(21205);
		when "0101001011010110" => data_out <= rom_array(21206);
		when "0101001011010111" => data_out <= rom_array(21207);
		when "0101001011011000" => data_out <= rom_array(21208);
		when "0101001011011001" => data_out <= rom_array(21209);
		when "0101001011011010" => data_out <= rom_array(21210);
		when "0101001011011011" => data_out <= rom_array(21211);
		when "0101001011011100" => data_out <= rom_array(21212);
		when "0101001011011101" => data_out <= rom_array(21213);
		when "0101001011011110" => data_out <= rom_array(21214);
		when "0101001011011111" => data_out <= rom_array(21215);
		when "0101001011100000" => data_out <= rom_array(21216);
		when "0101001011100001" => data_out <= rom_array(21217);
		when "0101001011100010" => data_out <= rom_array(21218);
		when "0101001011100011" => data_out <= rom_array(21219);
		when "0101001011100100" => data_out <= rom_array(21220);
		when "0101001011100101" => data_out <= rom_array(21221);
		when "0101001011100110" => data_out <= rom_array(21222);
		when "0101001011100111" => data_out <= rom_array(21223);
		when "0101001011101000" => data_out <= rom_array(21224);
		when "0101001011101001" => data_out <= rom_array(21225);
		when "0101001011101010" => data_out <= rom_array(21226);
		when "0101001011101011" => data_out <= rom_array(21227);
		when "0101001011101100" => data_out <= rom_array(21228);
		when "0101001011101101" => data_out <= rom_array(21229);
		when "0101001011101110" => data_out <= rom_array(21230);
		when "0101001011101111" => data_out <= rom_array(21231);
		when "0101001011110000" => data_out <= rom_array(21232);
		when "0101001011110001" => data_out <= rom_array(21233);
		when "0101001011110010" => data_out <= rom_array(21234);
		when "0101001011110011" => data_out <= rom_array(21235);
		when "0101001011110100" => data_out <= rom_array(21236);
		when "0101001011110101" => data_out <= rom_array(21237);
		when "0101001011110110" => data_out <= rom_array(21238);
		when "0101001011110111" => data_out <= rom_array(21239);
		when "0101001011111000" => data_out <= rom_array(21240);
		when "0101001011111001" => data_out <= rom_array(21241);
		when "0101001011111010" => data_out <= rom_array(21242);
		when "0101001011111011" => data_out <= rom_array(21243);
		when "0101001011111100" => data_out <= rom_array(21244);
		when "0101001011111101" => data_out <= rom_array(21245);
		when "0101001011111110" => data_out <= rom_array(21246);
		when "0101001011111111" => data_out <= rom_array(21247);
		when "0101001100000000" => data_out <= rom_array(21248);
		when "0101001100000001" => data_out <= rom_array(21249);
		when "0101001100000010" => data_out <= rom_array(21250);
		when "0101001100000011" => data_out <= rom_array(21251);
		when "0101001100000100" => data_out <= rom_array(21252);
		when "0101001100000101" => data_out <= rom_array(21253);
		when "0101001100000110" => data_out <= rom_array(21254);
		when "0101001100000111" => data_out <= rom_array(21255);
		when "0101001100001000" => data_out <= rom_array(21256);
		when "0101001100001001" => data_out <= rom_array(21257);
		when "0101001100001010" => data_out <= rom_array(21258);
		when "0101001100001011" => data_out <= rom_array(21259);
		when "0101001100001100" => data_out <= rom_array(21260);
		when "0101001100001101" => data_out <= rom_array(21261);
		when "0101001100001110" => data_out <= rom_array(21262);
		when "0101001100001111" => data_out <= rom_array(21263);
		when "0101001100010000" => data_out <= rom_array(21264);
		when "0101001100010001" => data_out <= rom_array(21265);
		when "0101001100010010" => data_out <= rom_array(21266);
		when "0101001100010011" => data_out <= rom_array(21267);
		when "0101001100010100" => data_out <= rom_array(21268);
		when "0101001100010101" => data_out <= rom_array(21269);
		when "0101001100010110" => data_out <= rom_array(21270);
		when "0101001100010111" => data_out <= rom_array(21271);
		when "0101001100011000" => data_out <= rom_array(21272);
		when "0101001100011001" => data_out <= rom_array(21273);
		when "0101001100011010" => data_out <= rom_array(21274);
		when "0101001100011011" => data_out <= rom_array(21275);
		when "0101001100011100" => data_out <= rom_array(21276);
		when "0101001100011101" => data_out <= rom_array(21277);
		when "0101001100011110" => data_out <= rom_array(21278);
		when "0101001100011111" => data_out <= rom_array(21279);
		when "0101001100100000" => data_out <= rom_array(21280);
		when "0101001100100001" => data_out <= rom_array(21281);
		when "0101001100100010" => data_out <= rom_array(21282);
		when "0101001100100011" => data_out <= rom_array(21283);
		when "0101001100100100" => data_out <= rom_array(21284);
		when "0101001100100101" => data_out <= rom_array(21285);
		when "0101001100100110" => data_out <= rom_array(21286);
		when "0101001100100111" => data_out <= rom_array(21287);
		when "0101001100101000" => data_out <= rom_array(21288);
		when "0101001100101001" => data_out <= rom_array(21289);
		when "0101001100101010" => data_out <= rom_array(21290);
		when "0101001100101011" => data_out <= rom_array(21291);
		when "0101001100101100" => data_out <= rom_array(21292);
		when "0101001100101101" => data_out <= rom_array(21293);
		when "0101001100101110" => data_out <= rom_array(21294);
		when "0101001100101111" => data_out <= rom_array(21295);
		when "0101001100110000" => data_out <= rom_array(21296);
		when "0101001100110001" => data_out <= rom_array(21297);
		when "0101001100110010" => data_out <= rom_array(21298);
		when "0101001100110011" => data_out <= rom_array(21299);
		when "0101001100110100" => data_out <= rom_array(21300);
		when "0101001100110101" => data_out <= rom_array(21301);
		when "0101001100110110" => data_out <= rom_array(21302);
		when "0101001100110111" => data_out <= rom_array(21303);
		when "0101001100111000" => data_out <= rom_array(21304);
		when "0101001100111001" => data_out <= rom_array(21305);
		when "0101001100111010" => data_out <= rom_array(21306);
		when "0101001100111011" => data_out <= rom_array(21307);
		when "0101001100111100" => data_out <= rom_array(21308);
		when "0101001100111101" => data_out <= rom_array(21309);
		when "0101001100111110" => data_out <= rom_array(21310);
		when "0101001100111111" => data_out <= rom_array(21311);
		when "0101001101000000" => data_out <= rom_array(21312);
		when "0101001101000001" => data_out <= rom_array(21313);
		when "0101001101000010" => data_out <= rom_array(21314);
		when "0101001101000011" => data_out <= rom_array(21315);
		when "0101001101000100" => data_out <= rom_array(21316);
		when "0101001101000101" => data_out <= rom_array(21317);
		when "0101001101000110" => data_out <= rom_array(21318);
		when "0101001101000111" => data_out <= rom_array(21319);
		when "0101001101001000" => data_out <= rom_array(21320);
		when "0101001101001001" => data_out <= rom_array(21321);
		when "0101001101001010" => data_out <= rom_array(21322);
		when "0101001101001011" => data_out <= rom_array(21323);
		when "0101001101001100" => data_out <= rom_array(21324);
		when "0101001101001101" => data_out <= rom_array(21325);
		when "0101001101001110" => data_out <= rom_array(21326);
		when "0101001101001111" => data_out <= rom_array(21327);
		when "0101001101010000" => data_out <= rom_array(21328);
		when "0101001101010001" => data_out <= rom_array(21329);
		when "0101001101010010" => data_out <= rom_array(21330);
		when "0101001101010011" => data_out <= rom_array(21331);
		when "0101001101010100" => data_out <= rom_array(21332);
		when "0101001101010101" => data_out <= rom_array(21333);
		when "0101001101010110" => data_out <= rom_array(21334);
		when "0101001101010111" => data_out <= rom_array(21335);
		when "0101001101011000" => data_out <= rom_array(21336);
		when "0101001101011001" => data_out <= rom_array(21337);
		when "0101001101011010" => data_out <= rom_array(21338);
		when "0101001101011011" => data_out <= rom_array(21339);
		when "0101001101011100" => data_out <= rom_array(21340);
		when "0101001101011101" => data_out <= rom_array(21341);
		when "0101001101011110" => data_out <= rom_array(21342);
		when "0101001101011111" => data_out <= rom_array(21343);
		when "0101001101100000" => data_out <= rom_array(21344);
		when "0101001101100001" => data_out <= rom_array(21345);
		when "0101001101100010" => data_out <= rom_array(21346);
		when "0101001101100011" => data_out <= rom_array(21347);
		when "0101001101100100" => data_out <= rom_array(21348);
		when "0101001101100101" => data_out <= rom_array(21349);
		when "0101001101100110" => data_out <= rom_array(21350);
		when "0101001101100111" => data_out <= rom_array(21351);
		when "0101001101101000" => data_out <= rom_array(21352);
		when "0101001101101001" => data_out <= rom_array(21353);
		when "0101001101101010" => data_out <= rom_array(21354);
		when "0101001101101011" => data_out <= rom_array(21355);
		when "0101001101101100" => data_out <= rom_array(21356);
		when "0101001101101101" => data_out <= rom_array(21357);
		when "0101001101101110" => data_out <= rom_array(21358);
		when "0101001101101111" => data_out <= rom_array(21359);
		when "0101001101110000" => data_out <= rom_array(21360);
		when "0101001101110001" => data_out <= rom_array(21361);
		when "0101001101110010" => data_out <= rom_array(21362);
		when "0101001101110011" => data_out <= rom_array(21363);
		when "0101001101110100" => data_out <= rom_array(21364);
		when "0101001101110101" => data_out <= rom_array(21365);
		when "0101001101110110" => data_out <= rom_array(21366);
		when "0101001101110111" => data_out <= rom_array(21367);
		when "0101001101111000" => data_out <= rom_array(21368);
		when "0101001101111001" => data_out <= rom_array(21369);
		when "0101001101111010" => data_out <= rom_array(21370);
		when "0101001101111011" => data_out <= rom_array(21371);
		when "0101001101111100" => data_out <= rom_array(21372);
		when "0101001101111101" => data_out <= rom_array(21373);
		when "0101001101111110" => data_out <= rom_array(21374);
		when "0101001101111111" => data_out <= rom_array(21375);
		when "0101001110000000" => data_out <= rom_array(21376);
		when "0101001110000001" => data_out <= rom_array(21377);
		when "0101001110000010" => data_out <= rom_array(21378);
		when "0101001110000011" => data_out <= rom_array(21379);
		when "0101001110000100" => data_out <= rom_array(21380);
		when "0101001110000101" => data_out <= rom_array(21381);
		when "0101001110000110" => data_out <= rom_array(21382);
		when "0101001110000111" => data_out <= rom_array(21383);
		when "0101001110001000" => data_out <= rom_array(21384);
		when "0101001110001001" => data_out <= rom_array(21385);
		when "0101001110001010" => data_out <= rom_array(21386);
		when "0101001110001011" => data_out <= rom_array(21387);
		when "0101001110001100" => data_out <= rom_array(21388);
		when "0101001110001101" => data_out <= rom_array(21389);
		when "0101001110001110" => data_out <= rom_array(21390);
		when "0101001110001111" => data_out <= rom_array(21391);
		when "0101001110010000" => data_out <= rom_array(21392);
		when "0101001110010001" => data_out <= rom_array(21393);
		when "0101001110010010" => data_out <= rom_array(21394);
		when "0101001110010011" => data_out <= rom_array(21395);
		when "0101001110010100" => data_out <= rom_array(21396);
		when "0101001110010101" => data_out <= rom_array(21397);
		when "0101001110010110" => data_out <= rom_array(21398);
		when "0101001110010111" => data_out <= rom_array(21399);
		when "0101001110011000" => data_out <= rom_array(21400);
		when "0101001110011001" => data_out <= rom_array(21401);
		when "0101001110011010" => data_out <= rom_array(21402);
		when "0101001110011011" => data_out <= rom_array(21403);
		when "0101001110011100" => data_out <= rom_array(21404);
		when "0101001110011101" => data_out <= rom_array(21405);
		when "0101001110011110" => data_out <= rom_array(21406);
		when "0101001110011111" => data_out <= rom_array(21407);
		when "0101001110100000" => data_out <= rom_array(21408);
		when "0101001110100001" => data_out <= rom_array(21409);
		when "0101001110100010" => data_out <= rom_array(21410);
		when "0101001110100011" => data_out <= rom_array(21411);
		when "0101001110100100" => data_out <= rom_array(21412);
		when "0101001110100101" => data_out <= rom_array(21413);
		when "0101001110100110" => data_out <= rom_array(21414);
		when "0101001110100111" => data_out <= rom_array(21415);
		when "0101001110101000" => data_out <= rom_array(21416);
		when "0101001110101001" => data_out <= rom_array(21417);
		when "0101001110101010" => data_out <= rom_array(21418);
		when "0101001110101011" => data_out <= rom_array(21419);
		when "0101001110101100" => data_out <= rom_array(21420);
		when "0101001110101101" => data_out <= rom_array(21421);
		when "0101001110101110" => data_out <= rom_array(21422);
		when "0101001110101111" => data_out <= rom_array(21423);
		when "0101001110110000" => data_out <= rom_array(21424);
		when "0101001110110001" => data_out <= rom_array(21425);
		when "0101001110110010" => data_out <= rom_array(21426);
		when "0101001110110011" => data_out <= rom_array(21427);
		when "0101001110110100" => data_out <= rom_array(21428);
		when "0101001110110101" => data_out <= rom_array(21429);
		when "0101001110110110" => data_out <= rom_array(21430);
		when "0101001110110111" => data_out <= rom_array(21431);
		when "0101001110111000" => data_out <= rom_array(21432);
		when "0101001110111001" => data_out <= rom_array(21433);
		when "0101001110111010" => data_out <= rom_array(21434);
		when "0101001110111011" => data_out <= rom_array(21435);
		when "0101001110111100" => data_out <= rom_array(21436);
		when "0101001110111101" => data_out <= rom_array(21437);
		when "0101001110111110" => data_out <= rom_array(21438);
		when "0101001110111111" => data_out <= rom_array(21439);
		when "0101001111000000" => data_out <= rom_array(21440);
		when "0101001111000001" => data_out <= rom_array(21441);
		when "0101001111000010" => data_out <= rom_array(21442);
		when "0101001111000011" => data_out <= rom_array(21443);
		when "0101001111000100" => data_out <= rom_array(21444);
		when "0101001111000101" => data_out <= rom_array(21445);
		when "0101001111000110" => data_out <= rom_array(21446);
		when "0101001111000111" => data_out <= rom_array(21447);
		when "0101001111001000" => data_out <= rom_array(21448);
		when "0101001111001001" => data_out <= rom_array(21449);
		when "0101001111001010" => data_out <= rom_array(21450);
		when "0101001111001011" => data_out <= rom_array(21451);
		when "0101001111001100" => data_out <= rom_array(21452);
		when "0101001111001101" => data_out <= rom_array(21453);
		when "0101001111001110" => data_out <= rom_array(21454);
		when "0101001111001111" => data_out <= rom_array(21455);
		when "0101001111010000" => data_out <= rom_array(21456);
		when "0101001111010001" => data_out <= rom_array(21457);
		when "0101001111010010" => data_out <= rom_array(21458);
		when "0101001111010011" => data_out <= rom_array(21459);
		when "0101001111010100" => data_out <= rom_array(21460);
		when "0101001111010101" => data_out <= rom_array(21461);
		when "0101001111010110" => data_out <= rom_array(21462);
		when "0101001111010111" => data_out <= rom_array(21463);
		when "0101001111011000" => data_out <= rom_array(21464);
		when "0101001111011001" => data_out <= rom_array(21465);
		when "0101001111011010" => data_out <= rom_array(21466);
		when "0101001111011011" => data_out <= rom_array(21467);
		when "0101001111011100" => data_out <= rom_array(21468);
		when "0101001111011101" => data_out <= rom_array(21469);
		when "0101001111011110" => data_out <= rom_array(21470);
		when "0101001111011111" => data_out <= rom_array(21471);
		when "0101001111100000" => data_out <= rom_array(21472);
		when "0101001111100001" => data_out <= rom_array(21473);
		when "0101001111100010" => data_out <= rom_array(21474);
		when "0101001111100011" => data_out <= rom_array(21475);
		when "0101001111100100" => data_out <= rom_array(21476);
		when "0101001111100101" => data_out <= rom_array(21477);
		when "0101001111100110" => data_out <= rom_array(21478);
		when "0101001111100111" => data_out <= rom_array(21479);
		when "0101001111101000" => data_out <= rom_array(21480);
		when "0101001111101001" => data_out <= rom_array(21481);
		when "0101001111101010" => data_out <= rom_array(21482);
		when "0101001111101011" => data_out <= rom_array(21483);
		when "0101001111101100" => data_out <= rom_array(21484);
		when "0101001111101101" => data_out <= rom_array(21485);
		when "0101001111101110" => data_out <= rom_array(21486);
		when "0101001111101111" => data_out <= rom_array(21487);
		when "0101001111110000" => data_out <= rom_array(21488);
		when "0101001111110001" => data_out <= rom_array(21489);
		when "0101001111110010" => data_out <= rom_array(21490);
		when "0101001111110011" => data_out <= rom_array(21491);
		when "0101001111110100" => data_out <= rom_array(21492);
		when "0101001111110101" => data_out <= rom_array(21493);
		when "0101001111110110" => data_out <= rom_array(21494);
		when "0101001111110111" => data_out <= rom_array(21495);
		when "0101001111111000" => data_out <= rom_array(21496);
		when "0101001111111001" => data_out <= rom_array(21497);
		when "0101001111111010" => data_out <= rom_array(21498);
		when "0101001111111011" => data_out <= rom_array(21499);
		when "0101001111111100" => data_out <= rom_array(21500);
		when "0101001111111101" => data_out <= rom_array(21501);
		when "0101001111111110" => data_out <= rom_array(21502);
		when "0101001111111111" => data_out <= rom_array(21503);
		when "0101010000000000" => data_out <= rom_array(21504);
		when "0101010000000001" => data_out <= rom_array(21505);
		when "0101010000000010" => data_out <= rom_array(21506);
		when "0101010000000011" => data_out <= rom_array(21507);
		when "0101010000000100" => data_out <= rom_array(21508);
		when "0101010000000101" => data_out <= rom_array(21509);
		when "0101010000000110" => data_out <= rom_array(21510);
		when "0101010000000111" => data_out <= rom_array(21511);
		when "0101010000001000" => data_out <= rom_array(21512);
		when "0101010000001001" => data_out <= rom_array(21513);
		when "0101010000001010" => data_out <= rom_array(21514);
		when "0101010000001011" => data_out <= rom_array(21515);
		when "0101010000001100" => data_out <= rom_array(21516);
		when "0101010000001101" => data_out <= rom_array(21517);
		when "0101010000001110" => data_out <= rom_array(21518);
		when "0101010000001111" => data_out <= rom_array(21519);
		when "0101010000010000" => data_out <= rom_array(21520);
		when "0101010000010001" => data_out <= rom_array(21521);
		when "0101010000010010" => data_out <= rom_array(21522);
		when "0101010000010011" => data_out <= rom_array(21523);
		when "0101010000010100" => data_out <= rom_array(21524);
		when "0101010000010101" => data_out <= rom_array(21525);
		when "0101010000010110" => data_out <= rom_array(21526);
		when "0101010000010111" => data_out <= rom_array(21527);
		when "0101010000011000" => data_out <= rom_array(21528);
		when "0101010000011001" => data_out <= rom_array(21529);
		when "0101010000011010" => data_out <= rom_array(21530);
		when "0101010000011011" => data_out <= rom_array(21531);
		when "0101010000011100" => data_out <= rom_array(21532);
		when "0101010000011101" => data_out <= rom_array(21533);
		when "0101010000011110" => data_out <= rom_array(21534);
		when "0101010000011111" => data_out <= rom_array(21535);
		when "0101010000100000" => data_out <= rom_array(21536);
		when "0101010000100001" => data_out <= rom_array(21537);
		when "0101010000100010" => data_out <= rom_array(21538);
		when "0101010000100011" => data_out <= rom_array(21539);
		when "0101010000100100" => data_out <= rom_array(21540);
		when "0101010000100101" => data_out <= rom_array(21541);
		when "0101010000100110" => data_out <= rom_array(21542);
		when "0101010000100111" => data_out <= rom_array(21543);
		when "0101010000101000" => data_out <= rom_array(21544);
		when "0101010000101001" => data_out <= rom_array(21545);
		when "0101010000101010" => data_out <= rom_array(21546);
		when "0101010000101011" => data_out <= rom_array(21547);
		when "0101010000101100" => data_out <= rom_array(21548);
		when "0101010000101101" => data_out <= rom_array(21549);
		when "0101010000101110" => data_out <= rom_array(21550);
		when "0101010000101111" => data_out <= rom_array(21551);
		when "0101010000110000" => data_out <= rom_array(21552);
		when "0101010000110001" => data_out <= rom_array(21553);
		when "0101010000110010" => data_out <= rom_array(21554);
		when "0101010000110011" => data_out <= rom_array(21555);
		when "0101010000110100" => data_out <= rom_array(21556);
		when "0101010000110101" => data_out <= rom_array(21557);
		when "0101010000110110" => data_out <= rom_array(21558);
		when "0101010000110111" => data_out <= rom_array(21559);
		when "0101010000111000" => data_out <= rom_array(21560);
		when "0101010000111001" => data_out <= rom_array(21561);
		when "0101010000111010" => data_out <= rom_array(21562);
		when "0101010000111011" => data_out <= rom_array(21563);
		when "0101010000111100" => data_out <= rom_array(21564);
		when "0101010000111101" => data_out <= rom_array(21565);
		when "0101010000111110" => data_out <= rom_array(21566);
		when "0101010000111111" => data_out <= rom_array(21567);
		when "0101010001000000" => data_out <= rom_array(21568);
		when "0101010001000001" => data_out <= rom_array(21569);
		when "0101010001000010" => data_out <= rom_array(21570);
		when "0101010001000011" => data_out <= rom_array(21571);
		when "0101010001000100" => data_out <= rom_array(21572);
		when "0101010001000101" => data_out <= rom_array(21573);
		when "0101010001000110" => data_out <= rom_array(21574);
		when "0101010001000111" => data_out <= rom_array(21575);
		when "0101010001001000" => data_out <= rom_array(21576);
		when "0101010001001001" => data_out <= rom_array(21577);
		when "0101010001001010" => data_out <= rom_array(21578);
		when "0101010001001011" => data_out <= rom_array(21579);
		when "0101010001001100" => data_out <= rom_array(21580);
		when "0101010001001101" => data_out <= rom_array(21581);
		when "0101010001001110" => data_out <= rom_array(21582);
		when "0101010001001111" => data_out <= rom_array(21583);
		when "0101010001010000" => data_out <= rom_array(21584);
		when "0101010001010001" => data_out <= rom_array(21585);
		when "0101010001010010" => data_out <= rom_array(21586);
		when "0101010001010011" => data_out <= rom_array(21587);
		when "0101010001010100" => data_out <= rom_array(21588);
		when "0101010001010101" => data_out <= rom_array(21589);
		when "0101010001010110" => data_out <= rom_array(21590);
		when "0101010001010111" => data_out <= rom_array(21591);
		when "0101010001011000" => data_out <= rom_array(21592);
		when "0101010001011001" => data_out <= rom_array(21593);
		when "0101010001011010" => data_out <= rom_array(21594);
		when "0101010001011011" => data_out <= rom_array(21595);
		when "0101010001011100" => data_out <= rom_array(21596);
		when "0101010001011101" => data_out <= rom_array(21597);
		when "0101010001011110" => data_out <= rom_array(21598);
		when "0101010001011111" => data_out <= rom_array(21599);
		when "0101010001100000" => data_out <= rom_array(21600);
		when "0101010001100001" => data_out <= rom_array(21601);
		when "0101010001100010" => data_out <= rom_array(21602);
		when "0101010001100011" => data_out <= rom_array(21603);
		when "0101010001100100" => data_out <= rom_array(21604);
		when "0101010001100101" => data_out <= rom_array(21605);
		when "0101010001100110" => data_out <= rom_array(21606);
		when "0101010001100111" => data_out <= rom_array(21607);
		when "0101010001101000" => data_out <= rom_array(21608);
		when "0101010001101001" => data_out <= rom_array(21609);
		when "0101010001101010" => data_out <= rom_array(21610);
		when "0101010001101011" => data_out <= rom_array(21611);
		when "0101010001101100" => data_out <= rom_array(21612);
		when "0101010001101101" => data_out <= rom_array(21613);
		when "0101010001101110" => data_out <= rom_array(21614);
		when "0101010001101111" => data_out <= rom_array(21615);
		when "0101010001110000" => data_out <= rom_array(21616);
		when "0101010001110001" => data_out <= rom_array(21617);
		when "0101010001110010" => data_out <= rom_array(21618);
		when "0101010001110011" => data_out <= rom_array(21619);
		when "0101010001110100" => data_out <= rom_array(21620);
		when "0101010001110101" => data_out <= rom_array(21621);
		when "0101010001110110" => data_out <= rom_array(21622);
		when "0101010001110111" => data_out <= rom_array(21623);
		when "0101010001111000" => data_out <= rom_array(21624);
		when "0101010001111001" => data_out <= rom_array(21625);
		when "0101010001111010" => data_out <= rom_array(21626);
		when "0101010001111011" => data_out <= rom_array(21627);
		when "0101010001111100" => data_out <= rom_array(21628);
		when "0101010001111101" => data_out <= rom_array(21629);
		when "0101010001111110" => data_out <= rom_array(21630);
		when "0101010001111111" => data_out <= rom_array(21631);
		when "0101010010000000" => data_out <= rom_array(21632);
		when "0101010010000001" => data_out <= rom_array(21633);
		when "0101010010000010" => data_out <= rom_array(21634);
		when "0101010010000011" => data_out <= rom_array(21635);
		when "0101010010000100" => data_out <= rom_array(21636);
		when "0101010010000101" => data_out <= rom_array(21637);
		when "0101010010000110" => data_out <= rom_array(21638);
		when "0101010010000111" => data_out <= rom_array(21639);
		when "0101010010001000" => data_out <= rom_array(21640);
		when "0101010010001001" => data_out <= rom_array(21641);
		when "0101010010001010" => data_out <= rom_array(21642);
		when "0101010010001011" => data_out <= rom_array(21643);
		when "0101010010001100" => data_out <= rom_array(21644);
		when "0101010010001101" => data_out <= rom_array(21645);
		when "0101010010001110" => data_out <= rom_array(21646);
		when "0101010010001111" => data_out <= rom_array(21647);
		when "0101010010010000" => data_out <= rom_array(21648);
		when "0101010010010001" => data_out <= rom_array(21649);
		when "0101010010010010" => data_out <= rom_array(21650);
		when "0101010010010011" => data_out <= rom_array(21651);
		when "0101010010010100" => data_out <= rom_array(21652);
		when "0101010010010101" => data_out <= rom_array(21653);
		when "0101010010010110" => data_out <= rom_array(21654);
		when "0101010010010111" => data_out <= rom_array(21655);
		when "0101010010011000" => data_out <= rom_array(21656);
		when "0101010010011001" => data_out <= rom_array(21657);
		when "0101010010011010" => data_out <= rom_array(21658);
		when "0101010010011011" => data_out <= rom_array(21659);
		when "0101010010011100" => data_out <= rom_array(21660);
		when "0101010010011101" => data_out <= rom_array(21661);
		when "0101010010011110" => data_out <= rom_array(21662);
		when "0101010010011111" => data_out <= rom_array(21663);
		when "0101010010100000" => data_out <= rom_array(21664);
		when "0101010010100001" => data_out <= rom_array(21665);
		when "0101010010100010" => data_out <= rom_array(21666);
		when "0101010010100011" => data_out <= rom_array(21667);
		when "0101010010100100" => data_out <= rom_array(21668);
		when "0101010010100101" => data_out <= rom_array(21669);
		when "0101010010100110" => data_out <= rom_array(21670);
		when "0101010010100111" => data_out <= rom_array(21671);
		when "0101010010101000" => data_out <= rom_array(21672);
		when "0101010010101001" => data_out <= rom_array(21673);
		when "0101010010101010" => data_out <= rom_array(21674);
		when "0101010010101011" => data_out <= rom_array(21675);
		when "0101010010101100" => data_out <= rom_array(21676);
		when "0101010010101101" => data_out <= rom_array(21677);
		when "0101010010101110" => data_out <= rom_array(21678);
		when "0101010010101111" => data_out <= rom_array(21679);
		when "0101010010110000" => data_out <= rom_array(21680);
		when "0101010010110001" => data_out <= rom_array(21681);
		when "0101010010110010" => data_out <= rom_array(21682);
		when "0101010010110011" => data_out <= rom_array(21683);
		when "0101010010110100" => data_out <= rom_array(21684);
		when "0101010010110101" => data_out <= rom_array(21685);
		when "0101010010110110" => data_out <= rom_array(21686);
		when "0101010010110111" => data_out <= rom_array(21687);
		when "0101010010111000" => data_out <= rom_array(21688);
		when "0101010010111001" => data_out <= rom_array(21689);
		when "0101010010111010" => data_out <= rom_array(21690);
		when "0101010010111011" => data_out <= rom_array(21691);
		when "0101010010111100" => data_out <= rom_array(21692);
		when "0101010010111101" => data_out <= rom_array(21693);
		when "0101010010111110" => data_out <= rom_array(21694);
		when "0101010010111111" => data_out <= rom_array(21695);
		when "0101010011000000" => data_out <= rom_array(21696);
		when "0101010011000001" => data_out <= rom_array(21697);
		when "0101010011000010" => data_out <= rom_array(21698);
		when "0101010011000011" => data_out <= rom_array(21699);
		when "0101010011000100" => data_out <= rom_array(21700);
		when "0101010011000101" => data_out <= rom_array(21701);
		when "0101010011000110" => data_out <= rom_array(21702);
		when "0101010011000111" => data_out <= rom_array(21703);
		when "0101010011001000" => data_out <= rom_array(21704);
		when "0101010011001001" => data_out <= rom_array(21705);
		when "0101010011001010" => data_out <= rom_array(21706);
		when "0101010011001011" => data_out <= rom_array(21707);
		when "0101010011001100" => data_out <= rom_array(21708);
		when "0101010011001101" => data_out <= rom_array(21709);
		when "0101010011001110" => data_out <= rom_array(21710);
		when "0101010011001111" => data_out <= rom_array(21711);
		when "0101010011010000" => data_out <= rom_array(21712);
		when "0101010011010001" => data_out <= rom_array(21713);
		when "0101010011010010" => data_out <= rom_array(21714);
		when "0101010011010011" => data_out <= rom_array(21715);
		when "0101010011010100" => data_out <= rom_array(21716);
		when "0101010011010101" => data_out <= rom_array(21717);
		when "0101010011010110" => data_out <= rom_array(21718);
		when "0101010011010111" => data_out <= rom_array(21719);
		when "0101010011011000" => data_out <= rom_array(21720);
		when "0101010011011001" => data_out <= rom_array(21721);
		when "0101010011011010" => data_out <= rom_array(21722);
		when "0101010011011011" => data_out <= rom_array(21723);
		when "0101010011011100" => data_out <= rom_array(21724);
		when "0101010011011101" => data_out <= rom_array(21725);
		when "0101010011011110" => data_out <= rom_array(21726);
		when "0101010011011111" => data_out <= rom_array(21727);
		when "0101010011100000" => data_out <= rom_array(21728);
		when "0101010011100001" => data_out <= rom_array(21729);
		when "0101010011100010" => data_out <= rom_array(21730);
		when "0101010011100011" => data_out <= rom_array(21731);
		when "0101010011100100" => data_out <= rom_array(21732);
		when "0101010011100101" => data_out <= rom_array(21733);
		when "0101010011100110" => data_out <= rom_array(21734);
		when "0101010011100111" => data_out <= rom_array(21735);
		when "0101010011101000" => data_out <= rom_array(21736);
		when "0101010011101001" => data_out <= rom_array(21737);
		when "0101010011101010" => data_out <= rom_array(21738);
		when "0101010011101011" => data_out <= rom_array(21739);
		when "0101010011101100" => data_out <= rom_array(21740);
		when "0101010011101101" => data_out <= rom_array(21741);
		when "0101010011101110" => data_out <= rom_array(21742);
		when "0101010011101111" => data_out <= rom_array(21743);
		when "0101010011110000" => data_out <= rom_array(21744);
		when "0101010011110001" => data_out <= rom_array(21745);
		when "0101010011110010" => data_out <= rom_array(21746);
		when "0101010011110011" => data_out <= rom_array(21747);
		when "0101010011110100" => data_out <= rom_array(21748);
		when "0101010011110101" => data_out <= rom_array(21749);
		when "0101010011110110" => data_out <= rom_array(21750);
		when "0101010011110111" => data_out <= rom_array(21751);
		when "0101010011111000" => data_out <= rom_array(21752);
		when "0101010011111001" => data_out <= rom_array(21753);
		when "0101010011111010" => data_out <= rom_array(21754);
		when "0101010011111011" => data_out <= rom_array(21755);
		when "0101010011111100" => data_out <= rom_array(21756);
		when "0101010011111101" => data_out <= rom_array(21757);
		when "0101010011111110" => data_out <= rom_array(21758);
		when "0101010011111111" => data_out <= rom_array(21759);
		when "0101010100000000" => data_out <= rom_array(21760);
		when "0101010100000001" => data_out <= rom_array(21761);
		when "0101010100000010" => data_out <= rom_array(21762);
		when "0101010100000011" => data_out <= rom_array(21763);
		when "0101010100000100" => data_out <= rom_array(21764);
		when "0101010100000101" => data_out <= rom_array(21765);
		when "0101010100000110" => data_out <= rom_array(21766);
		when "0101010100000111" => data_out <= rom_array(21767);
		when "0101010100001000" => data_out <= rom_array(21768);
		when "0101010100001001" => data_out <= rom_array(21769);
		when "0101010100001010" => data_out <= rom_array(21770);
		when "0101010100001011" => data_out <= rom_array(21771);
		when "0101010100001100" => data_out <= rom_array(21772);
		when "0101010100001101" => data_out <= rom_array(21773);
		when "0101010100001110" => data_out <= rom_array(21774);
		when "0101010100001111" => data_out <= rom_array(21775);
		when "0101010100010000" => data_out <= rom_array(21776);
		when "0101010100010001" => data_out <= rom_array(21777);
		when "0101010100010010" => data_out <= rom_array(21778);
		when "0101010100010011" => data_out <= rom_array(21779);
		when "0101010100010100" => data_out <= rom_array(21780);
		when "0101010100010101" => data_out <= rom_array(21781);
		when "0101010100010110" => data_out <= rom_array(21782);
		when "0101010100010111" => data_out <= rom_array(21783);
		when "0101010100011000" => data_out <= rom_array(21784);
		when "0101010100011001" => data_out <= rom_array(21785);
		when "0101010100011010" => data_out <= rom_array(21786);
		when "0101010100011011" => data_out <= rom_array(21787);
		when "0101010100011100" => data_out <= rom_array(21788);
		when "0101010100011101" => data_out <= rom_array(21789);
		when "0101010100011110" => data_out <= rom_array(21790);
		when "0101010100011111" => data_out <= rom_array(21791);
		when "0101010100100000" => data_out <= rom_array(21792);
		when "0101010100100001" => data_out <= rom_array(21793);
		when "0101010100100010" => data_out <= rom_array(21794);
		when "0101010100100011" => data_out <= rom_array(21795);
		when "0101010100100100" => data_out <= rom_array(21796);
		when "0101010100100101" => data_out <= rom_array(21797);
		when "0101010100100110" => data_out <= rom_array(21798);
		when "0101010100100111" => data_out <= rom_array(21799);
		when "0101010100101000" => data_out <= rom_array(21800);
		when "0101010100101001" => data_out <= rom_array(21801);
		when "0101010100101010" => data_out <= rom_array(21802);
		when "0101010100101011" => data_out <= rom_array(21803);
		when "0101010100101100" => data_out <= rom_array(21804);
		when "0101010100101101" => data_out <= rom_array(21805);
		when "0101010100101110" => data_out <= rom_array(21806);
		when "0101010100101111" => data_out <= rom_array(21807);
		when "0101010100110000" => data_out <= rom_array(21808);
		when "0101010100110001" => data_out <= rom_array(21809);
		when "0101010100110010" => data_out <= rom_array(21810);
		when "0101010100110011" => data_out <= rom_array(21811);
		when "0101010100110100" => data_out <= rom_array(21812);
		when "0101010100110101" => data_out <= rom_array(21813);
		when "0101010100110110" => data_out <= rom_array(21814);
		when "0101010100110111" => data_out <= rom_array(21815);
		when "0101010100111000" => data_out <= rom_array(21816);
		when "0101010100111001" => data_out <= rom_array(21817);
		when "0101010100111010" => data_out <= rom_array(21818);
		when "0101010100111011" => data_out <= rom_array(21819);
		when "0101010100111100" => data_out <= rom_array(21820);
		when "0101010100111101" => data_out <= rom_array(21821);
		when "0101010100111110" => data_out <= rom_array(21822);
		when "0101010100111111" => data_out <= rom_array(21823);
		when "0101010101000000" => data_out <= rom_array(21824);
		when "0101010101000001" => data_out <= rom_array(21825);
		when "0101010101000010" => data_out <= rom_array(21826);
		when "0101010101000011" => data_out <= rom_array(21827);
		when "0101010101000100" => data_out <= rom_array(21828);
		when "0101010101000101" => data_out <= rom_array(21829);
		when "0101010101000110" => data_out <= rom_array(21830);
		when "0101010101000111" => data_out <= rom_array(21831);
		when "0101010101001000" => data_out <= rom_array(21832);
		when "0101010101001001" => data_out <= rom_array(21833);
		when "0101010101001010" => data_out <= rom_array(21834);
		when "0101010101001011" => data_out <= rom_array(21835);
		when "0101010101001100" => data_out <= rom_array(21836);
		when "0101010101001101" => data_out <= rom_array(21837);
		when "0101010101001110" => data_out <= rom_array(21838);
		when "0101010101001111" => data_out <= rom_array(21839);
		when "0101010101010000" => data_out <= rom_array(21840);
		when "0101010101010001" => data_out <= rom_array(21841);
		when "0101010101010010" => data_out <= rom_array(21842);
		when "0101010101010011" => data_out <= rom_array(21843);
		when "0101010101010100" => data_out <= rom_array(21844);
		when "0101010101010101" => data_out <= rom_array(21845);
		when "0101010101010110" => data_out <= rom_array(21846);
		when "0101010101010111" => data_out <= rom_array(21847);
		when "0101010101011000" => data_out <= rom_array(21848);
		when "0101010101011001" => data_out <= rom_array(21849);
		when "0101010101011010" => data_out <= rom_array(21850);
		when "0101010101011011" => data_out <= rom_array(21851);
		when "0101010101011100" => data_out <= rom_array(21852);
		when "0101010101011101" => data_out <= rom_array(21853);
		when "0101010101011110" => data_out <= rom_array(21854);
		when "0101010101011111" => data_out <= rom_array(21855);
		when "0101010101100000" => data_out <= rom_array(21856);
		when "0101010101100001" => data_out <= rom_array(21857);
		when "0101010101100010" => data_out <= rom_array(21858);
		when "0101010101100011" => data_out <= rom_array(21859);
		when "0101010101100100" => data_out <= rom_array(21860);
		when "0101010101100101" => data_out <= rom_array(21861);
		when "0101010101100110" => data_out <= rom_array(21862);
		when "0101010101100111" => data_out <= rom_array(21863);
		when "0101010101101000" => data_out <= rom_array(21864);
		when "0101010101101001" => data_out <= rom_array(21865);
		when "0101010101101010" => data_out <= rom_array(21866);
		when "0101010101101011" => data_out <= rom_array(21867);
		when "0101010101101100" => data_out <= rom_array(21868);
		when "0101010101101101" => data_out <= rom_array(21869);
		when "0101010101101110" => data_out <= rom_array(21870);
		when "0101010101101111" => data_out <= rom_array(21871);
		when "0101010101110000" => data_out <= rom_array(21872);
		when "0101010101110001" => data_out <= rom_array(21873);
		when "0101010101110010" => data_out <= rom_array(21874);
		when "0101010101110011" => data_out <= rom_array(21875);
		when "0101010101110100" => data_out <= rom_array(21876);
		when "0101010101110101" => data_out <= rom_array(21877);
		when "0101010101110110" => data_out <= rom_array(21878);
		when "0101010101110111" => data_out <= rom_array(21879);
		when "0101010101111000" => data_out <= rom_array(21880);
		when "0101010101111001" => data_out <= rom_array(21881);
		when "0101010101111010" => data_out <= rom_array(21882);
		when "0101010101111011" => data_out <= rom_array(21883);
		when "0101010101111100" => data_out <= rom_array(21884);
		when "0101010101111101" => data_out <= rom_array(21885);
		when "0101010101111110" => data_out <= rom_array(21886);
		when "0101010101111111" => data_out <= rom_array(21887);
		when "0101010110000000" => data_out <= rom_array(21888);
		when "0101010110000001" => data_out <= rom_array(21889);
		when "0101010110000010" => data_out <= rom_array(21890);
		when "0101010110000011" => data_out <= rom_array(21891);
		when "0101010110000100" => data_out <= rom_array(21892);
		when "0101010110000101" => data_out <= rom_array(21893);
		when "0101010110000110" => data_out <= rom_array(21894);
		when "0101010110000111" => data_out <= rom_array(21895);
		when "0101010110001000" => data_out <= rom_array(21896);
		when "0101010110001001" => data_out <= rom_array(21897);
		when "0101010110001010" => data_out <= rom_array(21898);
		when "0101010110001011" => data_out <= rom_array(21899);
		when "0101010110001100" => data_out <= rom_array(21900);
		when "0101010110001101" => data_out <= rom_array(21901);
		when "0101010110001110" => data_out <= rom_array(21902);
		when "0101010110001111" => data_out <= rom_array(21903);
		when "0101010110010000" => data_out <= rom_array(21904);
		when "0101010110010001" => data_out <= rom_array(21905);
		when "0101010110010010" => data_out <= rom_array(21906);
		when "0101010110010011" => data_out <= rom_array(21907);
		when "0101010110010100" => data_out <= rom_array(21908);
		when "0101010110010101" => data_out <= rom_array(21909);
		when "0101010110010110" => data_out <= rom_array(21910);
		when "0101010110010111" => data_out <= rom_array(21911);
		when "0101010110011000" => data_out <= rom_array(21912);
		when "0101010110011001" => data_out <= rom_array(21913);
		when "0101010110011010" => data_out <= rom_array(21914);
		when "0101010110011011" => data_out <= rom_array(21915);
		when "0101010110011100" => data_out <= rom_array(21916);
		when "0101010110011101" => data_out <= rom_array(21917);
		when "0101010110011110" => data_out <= rom_array(21918);
		when "0101010110011111" => data_out <= rom_array(21919);
		when "0101010110100000" => data_out <= rom_array(21920);
		when "0101010110100001" => data_out <= rom_array(21921);
		when "0101010110100010" => data_out <= rom_array(21922);
		when "0101010110100011" => data_out <= rom_array(21923);
		when "0101010110100100" => data_out <= rom_array(21924);
		when "0101010110100101" => data_out <= rom_array(21925);
		when "0101010110100110" => data_out <= rom_array(21926);
		when "0101010110100111" => data_out <= rom_array(21927);
		when "0101010110101000" => data_out <= rom_array(21928);
		when "0101010110101001" => data_out <= rom_array(21929);
		when "0101010110101010" => data_out <= rom_array(21930);
		when "0101010110101011" => data_out <= rom_array(21931);
		when "0101010110101100" => data_out <= rom_array(21932);
		when "0101010110101101" => data_out <= rom_array(21933);
		when "0101010110101110" => data_out <= rom_array(21934);
		when "0101010110101111" => data_out <= rom_array(21935);
		when "0101010110110000" => data_out <= rom_array(21936);
		when "0101010110110001" => data_out <= rom_array(21937);
		when "0101010110110010" => data_out <= rom_array(21938);
		when "0101010110110011" => data_out <= rom_array(21939);
		when "0101010110110100" => data_out <= rom_array(21940);
		when "0101010110110101" => data_out <= rom_array(21941);
		when "0101010110110110" => data_out <= rom_array(21942);
		when "0101010110110111" => data_out <= rom_array(21943);
		when "0101010110111000" => data_out <= rom_array(21944);
		when "0101010110111001" => data_out <= rom_array(21945);
		when "0101010110111010" => data_out <= rom_array(21946);
		when "0101010110111011" => data_out <= rom_array(21947);
		when "0101010110111100" => data_out <= rom_array(21948);
		when "0101010110111101" => data_out <= rom_array(21949);
		when "0101010110111110" => data_out <= rom_array(21950);
		when "0101010110111111" => data_out <= rom_array(21951);
		when "0101010111000000" => data_out <= rom_array(21952);
		when "0101010111000001" => data_out <= rom_array(21953);
		when "0101010111000010" => data_out <= rom_array(21954);
		when "0101010111000011" => data_out <= rom_array(21955);
		when "0101010111000100" => data_out <= rom_array(21956);
		when "0101010111000101" => data_out <= rom_array(21957);
		when "0101010111000110" => data_out <= rom_array(21958);
		when "0101010111000111" => data_out <= rom_array(21959);
		when "0101010111001000" => data_out <= rom_array(21960);
		when "0101010111001001" => data_out <= rom_array(21961);
		when "0101010111001010" => data_out <= rom_array(21962);
		when "0101010111001011" => data_out <= rom_array(21963);
		when "0101010111001100" => data_out <= rom_array(21964);
		when "0101010111001101" => data_out <= rom_array(21965);
		when "0101010111001110" => data_out <= rom_array(21966);
		when "0101010111001111" => data_out <= rom_array(21967);
		when "0101010111010000" => data_out <= rom_array(21968);
		when "0101010111010001" => data_out <= rom_array(21969);
		when "0101010111010010" => data_out <= rom_array(21970);
		when "0101010111010011" => data_out <= rom_array(21971);
		when "0101010111010100" => data_out <= rom_array(21972);
		when "0101010111010101" => data_out <= rom_array(21973);
		when "0101010111010110" => data_out <= rom_array(21974);
		when "0101010111010111" => data_out <= rom_array(21975);
		when "0101010111011000" => data_out <= rom_array(21976);
		when "0101010111011001" => data_out <= rom_array(21977);
		when "0101010111011010" => data_out <= rom_array(21978);
		when "0101010111011011" => data_out <= rom_array(21979);
		when "0101010111011100" => data_out <= rom_array(21980);
		when "0101010111011101" => data_out <= rom_array(21981);
		when "0101010111011110" => data_out <= rom_array(21982);
		when "0101010111011111" => data_out <= rom_array(21983);
		when "0101010111100000" => data_out <= rom_array(21984);
		when "0101010111100001" => data_out <= rom_array(21985);
		when "0101010111100010" => data_out <= rom_array(21986);
		when "0101010111100011" => data_out <= rom_array(21987);
		when "0101010111100100" => data_out <= rom_array(21988);
		when "0101010111100101" => data_out <= rom_array(21989);
		when "0101010111100110" => data_out <= rom_array(21990);
		when "0101010111100111" => data_out <= rom_array(21991);
		when "0101010111101000" => data_out <= rom_array(21992);
		when "0101010111101001" => data_out <= rom_array(21993);
		when "0101010111101010" => data_out <= rom_array(21994);
		when "0101010111101011" => data_out <= rom_array(21995);
		when "0101010111101100" => data_out <= rom_array(21996);
		when "0101010111101101" => data_out <= rom_array(21997);
		when "0101010111101110" => data_out <= rom_array(21998);
		when "0101010111101111" => data_out <= rom_array(21999);
		when "0101010111110000" => data_out <= rom_array(22000);
		when "0101010111110001" => data_out <= rom_array(22001);
		when "0101010111110010" => data_out <= rom_array(22002);
		when "0101010111110011" => data_out <= rom_array(22003);
		when "0101010111110100" => data_out <= rom_array(22004);
		when "0101010111110101" => data_out <= rom_array(22005);
		when "0101010111110110" => data_out <= rom_array(22006);
		when "0101010111110111" => data_out <= rom_array(22007);
		when "0101010111111000" => data_out <= rom_array(22008);
		when "0101010111111001" => data_out <= rom_array(22009);
		when "0101010111111010" => data_out <= rom_array(22010);
		when "0101010111111011" => data_out <= rom_array(22011);
		when "0101010111111100" => data_out <= rom_array(22012);
		when "0101010111111101" => data_out <= rom_array(22013);
		when "0101010111111110" => data_out <= rom_array(22014);
		when "0101010111111111" => data_out <= rom_array(22015);
		when "0101011000000000" => data_out <= rom_array(22016);
		when "0101011000000001" => data_out <= rom_array(22017);
		when "0101011000000010" => data_out <= rom_array(22018);
		when "0101011000000011" => data_out <= rom_array(22019);
		when "0101011000000100" => data_out <= rom_array(22020);
		when "0101011000000101" => data_out <= rom_array(22021);
		when "0101011000000110" => data_out <= rom_array(22022);
		when "0101011000000111" => data_out <= rom_array(22023);
		when "0101011000001000" => data_out <= rom_array(22024);
		when "0101011000001001" => data_out <= rom_array(22025);
		when "0101011000001010" => data_out <= rom_array(22026);
		when "0101011000001011" => data_out <= rom_array(22027);
		when "0101011000001100" => data_out <= rom_array(22028);
		when "0101011000001101" => data_out <= rom_array(22029);
		when "0101011000001110" => data_out <= rom_array(22030);
		when "0101011000001111" => data_out <= rom_array(22031);
		when "0101011000010000" => data_out <= rom_array(22032);
		when "0101011000010001" => data_out <= rom_array(22033);
		when "0101011000010010" => data_out <= rom_array(22034);
		when "0101011000010011" => data_out <= rom_array(22035);
		when "0101011000010100" => data_out <= rom_array(22036);
		when "0101011000010101" => data_out <= rom_array(22037);
		when "0101011000010110" => data_out <= rom_array(22038);
		when "0101011000010111" => data_out <= rom_array(22039);
		when "0101011000011000" => data_out <= rom_array(22040);
		when "0101011000011001" => data_out <= rom_array(22041);
		when "0101011000011010" => data_out <= rom_array(22042);
		when "0101011000011011" => data_out <= rom_array(22043);
		when "0101011000011100" => data_out <= rom_array(22044);
		when "0101011000011101" => data_out <= rom_array(22045);
		when "0101011000011110" => data_out <= rom_array(22046);
		when "0101011000011111" => data_out <= rom_array(22047);
		when "0101011000100000" => data_out <= rom_array(22048);
		when "0101011000100001" => data_out <= rom_array(22049);
		when "0101011000100010" => data_out <= rom_array(22050);
		when "0101011000100011" => data_out <= rom_array(22051);
		when "0101011000100100" => data_out <= rom_array(22052);
		when "0101011000100101" => data_out <= rom_array(22053);
		when "0101011000100110" => data_out <= rom_array(22054);
		when "0101011000100111" => data_out <= rom_array(22055);
		when "0101011000101000" => data_out <= rom_array(22056);
		when "0101011000101001" => data_out <= rom_array(22057);
		when "0101011000101010" => data_out <= rom_array(22058);
		when "0101011000101011" => data_out <= rom_array(22059);
		when "0101011000101100" => data_out <= rom_array(22060);
		when "0101011000101101" => data_out <= rom_array(22061);
		when "0101011000101110" => data_out <= rom_array(22062);
		when "0101011000101111" => data_out <= rom_array(22063);
		when "0101011000110000" => data_out <= rom_array(22064);
		when "0101011000110001" => data_out <= rom_array(22065);
		when "0101011000110010" => data_out <= rom_array(22066);
		when "0101011000110011" => data_out <= rom_array(22067);
		when "0101011000110100" => data_out <= rom_array(22068);
		when "0101011000110101" => data_out <= rom_array(22069);
		when "0101011000110110" => data_out <= rom_array(22070);
		when "0101011000110111" => data_out <= rom_array(22071);
		when "0101011000111000" => data_out <= rom_array(22072);
		when "0101011000111001" => data_out <= rom_array(22073);
		when "0101011000111010" => data_out <= rom_array(22074);
		when "0101011000111011" => data_out <= rom_array(22075);
		when "0101011000111100" => data_out <= rom_array(22076);
		when "0101011000111101" => data_out <= rom_array(22077);
		when "0101011000111110" => data_out <= rom_array(22078);
		when "0101011000111111" => data_out <= rom_array(22079);
		when "0101011001000000" => data_out <= rom_array(22080);
		when "0101011001000001" => data_out <= rom_array(22081);
		when "0101011001000010" => data_out <= rom_array(22082);
		when "0101011001000011" => data_out <= rom_array(22083);
		when "0101011001000100" => data_out <= rom_array(22084);
		when "0101011001000101" => data_out <= rom_array(22085);
		when "0101011001000110" => data_out <= rom_array(22086);
		when "0101011001000111" => data_out <= rom_array(22087);
		when "0101011001001000" => data_out <= rom_array(22088);
		when "0101011001001001" => data_out <= rom_array(22089);
		when "0101011001001010" => data_out <= rom_array(22090);
		when "0101011001001011" => data_out <= rom_array(22091);
		when "0101011001001100" => data_out <= rom_array(22092);
		when "0101011001001101" => data_out <= rom_array(22093);
		when "0101011001001110" => data_out <= rom_array(22094);
		when "0101011001001111" => data_out <= rom_array(22095);
		when "0101011001010000" => data_out <= rom_array(22096);
		when "0101011001010001" => data_out <= rom_array(22097);
		when "0101011001010010" => data_out <= rom_array(22098);
		when "0101011001010011" => data_out <= rom_array(22099);
		when "0101011001010100" => data_out <= rom_array(22100);
		when "0101011001010101" => data_out <= rom_array(22101);
		when "0101011001010110" => data_out <= rom_array(22102);
		when "0101011001010111" => data_out <= rom_array(22103);
		when "0101011001011000" => data_out <= rom_array(22104);
		when "0101011001011001" => data_out <= rom_array(22105);
		when "0101011001011010" => data_out <= rom_array(22106);
		when "0101011001011011" => data_out <= rom_array(22107);
		when "0101011001011100" => data_out <= rom_array(22108);
		when "0101011001011101" => data_out <= rom_array(22109);
		when "0101011001011110" => data_out <= rom_array(22110);
		when "0101011001011111" => data_out <= rom_array(22111);
		when "0101011001100000" => data_out <= rom_array(22112);
		when "0101011001100001" => data_out <= rom_array(22113);
		when "0101011001100010" => data_out <= rom_array(22114);
		when "0101011001100011" => data_out <= rom_array(22115);
		when "0101011001100100" => data_out <= rom_array(22116);
		when "0101011001100101" => data_out <= rom_array(22117);
		when "0101011001100110" => data_out <= rom_array(22118);
		when "0101011001100111" => data_out <= rom_array(22119);
		when "0101011001101000" => data_out <= rom_array(22120);
		when "0101011001101001" => data_out <= rom_array(22121);
		when "0101011001101010" => data_out <= rom_array(22122);
		when "0101011001101011" => data_out <= rom_array(22123);
		when "0101011001101100" => data_out <= rom_array(22124);
		when "0101011001101101" => data_out <= rom_array(22125);
		when "0101011001101110" => data_out <= rom_array(22126);
		when "0101011001101111" => data_out <= rom_array(22127);
		when "0101011001110000" => data_out <= rom_array(22128);
		when "0101011001110001" => data_out <= rom_array(22129);
		when "0101011001110010" => data_out <= rom_array(22130);
		when "0101011001110011" => data_out <= rom_array(22131);
		when "0101011001110100" => data_out <= rom_array(22132);
		when "0101011001110101" => data_out <= rom_array(22133);
		when "0101011001110110" => data_out <= rom_array(22134);
		when "0101011001110111" => data_out <= rom_array(22135);
		when "0101011001111000" => data_out <= rom_array(22136);
		when "0101011001111001" => data_out <= rom_array(22137);
		when "0101011001111010" => data_out <= rom_array(22138);
		when "0101011001111011" => data_out <= rom_array(22139);
		when "0101011001111100" => data_out <= rom_array(22140);
		when "0101011001111101" => data_out <= rom_array(22141);
		when "0101011001111110" => data_out <= rom_array(22142);
		when "0101011001111111" => data_out <= rom_array(22143);
		when "0101011010000000" => data_out <= rom_array(22144);
		when "0101011010000001" => data_out <= rom_array(22145);
		when "0101011010000010" => data_out <= rom_array(22146);
		when "0101011010000011" => data_out <= rom_array(22147);
		when "0101011010000100" => data_out <= rom_array(22148);
		when "0101011010000101" => data_out <= rom_array(22149);
		when "0101011010000110" => data_out <= rom_array(22150);
		when "0101011010000111" => data_out <= rom_array(22151);
		when "0101011010001000" => data_out <= rom_array(22152);
		when "0101011010001001" => data_out <= rom_array(22153);
		when "0101011010001010" => data_out <= rom_array(22154);
		when "0101011010001011" => data_out <= rom_array(22155);
		when "0101011010001100" => data_out <= rom_array(22156);
		when "0101011010001101" => data_out <= rom_array(22157);
		when "0101011010001110" => data_out <= rom_array(22158);
		when "0101011010001111" => data_out <= rom_array(22159);
		when "0101011010010000" => data_out <= rom_array(22160);
		when "0101011010010001" => data_out <= rom_array(22161);
		when "0101011010010010" => data_out <= rom_array(22162);
		when "0101011010010011" => data_out <= rom_array(22163);
		when "0101011010010100" => data_out <= rom_array(22164);
		when "0101011010010101" => data_out <= rom_array(22165);
		when "0101011010010110" => data_out <= rom_array(22166);
		when "0101011010010111" => data_out <= rom_array(22167);
		when "0101011010011000" => data_out <= rom_array(22168);
		when "0101011010011001" => data_out <= rom_array(22169);
		when "0101011010011010" => data_out <= rom_array(22170);
		when "0101011010011011" => data_out <= rom_array(22171);
		when "0101011010011100" => data_out <= rom_array(22172);
		when "0101011010011101" => data_out <= rom_array(22173);
		when "0101011010011110" => data_out <= rom_array(22174);
		when "0101011010011111" => data_out <= rom_array(22175);
		when "0101011010100000" => data_out <= rom_array(22176);
		when "0101011010100001" => data_out <= rom_array(22177);
		when "0101011010100010" => data_out <= rom_array(22178);
		when "0101011010100011" => data_out <= rom_array(22179);
		when "0101011010100100" => data_out <= rom_array(22180);
		when "0101011010100101" => data_out <= rom_array(22181);
		when "0101011010100110" => data_out <= rom_array(22182);
		when "0101011010100111" => data_out <= rom_array(22183);
		when "0101011010101000" => data_out <= rom_array(22184);
		when "0101011010101001" => data_out <= rom_array(22185);
		when "0101011010101010" => data_out <= rom_array(22186);
		when "0101011010101011" => data_out <= rom_array(22187);
		when "0101011010101100" => data_out <= rom_array(22188);
		when "0101011010101101" => data_out <= rom_array(22189);
		when "0101011010101110" => data_out <= rom_array(22190);
		when "0101011010101111" => data_out <= rom_array(22191);
		when "0101011010110000" => data_out <= rom_array(22192);
		when "0101011010110001" => data_out <= rom_array(22193);
		when "0101011010110010" => data_out <= rom_array(22194);
		when "0101011010110011" => data_out <= rom_array(22195);
		when "0101011010110100" => data_out <= rom_array(22196);
		when "0101011010110101" => data_out <= rom_array(22197);
		when "0101011010110110" => data_out <= rom_array(22198);
		when "0101011010110111" => data_out <= rom_array(22199);
		when "0101011010111000" => data_out <= rom_array(22200);
		when "0101011010111001" => data_out <= rom_array(22201);
		when "0101011010111010" => data_out <= rom_array(22202);
		when "0101011010111011" => data_out <= rom_array(22203);
		when "0101011010111100" => data_out <= rom_array(22204);
		when "0101011010111101" => data_out <= rom_array(22205);
		when "0101011010111110" => data_out <= rom_array(22206);
		when "0101011010111111" => data_out <= rom_array(22207);
		when "0101011011000000" => data_out <= rom_array(22208);
		when "0101011011000001" => data_out <= rom_array(22209);
		when "0101011011000010" => data_out <= rom_array(22210);
		when "0101011011000011" => data_out <= rom_array(22211);
		when "0101011011000100" => data_out <= rom_array(22212);
		when "0101011011000101" => data_out <= rom_array(22213);
		when "0101011011000110" => data_out <= rom_array(22214);
		when "0101011011000111" => data_out <= rom_array(22215);
		when "0101011011001000" => data_out <= rom_array(22216);
		when "0101011011001001" => data_out <= rom_array(22217);
		when "0101011011001010" => data_out <= rom_array(22218);
		when "0101011011001011" => data_out <= rom_array(22219);
		when "0101011011001100" => data_out <= rom_array(22220);
		when "0101011011001101" => data_out <= rom_array(22221);
		when "0101011011001110" => data_out <= rom_array(22222);
		when "0101011011001111" => data_out <= rom_array(22223);
		when "0101011011010000" => data_out <= rom_array(22224);
		when "0101011011010001" => data_out <= rom_array(22225);
		when "0101011011010010" => data_out <= rom_array(22226);
		when "0101011011010011" => data_out <= rom_array(22227);
		when "0101011011010100" => data_out <= rom_array(22228);
		when "0101011011010101" => data_out <= rom_array(22229);
		when "0101011011010110" => data_out <= rom_array(22230);
		when "0101011011010111" => data_out <= rom_array(22231);
		when "0101011011011000" => data_out <= rom_array(22232);
		when "0101011011011001" => data_out <= rom_array(22233);
		when "0101011011011010" => data_out <= rom_array(22234);
		when "0101011011011011" => data_out <= rom_array(22235);
		when "0101011011011100" => data_out <= rom_array(22236);
		when "0101011011011101" => data_out <= rom_array(22237);
		when "0101011011011110" => data_out <= rom_array(22238);
		when "0101011011011111" => data_out <= rom_array(22239);
		when "0101011011100000" => data_out <= rom_array(22240);
		when "0101011011100001" => data_out <= rom_array(22241);
		when "0101011011100010" => data_out <= rom_array(22242);
		when "0101011011100011" => data_out <= rom_array(22243);
		when "0101011011100100" => data_out <= rom_array(22244);
		when "0101011011100101" => data_out <= rom_array(22245);
		when "0101011011100110" => data_out <= rom_array(22246);
		when "0101011011100111" => data_out <= rom_array(22247);
		when "0101011011101000" => data_out <= rom_array(22248);
		when "0101011011101001" => data_out <= rom_array(22249);
		when "0101011011101010" => data_out <= rom_array(22250);
		when "0101011011101011" => data_out <= rom_array(22251);
		when "0101011011101100" => data_out <= rom_array(22252);
		when "0101011011101101" => data_out <= rom_array(22253);
		when "0101011011101110" => data_out <= rom_array(22254);
		when "0101011011101111" => data_out <= rom_array(22255);
		when "0101011011110000" => data_out <= rom_array(22256);
		when "0101011011110001" => data_out <= rom_array(22257);
		when "0101011011110010" => data_out <= rom_array(22258);
		when "0101011011110011" => data_out <= rom_array(22259);
		when "0101011011110100" => data_out <= rom_array(22260);
		when "0101011011110101" => data_out <= rom_array(22261);
		when "0101011011110110" => data_out <= rom_array(22262);
		when "0101011011110111" => data_out <= rom_array(22263);
		when "0101011011111000" => data_out <= rom_array(22264);
		when "0101011011111001" => data_out <= rom_array(22265);
		when "0101011011111010" => data_out <= rom_array(22266);
		when "0101011011111011" => data_out <= rom_array(22267);
		when "0101011011111100" => data_out <= rom_array(22268);
		when "0101011011111101" => data_out <= rom_array(22269);
		when "0101011011111110" => data_out <= rom_array(22270);
		when "0101011011111111" => data_out <= rom_array(22271);
		when "0101011100000000" => data_out <= rom_array(22272);
		when "0101011100000001" => data_out <= rom_array(22273);
		when "0101011100000010" => data_out <= rom_array(22274);
		when "0101011100000011" => data_out <= rom_array(22275);
		when "0101011100000100" => data_out <= rom_array(22276);
		when "0101011100000101" => data_out <= rom_array(22277);
		when "0101011100000110" => data_out <= rom_array(22278);
		when "0101011100000111" => data_out <= rom_array(22279);
		when "0101011100001000" => data_out <= rom_array(22280);
		when "0101011100001001" => data_out <= rom_array(22281);
		when "0101011100001010" => data_out <= rom_array(22282);
		when "0101011100001011" => data_out <= rom_array(22283);
		when "0101011100001100" => data_out <= rom_array(22284);
		when "0101011100001101" => data_out <= rom_array(22285);
		when "0101011100001110" => data_out <= rom_array(22286);
		when "0101011100001111" => data_out <= rom_array(22287);
		when "0101011100010000" => data_out <= rom_array(22288);
		when "0101011100010001" => data_out <= rom_array(22289);
		when "0101011100010010" => data_out <= rom_array(22290);
		when "0101011100010011" => data_out <= rom_array(22291);
		when "0101011100010100" => data_out <= rom_array(22292);
		when "0101011100010101" => data_out <= rom_array(22293);
		when "0101011100010110" => data_out <= rom_array(22294);
		when "0101011100010111" => data_out <= rom_array(22295);
		when "0101011100011000" => data_out <= rom_array(22296);
		when "0101011100011001" => data_out <= rom_array(22297);
		when "0101011100011010" => data_out <= rom_array(22298);
		when "0101011100011011" => data_out <= rom_array(22299);
		when "0101011100011100" => data_out <= rom_array(22300);
		when "0101011100011101" => data_out <= rom_array(22301);
		when "0101011100011110" => data_out <= rom_array(22302);
		when "0101011100011111" => data_out <= rom_array(22303);
		when "0101011100100000" => data_out <= rom_array(22304);
		when "0101011100100001" => data_out <= rom_array(22305);
		when "0101011100100010" => data_out <= rom_array(22306);
		when "0101011100100011" => data_out <= rom_array(22307);
		when "0101011100100100" => data_out <= rom_array(22308);
		when "0101011100100101" => data_out <= rom_array(22309);
		when "0101011100100110" => data_out <= rom_array(22310);
		when "0101011100100111" => data_out <= rom_array(22311);
		when "0101011100101000" => data_out <= rom_array(22312);
		when "0101011100101001" => data_out <= rom_array(22313);
		when "0101011100101010" => data_out <= rom_array(22314);
		when "0101011100101011" => data_out <= rom_array(22315);
		when "0101011100101100" => data_out <= rom_array(22316);
		when "0101011100101101" => data_out <= rom_array(22317);
		when "0101011100101110" => data_out <= rom_array(22318);
		when "0101011100101111" => data_out <= rom_array(22319);
		when "0101011100110000" => data_out <= rom_array(22320);
		when "0101011100110001" => data_out <= rom_array(22321);
		when "0101011100110010" => data_out <= rom_array(22322);
		when "0101011100110011" => data_out <= rom_array(22323);
		when "0101011100110100" => data_out <= rom_array(22324);
		when "0101011100110101" => data_out <= rom_array(22325);
		when "0101011100110110" => data_out <= rom_array(22326);
		when "0101011100110111" => data_out <= rom_array(22327);
		when "0101011100111000" => data_out <= rom_array(22328);
		when "0101011100111001" => data_out <= rom_array(22329);
		when "0101011100111010" => data_out <= rom_array(22330);
		when "0101011100111011" => data_out <= rom_array(22331);
		when "0101011100111100" => data_out <= rom_array(22332);
		when "0101011100111101" => data_out <= rom_array(22333);
		when "0101011100111110" => data_out <= rom_array(22334);
		when "0101011100111111" => data_out <= rom_array(22335);
		when "0101011101000000" => data_out <= rom_array(22336);
		when "0101011101000001" => data_out <= rom_array(22337);
		when "0101011101000010" => data_out <= rom_array(22338);
		when "0101011101000011" => data_out <= rom_array(22339);
		when "0101011101000100" => data_out <= rom_array(22340);
		when "0101011101000101" => data_out <= rom_array(22341);
		when "0101011101000110" => data_out <= rom_array(22342);
		when "0101011101000111" => data_out <= rom_array(22343);
		when "0101011101001000" => data_out <= rom_array(22344);
		when "0101011101001001" => data_out <= rom_array(22345);
		when "0101011101001010" => data_out <= rom_array(22346);
		when "0101011101001011" => data_out <= rom_array(22347);
		when "0101011101001100" => data_out <= rom_array(22348);
		when "0101011101001101" => data_out <= rom_array(22349);
		when "0101011101001110" => data_out <= rom_array(22350);
		when "0101011101001111" => data_out <= rom_array(22351);
		when "0101011101010000" => data_out <= rom_array(22352);
		when "0101011101010001" => data_out <= rom_array(22353);
		when "0101011101010010" => data_out <= rom_array(22354);
		when "0101011101010011" => data_out <= rom_array(22355);
		when "0101011101010100" => data_out <= rom_array(22356);
		when "0101011101010101" => data_out <= rom_array(22357);
		when "0101011101010110" => data_out <= rom_array(22358);
		when "0101011101010111" => data_out <= rom_array(22359);
		when "0101011101011000" => data_out <= rom_array(22360);
		when "0101011101011001" => data_out <= rom_array(22361);
		when "0101011101011010" => data_out <= rom_array(22362);
		when "0101011101011011" => data_out <= rom_array(22363);
		when "0101011101011100" => data_out <= rom_array(22364);
		when "0101011101011101" => data_out <= rom_array(22365);
		when "0101011101011110" => data_out <= rom_array(22366);
		when "0101011101011111" => data_out <= rom_array(22367);
		when "0101011101100000" => data_out <= rom_array(22368);
		when "0101011101100001" => data_out <= rom_array(22369);
		when "0101011101100010" => data_out <= rom_array(22370);
		when "0101011101100011" => data_out <= rom_array(22371);
		when "0101011101100100" => data_out <= rom_array(22372);
		when "0101011101100101" => data_out <= rom_array(22373);
		when "0101011101100110" => data_out <= rom_array(22374);
		when "0101011101100111" => data_out <= rom_array(22375);
		when "0101011101101000" => data_out <= rom_array(22376);
		when "0101011101101001" => data_out <= rom_array(22377);
		when "0101011101101010" => data_out <= rom_array(22378);
		when "0101011101101011" => data_out <= rom_array(22379);
		when "0101011101101100" => data_out <= rom_array(22380);
		when "0101011101101101" => data_out <= rom_array(22381);
		when "0101011101101110" => data_out <= rom_array(22382);
		when "0101011101101111" => data_out <= rom_array(22383);
		when "0101011101110000" => data_out <= rom_array(22384);
		when "0101011101110001" => data_out <= rom_array(22385);
		when "0101011101110010" => data_out <= rom_array(22386);
		when "0101011101110011" => data_out <= rom_array(22387);
		when "0101011101110100" => data_out <= rom_array(22388);
		when "0101011101110101" => data_out <= rom_array(22389);
		when "0101011101110110" => data_out <= rom_array(22390);
		when "0101011101110111" => data_out <= rom_array(22391);
		when "0101011101111000" => data_out <= rom_array(22392);
		when "0101011101111001" => data_out <= rom_array(22393);
		when "0101011101111010" => data_out <= rom_array(22394);
		when "0101011101111011" => data_out <= rom_array(22395);
		when "0101011101111100" => data_out <= rom_array(22396);
		when "0101011101111101" => data_out <= rom_array(22397);
		when "0101011101111110" => data_out <= rom_array(22398);
		when "0101011101111111" => data_out <= rom_array(22399);
		when "0101011110000000" => data_out <= rom_array(22400);
		when "0101011110000001" => data_out <= rom_array(22401);
		when "0101011110000010" => data_out <= rom_array(22402);
		when "0101011110000011" => data_out <= rom_array(22403);
		when "0101011110000100" => data_out <= rom_array(22404);
		when "0101011110000101" => data_out <= rom_array(22405);
		when "0101011110000110" => data_out <= rom_array(22406);
		when "0101011110000111" => data_out <= rom_array(22407);
		when "0101011110001000" => data_out <= rom_array(22408);
		when "0101011110001001" => data_out <= rom_array(22409);
		when "0101011110001010" => data_out <= rom_array(22410);
		when "0101011110001011" => data_out <= rom_array(22411);
		when "0101011110001100" => data_out <= rom_array(22412);
		when "0101011110001101" => data_out <= rom_array(22413);
		when "0101011110001110" => data_out <= rom_array(22414);
		when "0101011110001111" => data_out <= rom_array(22415);
		when "0101011110010000" => data_out <= rom_array(22416);
		when "0101011110010001" => data_out <= rom_array(22417);
		when "0101011110010010" => data_out <= rom_array(22418);
		when "0101011110010011" => data_out <= rom_array(22419);
		when "0101011110010100" => data_out <= rom_array(22420);
		when "0101011110010101" => data_out <= rom_array(22421);
		when "0101011110010110" => data_out <= rom_array(22422);
		when "0101011110010111" => data_out <= rom_array(22423);
		when "0101011110011000" => data_out <= rom_array(22424);
		when "0101011110011001" => data_out <= rom_array(22425);
		when "0101011110011010" => data_out <= rom_array(22426);
		when "0101011110011011" => data_out <= rom_array(22427);
		when "0101011110011100" => data_out <= rom_array(22428);
		when "0101011110011101" => data_out <= rom_array(22429);
		when "0101011110011110" => data_out <= rom_array(22430);
		when "0101011110011111" => data_out <= rom_array(22431);
		when "0101011110100000" => data_out <= rom_array(22432);
		when "0101011110100001" => data_out <= rom_array(22433);
		when "0101011110100010" => data_out <= rom_array(22434);
		when "0101011110100011" => data_out <= rom_array(22435);
		when "0101011110100100" => data_out <= rom_array(22436);
		when "0101011110100101" => data_out <= rom_array(22437);
		when "0101011110100110" => data_out <= rom_array(22438);
		when "0101011110100111" => data_out <= rom_array(22439);
		when "0101011110101000" => data_out <= rom_array(22440);
		when "0101011110101001" => data_out <= rom_array(22441);
		when "0101011110101010" => data_out <= rom_array(22442);
		when "0101011110101011" => data_out <= rom_array(22443);
		when "0101011110101100" => data_out <= rom_array(22444);
		when "0101011110101101" => data_out <= rom_array(22445);
		when "0101011110101110" => data_out <= rom_array(22446);
		when "0101011110101111" => data_out <= rom_array(22447);
		when "0101011110110000" => data_out <= rom_array(22448);
		when "0101011110110001" => data_out <= rom_array(22449);
		when "0101011110110010" => data_out <= rom_array(22450);
		when "0101011110110011" => data_out <= rom_array(22451);
		when "0101011110110100" => data_out <= rom_array(22452);
		when "0101011110110101" => data_out <= rom_array(22453);
		when "0101011110110110" => data_out <= rom_array(22454);
		when "0101011110110111" => data_out <= rom_array(22455);
		when "0101011110111000" => data_out <= rom_array(22456);
		when "0101011110111001" => data_out <= rom_array(22457);
		when "0101011110111010" => data_out <= rom_array(22458);
		when "0101011110111011" => data_out <= rom_array(22459);
		when "0101011110111100" => data_out <= rom_array(22460);
		when "0101011110111101" => data_out <= rom_array(22461);
		when "0101011110111110" => data_out <= rom_array(22462);
		when "0101011110111111" => data_out <= rom_array(22463);
		when "0101011111000000" => data_out <= rom_array(22464);
		when "0101011111000001" => data_out <= rom_array(22465);
		when "0101011111000010" => data_out <= rom_array(22466);
		when "0101011111000011" => data_out <= rom_array(22467);
		when "0101011111000100" => data_out <= rom_array(22468);
		when "0101011111000101" => data_out <= rom_array(22469);
		when "0101011111000110" => data_out <= rom_array(22470);
		when "0101011111000111" => data_out <= rom_array(22471);
		when "0101011111001000" => data_out <= rom_array(22472);
		when "0101011111001001" => data_out <= rom_array(22473);
		when "0101011111001010" => data_out <= rom_array(22474);
		when "0101011111001011" => data_out <= rom_array(22475);
		when "0101011111001100" => data_out <= rom_array(22476);
		when "0101011111001101" => data_out <= rom_array(22477);
		when "0101011111001110" => data_out <= rom_array(22478);
		when "0101011111001111" => data_out <= rom_array(22479);
		when "0101011111010000" => data_out <= rom_array(22480);
		when "0101011111010001" => data_out <= rom_array(22481);
		when "0101011111010010" => data_out <= rom_array(22482);
		when "0101011111010011" => data_out <= rom_array(22483);
		when "0101011111010100" => data_out <= rom_array(22484);
		when "0101011111010101" => data_out <= rom_array(22485);
		when "0101011111010110" => data_out <= rom_array(22486);
		when "0101011111010111" => data_out <= rom_array(22487);
		when "0101011111011000" => data_out <= rom_array(22488);
		when "0101011111011001" => data_out <= rom_array(22489);
		when "0101011111011010" => data_out <= rom_array(22490);
		when "0101011111011011" => data_out <= rom_array(22491);
		when "0101011111011100" => data_out <= rom_array(22492);
		when "0101011111011101" => data_out <= rom_array(22493);
		when "0101011111011110" => data_out <= rom_array(22494);
		when "0101011111011111" => data_out <= rom_array(22495);
		when "0101011111100000" => data_out <= rom_array(22496);
		when "0101011111100001" => data_out <= rom_array(22497);
		when "0101011111100010" => data_out <= rom_array(22498);
		when "0101011111100011" => data_out <= rom_array(22499);
		when "0101011111100100" => data_out <= rom_array(22500);
		when "0101011111100101" => data_out <= rom_array(22501);
		when "0101011111100110" => data_out <= rom_array(22502);
		when "0101011111100111" => data_out <= rom_array(22503);
		when "0101011111101000" => data_out <= rom_array(22504);
		when "0101011111101001" => data_out <= rom_array(22505);
		when "0101011111101010" => data_out <= rom_array(22506);
		when "0101011111101011" => data_out <= rom_array(22507);
		when "0101011111101100" => data_out <= rom_array(22508);
		when "0101011111101101" => data_out <= rom_array(22509);
		when "0101011111101110" => data_out <= rom_array(22510);
		when "0101011111101111" => data_out <= rom_array(22511);
		when "0101011111110000" => data_out <= rom_array(22512);
		when "0101011111110001" => data_out <= rom_array(22513);
		when "0101011111110010" => data_out <= rom_array(22514);
		when "0101011111110011" => data_out <= rom_array(22515);
		when "0101011111110100" => data_out <= rom_array(22516);
		when "0101011111110101" => data_out <= rom_array(22517);
		when "0101011111110110" => data_out <= rom_array(22518);
		when "0101011111110111" => data_out <= rom_array(22519);
		when "0101011111111000" => data_out <= rom_array(22520);
		when "0101011111111001" => data_out <= rom_array(22521);
		when "0101011111111010" => data_out <= rom_array(22522);
		when "0101011111111011" => data_out <= rom_array(22523);
		when "0101011111111100" => data_out <= rom_array(22524);
		when "0101011111111101" => data_out <= rom_array(22525);
		when "0101011111111110" => data_out <= rom_array(22526);
		when "0101011111111111" => data_out <= rom_array(22527);
		when "0101100000000000" => data_out <= rom_array(22528);
		when "0101100000000001" => data_out <= rom_array(22529);
		when "0101100000000010" => data_out <= rom_array(22530);
		when "0101100000000011" => data_out <= rom_array(22531);
		when "0101100000000100" => data_out <= rom_array(22532);
		when "0101100000000101" => data_out <= rom_array(22533);
		when "0101100000000110" => data_out <= rom_array(22534);
		when "0101100000000111" => data_out <= rom_array(22535);
		when "0101100000001000" => data_out <= rom_array(22536);
		when "0101100000001001" => data_out <= rom_array(22537);
		when "0101100000001010" => data_out <= rom_array(22538);
		when "0101100000001011" => data_out <= rom_array(22539);
		when "0101100000001100" => data_out <= rom_array(22540);
		when "0101100000001101" => data_out <= rom_array(22541);
		when "0101100000001110" => data_out <= rom_array(22542);
		when "0101100000001111" => data_out <= rom_array(22543);
		when "0101100000010000" => data_out <= rom_array(22544);
		when "0101100000010001" => data_out <= rom_array(22545);
		when "0101100000010010" => data_out <= rom_array(22546);
		when "0101100000010011" => data_out <= rom_array(22547);
		when "0101100000010100" => data_out <= rom_array(22548);
		when "0101100000010101" => data_out <= rom_array(22549);
		when "0101100000010110" => data_out <= rom_array(22550);
		when "0101100000010111" => data_out <= rom_array(22551);
		when "0101100000011000" => data_out <= rom_array(22552);
		when "0101100000011001" => data_out <= rom_array(22553);
		when "0101100000011010" => data_out <= rom_array(22554);
		when "0101100000011011" => data_out <= rom_array(22555);
		when "0101100000011100" => data_out <= rom_array(22556);
		when "0101100000011101" => data_out <= rom_array(22557);
		when "0101100000011110" => data_out <= rom_array(22558);
		when "0101100000011111" => data_out <= rom_array(22559);
		when "0101100000100000" => data_out <= rom_array(22560);
		when "0101100000100001" => data_out <= rom_array(22561);
		when "0101100000100010" => data_out <= rom_array(22562);
		when "0101100000100011" => data_out <= rom_array(22563);
		when "0101100000100100" => data_out <= rom_array(22564);
		when "0101100000100101" => data_out <= rom_array(22565);
		when "0101100000100110" => data_out <= rom_array(22566);
		when "0101100000100111" => data_out <= rom_array(22567);
		when "0101100000101000" => data_out <= rom_array(22568);
		when "0101100000101001" => data_out <= rom_array(22569);
		when "0101100000101010" => data_out <= rom_array(22570);
		when "0101100000101011" => data_out <= rom_array(22571);
		when "0101100000101100" => data_out <= rom_array(22572);
		when "0101100000101101" => data_out <= rom_array(22573);
		when "0101100000101110" => data_out <= rom_array(22574);
		when "0101100000101111" => data_out <= rom_array(22575);
		when "0101100000110000" => data_out <= rom_array(22576);
		when "0101100000110001" => data_out <= rom_array(22577);
		when "0101100000110010" => data_out <= rom_array(22578);
		when "0101100000110011" => data_out <= rom_array(22579);
		when "0101100000110100" => data_out <= rom_array(22580);
		when "0101100000110101" => data_out <= rom_array(22581);
		when "0101100000110110" => data_out <= rom_array(22582);
		when "0101100000110111" => data_out <= rom_array(22583);
		when "0101100000111000" => data_out <= rom_array(22584);
		when "0101100000111001" => data_out <= rom_array(22585);
		when "0101100000111010" => data_out <= rom_array(22586);
		when "0101100000111011" => data_out <= rom_array(22587);
		when "0101100000111100" => data_out <= rom_array(22588);
		when "0101100000111101" => data_out <= rom_array(22589);
		when "0101100000111110" => data_out <= rom_array(22590);
		when "0101100000111111" => data_out <= rom_array(22591);
		when "0101100001000000" => data_out <= rom_array(22592);
		when "0101100001000001" => data_out <= rom_array(22593);
		when "0101100001000010" => data_out <= rom_array(22594);
		when "0101100001000011" => data_out <= rom_array(22595);
		when "0101100001000100" => data_out <= rom_array(22596);
		when "0101100001000101" => data_out <= rom_array(22597);
		when "0101100001000110" => data_out <= rom_array(22598);
		when "0101100001000111" => data_out <= rom_array(22599);
		when "0101100001001000" => data_out <= rom_array(22600);
		when "0101100001001001" => data_out <= rom_array(22601);
		when "0101100001001010" => data_out <= rom_array(22602);
		when "0101100001001011" => data_out <= rom_array(22603);
		when "0101100001001100" => data_out <= rom_array(22604);
		when "0101100001001101" => data_out <= rom_array(22605);
		when "0101100001001110" => data_out <= rom_array(22606);
		when "0101100001001111" => data_out <= rom_array(22607);
		when "0101100001010000" => data_out <= rom_array(22608);
		when "0101100001010001" => data_out <= rom_array(22609);
		when "0101100001010010" => data_out <= rom_array(22610);
		when "0101100001010011" => data_out <= rom_array(22611);
		when "0101100001010100" => data_out <= rom_array(22612);
		when "0101100001010101" => data_out <= rom_array(22613);
		when "0101100001010110" => data_out <= rom_array(22614);
		when "0101100001010111" => data_out <= rom_array(22615);
		when "0101100001011000" => data_out <= rom_array(22616);
		when "0101100001011001" => data_out <= rom_array(22617);
		when "0101100001011010" => data_out <= rom_array(22618);
		when "0101100001011011" => data_out <= rom_array(22619);
		when "0101100001011100" => data_out <= rom_array(22620);
		when "0101100001011101" => data_out <= rom_array(22621);
		when "0101100001011110" => data_out <= rom_array(22622);
		when "0101100001011111" => data_out <= rom_array(22623);
		when "0101100001100000" => data_out <= rom_array(22624);
		when "0101100001100001" => data_out <= rom_array(22625);
		when "0101100001100010" => data_out <= rom_array(22626);
		when "0101100001100011" => data_out <= rom_array(22627);
		when "0101100001100100" => data_out <= rom_array(22628);
		when "0101100001100101" => data_out <= rom_array(22629);
		when "0101100001100110" => data_out <= rom_array(22630);
		when "0101100001100111" => data_out <= rom_array(22631);
		when "0101100001101000" => data_out <= rom_array(22632);
		when "0101100001101001" => data_out <= rom_array(22633);
		when "0101100001101010" => data_out <= rom_array(22634);
		when "0101100001101011" => data_out <= rom_array(22635);
		when "0101100001101100" => data_out <= rom_array(22636);
		when "0101100001101101" => data_out <= rom_array(22637);
		when "0101100001101110" => data_out <= rom_array(22638);
		when "0101100001101111" => data_out <= rom_array(22639);
		when "0101100001110000" => data_out <= rom_array(22640);
		when "0101100001110001" => data_out <= rom_array(22641);
		when "0101100001110010" => data_out <= rom_array(22642);
		when "0101100001110011" => data_out <= rom_array(22643);
		when "0101100001110100" => data_out <= rom_array(22644);
		when "0101100001110101" => data_out <= rom_array(22645);
		when "0101100001110110" => data_out <= rom_array(22646);
		when "0101100001110111" => data_out <= rom_array(22647);
		when "0101100001111000" => data_out <= rom_array(22648);
		when "0101100001111001" => data_out <= rom_array(22649);
		when "0101100001111010" => data_out <= rom_array(22650);
		when "0101100001111011" => data_out <= rom_array(22651);
		when "0101100001111100" => data_out <= rom_array(22652);
		when "0101100001111101" => data_out <= rom_array(22653);
		when "0101100001111110" => data_out <= rom_array(22654);
		when "0101100001111111" => data_out <= rom_array(22655);
		when "0101100010000000" => data_out <= rom_array(22656);
		when "0101100010000001" => data_out <= rom_array(22657);
		when "0101100010000010" => data_out <= rom_array(22658);
		when "0101100010000011" => data_out <= rom_array(22659);
		when "0101100010000100" => data_out <= rom_array(22660);
		when "0101100010000101" => data_out <= rom_array(22661);
		when "0101100010000110" => data_out <= rom_array(22662);
		when "0101100010000111" => data_out <= rom_array(22663);
		when "0101100010001000" => data_out <= rom_array(22664);
		when "0101100010001001" => data_out <= rom_array(22665);
		when "0101100010001010" => data_out <= rom_array(22666);
		when "0101100010001011" => data_out <= rom_array(22667);
		when "0101100010001100" => data_out <= rom_array(22668);
		when "0101100010001101" => data_out <= rom_array(22669);
		when "0101100010001110" => data_out <= rom_array(22670);
		when "0101100010001111" => data_out <= rom_array(22671);
		when "0101100010010000" => data_out <= rom_array(22672);
		when "0101100010010001" => data_out <= rom_array(22673);
		when "0101100010010010" => data_out <= rom_array(22674);
		when "0101100010010011" => data_out <= rom_array(22675);
		when "0101100010010100" => data_out <= rom_array(22676);
		when "0101100010010101" => data_out <= rom_array(22677);
		when "0101100010010110" => data_out <= rom_array(22678);
		when "0101100010010111" => data_out <= rom_array(22679);
		when "0101100010011000" => data_out <= rom_array(22680);
		when "0101100010011001" => data_out <= rom_array(22681);
		when "0101100010011010" => data_out <= rom_array(22682);
		when "0101100010011011" => data_out <= rom_array(22683);
		when "0101100010011100" => data_out <= rom_array(22684);
		when "0101100010011101" => data_out <= rom_array(22685);
		when "0101100010011110" => data_out <= rom_array(22686);
		when "0101100010011111" => data_out <= rom_array(22687);
		when "0101100010100000" => data_out <= rom_array(22688);
		when "0101100010100001" => data_out <= rom_array(22689);
		when "0101100010100010" => data_out <= rom_array(22690);
		when "0101100010100011" => data_out <= rom_array(22691);
		when "0101100010100100" => data_out <= rom_array(22692);
		when "0101100010100101" => data_out <= rom_array(22693);
		when "0101100010100110" => data_out <= rom_array(22694);
		when "0101100010100111" => data_out <= rom_array(22695);
		when "0101100010101000" => data_out <= rom_array(22696);
		when "0101100010101001" => data_out <= rom_array(22697);
		when "0101100010101010" => data_out <= rom_array(22698);
		when "0101100010101011" => data_out <= rom_array(22699);
		when "0101100010101100" => data_out <= rom_array(22700);
		when "0101100010101101" => data_out <= rom_array(22701);
		when "0101100010101110" => data_out <= rom_array(22702);
		when "0101100010101111" => data_out <= rom_array(22703);
		when "0101100010110000" => data_out <= rom_array(22704);
		when "0101100010110001" => data_out <= rom_array(22705);
		when "0101100010110010" => data_out <= rom_array(22706);
		when "0101100010110011" => data_out <= rom_array(22707);
		when "0101100010110100" => data_out <= rom_array(22708);
		when "0101100010110101" => data_out <= rom_array(22709);
		when "0101100010110110" => data_out <= rom_array(22710);
		when "0101100010110111" => data_out <= rom_array(22711);
		when "0101100010111000" => data_out <= rom_array(22712);
		when "0101100010111001" => data_out <= rom_array(22713);
		when "0101100010111010" => data_out <= rom_array(22714);
		when "0101100010111011" => data_out <= rom_array(22715);
		when "0101100010111100" => data_out <= rom_array(22716);
		when "0101100010111101" => data_out <= rom_array(22717);
		when "0101100010111110" => data_out <= rom_array(22718);
		when "0101100010111111" => data_out <= rom_array(22719);
		when "0101100011000000" => data_out <= rom_array(22720);
		when "0101100011000001" => data_out <= rom_array(22721);
		when "0101100011000010" => data_out <= rom_array(22722);
		when "0101100011000011" => data_out <= rom_array(22723);
		when "0101100011000100" => data_out <= rom_array(22724);
		when "0101100011000101" => data_out <= rom_array(22725);
		when "0101100011000110" => data_out <= rom_array(22726);
		when "0101100011000111" => data_out <= rom_array(22727);
		when "0101100011001000" => data_out <= rom_array(22728);
		when "0101100011001001" => data_out <= rom_array(22729);
		when "0101100011001010" => data_out <= rom_array(22730);
		when "0101100011001011" => data_out <= rom_array(22731);
		when "0101100011001100" => data_out <= rom_array(22732);
		when "0101100011001101" => data_out <= rom_array(22733);
		when "0101100011001110" => data_out <= rom_array(22734);
		when "0101100011001111" => data_out <= rom_array(22735);
		when "0101100011010000" => data_out <= rom_array(22736);
		when "0101100011010001" => data_out <= rom_array(22737);
		when "0101100011010010" => data_out <= rom_array(22738);
		when "0101100011010011" => data_out <= rom_array(22739);
		when "0101100011010100" => data_out <= rom_array(22740);
		when "0101100011010101" => data_out <= rom_array(22741);
		when "0101100011010110" => data_out <= rom_array(22742);
		when "0101100011010111" => data_out <= rom_array(22743);
		when "0101100011011000" => data_out <= rom_array(22744);
		when "0101100011011001" => data_out <= rom_array(22745);
		when "0101100011011010" => data_out <= rom_array(22746);
		when "0101100011011011" => data_out <= rom_array(22747);
		when "0101100011011100" => data_out <= rom_array(22748);
		when "0101100011011101" => data_out <= rom_array(22749);
		when "0101100011011110" => data_out <= rom_array(22750);
		when "0101100011011111" => data_out <= rom_array(22751);
		when "0101100011100000" => data_out <= rom_array(22752);
		when "0101100011100001" => data_out <= rom_array(22753);
		when "0101100011100010" => data_out <= rom_array(22754);
		when "0101100011100011" => data_out <= rom_array(22755);
		when "0101100011100100" => data_out <= rom_array(22756);
		when "0101100011100101" => data_out <= rom_array(22757);
		when "0101100011100110" => data_out <= rom_array(22758);
		when "0101100011100111" => data_out <= rom_array(22759);
		when "0101100011101000" => data_out <= rom_array(22760);
		when "0101100011101001" => data_out <= rom_array(22761);
		when "0101100011101010" => data_out <= rom_array(22762);
		when "0101100011101011" => data_out <= rom_array(22763);
		when "0101100011101100" => data_out <= rom_array(22764);
		when "0101100011101101" => data_out <= rom_array(22765);
		when "0101100011101110" => data_out <= rom_array(22766);
		when "0101100011101111" => data_out <= rom_array(22767);
		when "0101100011110000" => data_out <= rom_array(22768);
		when "0101100011110001" => data_out <= rom_array(22769);
		when "0101100011110010" => data_out <= rom_array(22770);
		when "0101100011110011" => data_out <= rom_array(22771);
		when "0101100011110100" => data_out <= rom_array(22772);
		when "0101100011110101" => data_out <= rom_array(22773);
		when "0101100011110110" => data_out <= rom_array(22774);
		when "0101100011110111" => data_out <= rom_array(22775);
		when "0101100011111000" => data_out <= rom_array(22776);
		when "0101100011111001" => data_out <= rom_array(22777);
		when "0101100011111010" => data_out <= rom_array(22778);
		when "0101100011111011" => data_out <= rom_array(22779);
		when "0101100011111100" => data_out <= rom_array(22780);
		when "0101100011111101" => data_out <= rom_array(22781);
		when "0101100011111110" => data_out <= rom_array(22782);
		when "0101100011111111" => data_out <= rom_array(22783);
		when "0101100100000000" => data_out <= rom_array(22784);
		when "0101100100000001" => data_out <= rom_array(22785);
		when "0101100100000010" => data_out <= rom_array(22786);
		when "0101100100000011" => data_out <= rom_array(22787);
		when "0101100100000100" => data_out <= rom_array(22788);
		when "0101100100000101" => data_out <= rom_array(22789);
		when "0101100100000110" => data_out <= rom_array(22790);
		when "0101100100000111" => data_out <= rom_array(22791);
		when "0101100100001000" => data_out <= rom_array(22792);
		when "0101100100001001" => data_out <= rom_array(22793);
		when "0101100100001010" => data_out <= rom_array(22794);
		when "0101100100001011" => data_out <= rom_array(22795);
		when "0101100100001100" => data_out <= rom_array(22796);
		when "0101100100001101" => data_out <= rom_array(22797);
		when "0101100100001110" => data_out <= rom_array(22798);
		when "0101100100001111" => data_out <= rom_array(22799);
		when "0101100100010000" => data_out <= rom_array(22800);
		when "0101100100010001" => data_out <= rom_array(22801);
		when "0101100100010010" => data_out <= rom_array(22802);
		when "0101100100010011" => data_out <= rom_array(22803);
		when "0101100100010100" => data_out <= rom_array(22804);
		when "0101100100010101" => data_out <= rom_array(22805);
		when "0101100100010110" => data_out <= rom_array(22806);
		when "0101100100010111" => data_out <= rom_array(22807);
		when "0101100100011000" => data_out <= rom_array(22808);
		when "0101100100011001" => data_out <= rom_array(22809);
		when "0101100100011010" => data_out <= rom_array(22810);
		when "0101100100011011" => data_out <= rom_array(22811);
		when "0101100100011100" => data_out <= rom_array(22812);
		when "0101100100011101" => data_out <= rom_array(22813);
		when "0101100100011110" => data_out <= rom_array(22814);
		when "0101100100011111" => data_out <= rom_array(22815);
		when "0101100100100000" => data_out <= rom_array(22816);
		when "0101100100100001" => data_out <= rom_array(22817);
		when "0101100100100010" => data_out <= rom_array(22818);
		when "0101100100100011" => data_out <= rom_array(22819);
		when "0101100100100100" => data_out <= rom_array(22820);
		when "0101100100100101" => data_out <= rom_array(22821);
		when "0101100100100110" => data_out <= rom_array(22822);
		when "0101100100100111" => data_out <= rom_array(22823);
		when "0101100100101000" => data_out <= rom_array(22824);
		when "0101100100101001" => data_out <= rom_array(22825);
		when "0101100100101010" => data_out <= rom_array(22826);
		when "0101100100101011" => data_out <= rom_array(22827);
		when "0101100100101100" => data_out <= rom_array(22828);
		when "0101100100101101" => data_out <= rom_array(22829);
		when "0101100100101110" => data_out <= rom_array(22830);
		when "0101100100101111" => data_out <= rom_array(22831);
		when "0101100100110000" => data_out <= rom_array(22832);
		when "0101100100110001" => data_out <= rom_array(22833);
		when "0101100100110010" => data_out <= rom_array(22834);
		when "0101100100110011" => data_out <= rom_array(22835);
		when "0101100100110100" => data_out <= rom_array(22836);
		when "0101100100110101" => data_out <= rom_array(22837);
		when "0101100100110110" => data_out <= rom_array(22838);
		when "0101100100110111" => data_out <= rom_array(22839);
		when "0101100100111000" => data_out <= rom_array(22840);
		when "0101100100111001" => data_out <= rom_array(22841);
		when "0101100100111010" => data_out <= rom_array(22842);
		when "0101100100111011" => data_out <= rom_array(22843);
		when "0101100100111100" => data_out <= rom_array(22844);
		when "0101100100111101" => data_out <= rom_array(22845);
		when "0101100100111110" => data_out <= rom_array(22846);
		when "0101100100111111" => data_out <= rom_array(22847);
		when "0101100101000000" => data_out <= rom_array(22848);
		when "0101100101000001" => data_out <= rom_array(22849);
		when "0101100101000010" => data_out <= rom_array(22850);
		when "0101100101000011" => data_out <= rom_array(22851);
		when "0101100101000100" => data_out <= rom_array(22852);
		when "0101100101000101" => data_out <= rom_array(22853);
		when "0101100101000110" => data_out <= rom_array(22854);
		when "0101100101000111" => data_out <= rom_array(22855);
		when "0101100101001000" => data_out <= rom_array(22856);
		when "0101100101001001" => data_out <= rom_array(22857);
		when "0101100101001010" => data_out <= rom_array(22858);
		when "0101100101001011" => data_out <= rom_array(22859);
		when "0101100101001100" => data_out <= rom_array(22860);
		when "0101100101001101" => data_out <= rom_array(22861);
		when "0101100101001110" => data_out <= rom_array(22862);
		when "0101100101001111" => data_out <= rom_array(22863);
		when "0101100101010000" => data_out <= rom_array(22864);
		when "0101100101010001" => data_out <= rom_array(22865);
		when "0101100101010010" => data_out <= rom_array(22866);
		when "0101100101010011" => data_out <= rom_array(22867);
		when "0101100101010100" => data_out <= rom_array(22868);
		when "0101100101010101" => data_out <= rom_array(22869);
		when "0101100101010110" => data_out <= rom_array(22870);
		when "0101100101010111" => data_out <= rom_array(22871);
		when "0101100101011000" => data_out <= rom_array(22872);
		when "0101100101011001" => data_out <= rom_array(22873);
		when "0101100101011010" => data_out <= rom_array(22874);
		when "0101100101011011" => data_out <= rom_array(22875);
		when "0101100101011100" => data_out <= rom_array(22876);
		when "0101100101011101" => data_out <= rom_array(22877);
		when "0101100101011110" => data_out <= rom_array(22878);
		when "0101100101011111" => data_out <= rom_array(22879);
		when "0101100101100000" => data_out <= rom_array(22880);
		when "0101100101100001" => data_out <= rom_array(22881);
		when "0101100101100010" => data_out <= rom_array(22882);
		when "0101100101100011" => data_out <= rom_array(22883);
		when "0101100101100100" => data_out <= rom_array(22884);
		when "0101100101100101" => data_out <= rom_array(22885);
		when "0101100101100110" => data_out <= rom_array(22886);
		when "0101100101100111" => data_out <= rom_array(22887);
		when "0101100101101000" => data_out <= rom_array(22888);
		when "0101100101101001" => data_out <= rom_array(22889);
		when "0101100101101010" => data_out <= rom_array(22890);
		when "0101100101101011" => data_out <= rom_array(22891);
		when "0101100101101100" => data_out <= rom_array(22892);
		when "0101100101101101" => data_out <= rom_array(22893);
		when "0101100101101110" => data_out <= rom_array(22894);
		when "0101100101101111" => data_out <= rom_array(22895);
		when "0101100101110000" => data_out <= rom_array(22896);
		when "0101100101110001" => data_out <= rom_array(22897);
		when "0101100101110010" => data_out <= rom_array(22898);
		when "0101100101110011" => data_out <= rom_array(22899);
		when "0101100101110100" => data_out <= rom_array(22900);
		when "0101100101110101" => data_out <= rom_array(22901);
		when "0101100101110110" => data_out <= rom_array(22902);
		when "0101100101110111" => data_out <= rom_array(22903);
		when "0101100101111000" => data_out <= rom_array(22904);
		when "0101100101111001" => data_out <= rom_array(22905);
		when "0101100101111010" => data_out <= rom_array(22906);
		when "0101100101111011" => data_out <= rom_array(22907);
		when "0101100101111100" => data_out <= rom_array(22908);
		when "0101100101111101" => data_out <= rom_array(22909);
		when "0101100101111110" => data_out <= rom_array(22910);
		when "0101100101111111" => data_out <= rom_array(22911);
		when "0101100110000000" => data_out <= rom_array(22912);
		when "0101100110000001" => data_out <= rom_array(22913);
		when "0101100110000010" => data_out <= rom_array(22914);
		when "0101100110000011" => data_out <= rom_array(22915);
		when "0101100110000100" => data_out <= rom_array(22916);
		when "0101100110000101" => data_out <= rom_array(22917);
		when "0101100110000110" => data_out <= rom_array(22918);
		when "0101100110000111" => data_out <= rom_array(22919);
		when "0101100110001000" => data_out <= rom_array(22920);
		when "0101100110001001" => data_out <= rom_array(22921);
		when "0101100110001010" => data_out <= rom_array(22922);
		when "0101100110001011" => data_out <= rom_array(22923);
		when "0101100110001100" => data_out <= rom_array(22924);
		when "0101100110001101" => data_out <= rom_array(22925);
		when "0101100110001110" => data_out <= rom_array(22926);
		when "0101100110001111" => data_out <= rom_array(22927);
		when "0101100110010000" => data_out <= rom_array(22928);
		when "0101100110010001" => data_out <= rom_array(22929);
		when "0101100110010010" => data_out <= rom_array(22930);
		when "0101100110010011" => data_out <= rom_array(22931);
		when "0101100110010100" => data_out <= rom_array(22932);
		when "0101100110010101" => data_out <= rom_array(22933);
		when "0101100110010110" => data_out <= rom_array(22934);
		when "0101100110010111" => data_out <= rom_array(22935);
		when "0101100110011000" => data_out <= rom_array(22936);
		when "0101100110011001" => data_out <= rom_array(22937);
		when "0101100110011010" => data_out <= rom_array(22938);
		when "0101100110011011" => data_out <= rom_array(22939);
		when "0101100110011100" => data_out <= rom_array(22940);
		when "0101100110011101" => data_out <= rom_array(22941);
		when "0101100110011110" => data_out <= rom_array(22942);
		when "0101100110011111" => data_out <= rom_array(22943);
		when "0101100110100000" => data_out <= rom_array(22944);
		when "0101100110100001" => data_out <= rom_array(22945);
		when "0101100110100010" => data_out <= rom_array(22946);
		when "0101100110100011" => data_out <= rom_array(22947);
		when "0101100110100100" => data_out <= rom_array(22948);
		when "0101100110100101" => data_out <= rom_array(22949);
		when "0101100110100110" => data_out <= rom_array(22950);
		when "0101100110100111" => data_out <= rom_array(22951);
		when "0101100110101000" => data_out <= rom_array(22952);
		when "0101100110101001" => data_out <= rom_array(22953);
		when "0101100110101010" => data_out <= rom_array(22954);
		when "0101100110101011" => data_out <= rom_array(22955);
		when "0101100110101100" => data_out <= rom_array(22956);
		when "0101100110101101" => data_out <= rom_array(22957);
		when "0101100110101110" => data_out <= rom_array(22958);
		when "0101100110101111" => data_out <= rom_array(22959);
		when "0101100110110000" => data_out <= rom_array(22960);
		when "0101100110110001" => data_out <= rom_array(22961);
		when "0101100110110010" => data_out <= rom_array(22962);
		when "0101100110110011" => data_out <= rom_array(22963);
		when "0101100110110100" => data_out <= rom_array(22964);
		when "0101100110110101" => data_out <= rom_array(22965);
		when "0101100110110110" => data_out <= rom_array(22966);
		when "0101100110110111" => data_out <= rom_array(22967);
		when "0101100110111000" => data_out <= rom_array(22968);
		when "0101100110111001" => data_out <= rom_array(22969);
		when "0101100110111010" => data_out <= rom_array(22970);
		when "0101100110111011" => data_out <= rom_array(22971);
		when "0101100110111100" => data_out <= rom_array(22972);
		when "0101100110111101" => data_out <= rom_array(22973);
		when "0101100110111110" => data_out <= rom_array(22974);
		when "0101100110111111" => data_out <= rom_array(22975);
		when "0101100111000000" => data_out <= rom_array(22976);
		when "0101100111000001" => data_out <= rom_array(22977);
		when "0101100111000010" => data_out <= rom_array(22978);
		when "0101100111000011" => data_out <= rom_array(22979);
		when "0101100111000100" => data_out <= rom_array(22980);
		when "0101100111000101" => data_out <= rom_array(22981);
		when "0101100111000110" => data_out <= rom_array(22982);
		when "0101100111000111" => data_out <= rom_array(22983);
		when "0101100111001000" => data_out <= rom_array(22984);
		when "0101100111001001" => data_out <= rom_array(22985);
		when "0101100111001010" => data_out <= rom_array(22986);
		when "0101100111001011" => data_out <= rom_array(22987);
		when "0101100111001100" => data_out <= rom_array(22988);
		when "0101100111001101" => data_out <= rom_array(22989);
		when "0101100111001110" => data_out <= rom_array(22990);
		when "0101100111001111" => data_out <= rom_array(22991);
		when "0101100111010000" => data_out <= rom_array(22992);
		when "0101100111010001" => data_out <= rom_array(22993);
		when "0101100111010010" => data_out <= rom_array(22994);
		when "0101100111010011" => data_out <= rom_array(22995);
		when "0101100111010100" => data_out <= rom_array(22996);
		when "0101100111010101" => data_out <= rom_array(22997);
		when "0101100111010110" => data_out <= rom_array(22998);
		when "0101100111010111" => data_out <= rom_array(22999);
		when "0101100111011000" => data_out <= rom_array(23000);
		when "0101100111011001" => data_out <= rom_array(23001);
		when "0101100111011010" => data_out <= rom_array(23002);
		when "0101100111011011" => data_out <= rom_array(23003);
		when "0101100111011100" => data_out <= rom_array(23004);
		when "0101100111011101" => data_out <= rom_array(23005);
		when "0101100111011110" => data_out <= rom_array(23006);
		when "0101100111011111" => data_out <= rom_array(23007);
		when "0101100111100000" => data_out <= rom_array(23008);
		when "0101100111100001" => data_out <= rom_array(23009);
		when "0101100111100010" => data_out <= rom_array(23010);
		when "0101100111100011" => data_out <= rom_array(23011);
		when "0101100111100100" => data_out <= rom_array(23012);
		when "0101100111100101" => data_out <= rom_array(23013);
		when "0101100111100110" => data_out <= rom_array(23014);
		when "0101100111100111" => data_out <= rom_array(23015);
		when "0101100111101000" => data_out <= rom_array(23016);
		when "0101100111101001" => data_out <= rom_array(23017);
		when "0101100111101010" => data_out <= rom_array(23018);
		when "0101100111101011" => data_out <= rom_array(23019);
		when "0101100111101100" => data_out <= rom_array(23020);
		when "0101100111101101" => data_out <= rom_array(23021);
		when "0101100111101110" => data_out <= rom_array(23022);
		when "0101100111101111" => data_out <= rom_array(23023);
		when "0101100111110000" => data_out <= rom_array(23024);
		when "0101100111110001" => data_out <= rom_array(23025);
		when "0101100111110010" => data_out <= rom_array(23026);
		when "0101100111110011" => data_out <= rom_array(23027);
		when "0101100111110100" => data_out <= rom_array(23028);
		when "0101100111110101" => data_out <= rom_array(23029);
		when "0101100111110110" => data_out <= rom_array(23030);
		when "0101100111110111" => data_out <= rom_array(23031);
		when "0101100111111000" => data_out <= rom_array(23032);
		when "0101100111111001" => data_out <= rom_array(23033);
		when "0101100111111010" => data_out <= rom_array(23034);
		when "0101100111111011" => data_out <= rom_array(23035);
		when "0101100111111100" => data_out <= rom_array(23036);
		when "0101100111111101" => data_out <= rom_array(23037);
		when "0101100111111110" => data_out <= rom_array(23038);
		when "0101100111111111" => data_out <= rom_array(23039);
		when "0101101000000000" => data_out <= rom_array(23040);
		when "0101101000000001" => data_out <= rom_array(23041);
		when "0101101000000010" => data_out <= rom_array(23042);
		when "0101101000000011" => data_out <= rom_array(23043);
		when "0101101000000100" => data_out <= rom_array(23044);
		when "0101101000000101" => data_out <= rom_array(23045);
		when "0101101000000110" => data_out <= rom_array(23046);
		when "0101101000000111" => data_out <= rom_array(23047);
		when "0101101000001000" => data_out <= rom_array(23048);
		when "0101101000001001" => data_out <= rom_array(23049);
		when "0101101000001010" => data_out <= rom_array(23050);
		when "0101101000001011" => data_out <= rom_array(23051);
		when "0101101000001100" => data_out <= rom_array(23052);
		when "0101101000001101" => data_out <= rom_array(23053);
		when "0101101000001110" => data_out <= rom_array(23054);
		when "0101101000001111" => data_out <= rom_array(23055);
		when "0101101000010000" => data_out <= rom_array(23056);
		when "0101101000010001" => data_out <= rom_array(23057);
		when "0101101000010010" => data_out <= rom_array(23058);
		when "0101101000010011" => data_out <= rom_array(23059);
		when "0101101000010100" => data_out <= rom_array(23060);
		when "0101101000010101" => data_out <= rom_array(23061);
		when "0101101000010110" => data_out <= rom_array(23062);
		when "0101101000010111" => data_out <= rom_array(23063);
		when "0101101000011000" => data_out <= rom_array(23064);
		when "0101101000011001" => data_out <= rom_array(23065);
		when "0101101000011010" => data_out <= rom_array(23066);
		when "0101101000011011" => data_out <= rom_array(23067);
		when "0101101000011100" => data_out <= rom_array(23068);
		when "0101101000011101" => data_out <= rom_array(23069);
		when "0101101000011110" => data_out <= rom_array(23070);
		when "0101101000011111" => data_out <= rom_array(23071);
		when "0101101000100000" => data_out <= rom_array(23072);
		when "0101101000100001" => data_out <= rom_array(23073);
		when "0101101000100010" => data_out <= rom_array(23074);
		when "0101101000100011" => data_out <= rom_array(23075);
		when "0101101000100100" => data_out <= rom_array(23076);
		when "0101101000100101" => data_out <= rom_array(23077);
		when "0101101000100110" => data_out <= rom_array(23078);
		when "0101101000100111" => data_out <= rom_array(23079);
		when "0101101000101000" => data_out <= rom_array(23080);
		when "0101101000101001" => data_out <= rom_array(23081);
		when "0101101000101010" => data_out <= rom_array(23082);
		when "0101101000101011" => data_out <= rom_array(23083);
		when "0101101000101100" => data_out <= rom_array(23084);
		when "0101101000101101" => data_out <= rom_array(23085);
		when "0101101000101110" => data_out <= rom_array(23086);
		when "0101101000101111" => data_out <= rom_array(23087);
		when "0101101000110000" => data_out <= rom_array(23088);
		when "0101101000110001" => data_out <= rom_array(23089);
		when "0101101000110010" => data_out <= rom_array(23090);
		when "0101101000110011" => data_out <= rom_array(23091);
		when "0101101000110100" => data_out <= rom_array(23092);
		when "0101101000110101" => data_out <= rom_array(23093);
		when "0101101000110110" => data_out <= rom_array(23094);
		when "0101101000110111" => data_out <= rom_array(23095);
		when "0101101000111000" => data_out <= rom_array(23096);
		when "0101101000111001" => data_out <= rom_array(23097);
		when "0101101000111010" => data_out <= rom_array(23098);
		when "0101101000111011" => data_out <= rom_array(23099);
		when "0101101000111100" => data_out <= rom_array(23100);
		when "0101101000111101" => data_out <= rom_array(23101);
		when "0101101000111110" => data_out <= rom_array(23102);
		when "0101101000111111" => data_out <= rom_array(23103);
		when "0101101001000000" => data_out <= rom_array(23104);
		when "0101101001000001" => data_out <= rom_array(23105);
		when "0101101001000010" => data_out <= rom_array(23106);
		when "0101101001000011" => data_out <= rom_array(23107);
		when "0101101001000100" => data_out <= rom_array(23108);
		when "0101101001000101" => data_out <= rom_array(23109);
		when "0101101001000110" => data_out <= rom_array(23110);
		when "0101101001000111" => data_out <= rom_array(23111);
		when "0101101001001000" => data_out <= rom_array(23112);
		when "0101101001001001" => data_out <= rom_array(23113);
		when "0101101001001010" => data_out <= rom_array(23114);
		when "0101101001001011" => data_out <= rom_array(23115);
		when "0101101001001100" => data_out <= rom_array(23116);
		when "0101101001001101" => data_out <= rom_array(23117);
		when "0101101001001110" => data_out <= rom_array(23118);
		when "0101101001001111" => data_out <= rom_array(23119);
		when "0101101001010000" => data_out <= rom_array(23120);
		when "0101101001010001" => data_out <= rom_array(23121);
		when "0101101001010010" => data_out <= rom_array(23122);
		when "0101101001010011" => data_out <= rom_array(23123);
		when "0101101001010100" => data_out <= rom_array(23124);
		when "0101101001010101" => data_out <= rom_array(23125);
		when "0101101001010110" => data_out <= rom_array(23126);
		when "0101101001010111" => data_out <= rom_array(23127);
		when "0101101001011000" => data_out <= rom_array(23128);
		when "0101101001011001" => data_out <= rom_array(23129);
		when "0101101001011010" => data_out <= rom_array(23130);
		when "0101101001011011" => data_out <= rom_array(23131);
		when "0101101001011100" => data_out <= rom_array(23132);
		when "0101101001011101" => data_out <= rom_array(23133);
		when "0101101001011110" => data_out <= rom_array(23134);
		when "0101101001011111" => data_out <= rom_array(23135);
		when "0101101001100000" => data_out <= rom_array(23136);
		when "0101101001100001" => data_out <= rom_array(23137);
		when "0101101001100010" => data_out <= rom_array(23138);
		when "0101101001100011" => data_out <= rom_array(23139);
		when "0101101001100100" => data_out <= rom_array(23140);
		when "0101101001100101" => data_out <= rom_array(23141);
		when "0101101001100110" => data_out <= rom_array(23142);
		when "0101101001100111" => data_out <= rom_array(23143);
		when "0101101001101000" => data_out <= rom_array(23144);
		when "0101101001101001" => data_out <= rom_array(23145);
		when "0101101001101010" => data_out <= rom_array(23146);
		when "0101101001101011" => data_out <= rom_array(23147);
		when "0101101001101100" => data_out <= rom_array(23148);
		when "0101101001101101" => data_out <= rom_array(23149);
		when "0101101001101110" => data_out <= rom_array(23150);
		when "0101101001101111" => data_out <= rom_array(23151);
		when "0101101001110000" => data_out <= rom_array(23152);
		when "0101101001110001" => data_out <= rom_array(23153);
		when "0101101001110010" => data_out <= rom_array(23154);
		when "0101101001110011" => data_out <= rom_array(23155);
		when "0101101001110100" => data_out <= rom_array(23156);
		when "0101101001110101" => data_out <= rom_array(23157);
		when "0101101001110110" => data_out <= rom_array(23158);
		when "0101101001110111" => data_out <= rom_array(23159);
		when "0101101001111000" => data_out <= rom_array(23160);
		when "0101101001111001" => data_out <= rom_array(23161);
		when "0101101001111010" => data_out <= rom_array(23162);
		when "0101101001111011" => data_out <= rom_array(23163);
		when "0101101001111100" => data_out <= rom_array(23164);
		when "0101101001111101" => data_out <= rom_array(23165);
		when "0101101001111110" => data_out <= rom_array(23166);
		when "0101101001111111" => data_out <= rom_array(23167);
		when "0101101010000000" => data_out <= rom_array(23168);
		when "0101101010000001" => data_out <= rom_array(23169);
		when "0101101010000010" => data_out <= rom_array(23170);
		when "0101101010000011" => data_out <= rom_array(23171);
		when "0101101010000100" => data_out <= rom_array(23172);
		when "0101101010000101" => data_out <= rom_array(23173);
		when "0101101010000110" => data_out <= rom_array(23174);
		when "0101101010000111" => data_out <= rom_array(23175);
		when "0101101010001000" => data_out <= rom_array(23176);
		when "0101101010001001" => data_out <= rom_array(23177);
		when "0101101010001010" => data_out <= rom_array(23178);
		when "0101101010001011" => data_out <= rom_array(23179);
		when "0101101010001100" => data_out <= rom_array(23180);
		when "0101101010001101" => data_out <= rom_array(23181);
		when "0101101010001110" => data_out <= rom_array(23182);
		when "0101101010001111" => data_out <= rom_array(23183);
		when "0101101010010000" => data_out <= rom_array(23184);
		when "0101101010010001" => data_out <= rom_array(23185);
		when "0101101010010010" => data_out <= rom_array(23186);
		when "0101101010010011" => data_out <= rom_array(23187);
		when "0101101010010100" => data_out <= rom_array(23188);
		when "0101101010010101" => data_out <= rom_array(23189);
		when "0101101010010110" => data_out <= rom_array(23190);
		when "0101101010010111" => data_out <= rom_array(23191);
		when "0101101010011000" => data_out <= rom_array(23192);
		when "0101101010011001" => data_out <= rom_array(23193);
		when "0101101010011010" => data_out <= rom_array(23194);
		when "0101101010011011" => data_out <= rom_array(23195);
		when "0101101010011100" => data_out <= rom_array(23196);
		when "0101101010011101" => data_out <= rom_array(23197);
		when "0101101010011110" => data_out <= rom_array(23198);
		when "0101101010011111" => data_out <= rom_array(23199);
		when "0101101010100000" => data_out <= rom_array(23200);
		when "0101101010100001" => data_out <= rom_array(23201);
		when "0101101010100010" => data_out <= rom_array(23202);
		when "0101101010100011" => data_out <= rom_array(23203);
		when "0101101010100100" => data_out <= rom_array(23204);
		when "0101101010100101" => data_out <= rom_array(23205);
		when "0101101010100110" => data_out <= rom_array(23206);
		when "0101101010100111" => data_out <= rom_array(23207);
		when "0101101010101000" => data_out <= rom_array(23208);
		when "0101101010101001" => data_out <= rom_array(23209);
		when "0101101010101010" => data_out <= rom_array(23210);
		when "0101101010101011" => data_out <= rom_array(23211);
		when "0101101010101100" => data_out <= rom_array(23212);
		when "0101101010101101" => data_out <= rom_array(23213);
		when "0101101010101110" => data_out <= rom_array(23214);
		when "0101101010101111" => data_out <= rom_array(23215);
		when "0101101010110000" => data_out <= rom_array(23216);
		when "0101101010110001" => data_out <= rom_array(23217);
		when "0101101010110010" => data_out <= rom_array(23218);
		when "0101101010110011" => data_out <= rom_array(23219);
		when "0101101010110100" => data_out <= rom_array(23220);
		when "0101101010110101" => data_out <= rom_array(23221);
		when "0101101010110110" => data_out <= rom_array(23222);
		when "0101101010110111" => data_out <= rom_array(23223);
		when "0101101010111000" => data_out <= rom_array(23224);
		when "0101101010111001" => data_out <= rom_array(23225);
		when "0101101010111010" => data_out <= rom_array(23226);
		when "0101101010111011" => data_out <= rom_array(23227);
		when "0101101010111100" => data_out <= rom_array(23228);
		when "0101101010111101" => data_out <= rom_array(23229);
		when "0101101010111110" => data_out <= rom_array(23230);
		when "0101101010111111" => data_out <= rom_array(23231);
		when "0101101011000000" => data_out <= rom_array(23232);
		when "0101101011000001" => data_out <= rom_array(23233);
		when "0101101011000010" => data_out <= rom_array(23234);
		when "0101101011000011" => data_out <= rom_array(23235);
		when "0101101011000100" => data_out <= rom_array(23236);
		when "0101101011000101" => data_out <= rom_array(23237);
		when "0101101011000110" => data_out <= rom_array(23238);
		when "0101101011000111" => data_out <= rom_array(23239);
		when "0101101011001000" => data_out <= rom_array(23240);
		when "0101101011001001" => data_out <= rom_array(23241);
		when "0101101011001010" => data_out <= rom_array(23242);
		when "0101101011001011" => data_out <= rom_array(23243);
		when "0101101011001100" => data_out <= rom_array(23244);
		when "0101101011001101" => data_out <= rom_array(23245);
		when "0101101011001110" => data_out <= rom_array(23246);
		when "0101101011001111" => data_out <= rom_array(23247);
		when "0101101011010000" => data_out <= rom_array(23248);
		when "0101101011010001" => data_out <= rom_array(23249);
		when "0101101011010010" => data_out <= rom_array(23250);
		when "0101101011010011" => data_out <= rom_array(23251);
		when "0101101011010100" => data_out <= rom_array(23252);
		when "0101101011010101" => data_out <= rom_array(23253);
		when "0101101011010110" => data_out <= rom_array(23254);
		when "0101101011010111" => data_out <= rom_array(23255);
		when "0101101011011000" => data_out <= rom_array(23256);
		when "0101101011011001" => data_out <= rom_array(23257);
		when "0101101011011010" => data_out <= rom_array(23258);
		when "0101101011011011" => data_out <= rom_array(23259);
		when "0101101011011100" => data_out <= rom_array(23260);
		when "0101101011011101" => data_out <= rom_array(23261);
		when "0101101011011110" => data_out <= rom_array(23262);
		when "0101101011011111" => data_out <= rom_array(23263);
		when "0101101011100000" => data_out <= rom_array(23264);
		when "0101101011100001" => data_out <= rom_array(23265);
		when "0101101011100010" => data_out <= rom_array(23266);
		when "0101101011100011" => data_out <= rom_array(23267);
		when "0101101011100100" => data_out <= rom_array(23268);
		when "0101101011100101" => data_out <= rom_array(23269);
		when "0101101011100110" => data_out <= rom_array(23270);
		when "0101101011100111" => data_out <= rom_array(23271);
		when "0101101011101000" => data_out <= rom_array(23272);
		when "0101101011101001" => data_out <= rom_array(23273);
		when "0101101011101010" => data_out <= rom_array(23274);
		when "0101101011101011" => data_out <= rom_array(23275);
		when "0101101011101100" => data_out <= rom_array(23276);
		when "0101101011101101" => data_out <= rom_array(23277);
		when "0101101011101110" => data_out <= rom_array(23278);
		when "0101101011101111" => data_out <= rom_array(23279);
		when "0101101011110000" => data_out <= rom_array(23280);
		when "0101101011110001" => data_out <= rom_array(23281);
		when "0101101011110010" => data_out <= rom_array(23282);
		when "0101101011110011" => data_out <= rom_array(23283);
		when "0101101011110100" => data_out <= rom_array(23284);
		when "0101101011110101" => data_out <= rom_array(23285);
		when "0101101011110110" => data_out <= rom_array(23286);
		when "0101101011110111" => data_out <= rom_array(23287);
		when "0101101011111000" => data_out <= rom_array(23288);
		when "0101101011111001" => data_out <= rom_array(23289);
		when "0101101011111010" => data_out <= rom_array(23290);
		when "0101101011111011" => data_out <= rom_array(23291);
		when "0101101011111100" => data_out <= rom_array(23292);
		when "0101101011111101" => data_out <= rom_array(23293);
		when "0101101011111110" => data_out <= rom_array(23294);
		when "0101101011111111" => data_out <= rom_array(23295);
		when "0101101100000000" => data_out <= rom_array(23296);
		when "0101101100000001" => data_out <= rom_array(23297);
		when "0101101100000010" => data_out <= rom_array(23298);
		when "0101101100000011" => data_out <= rom_array(23299);
		when "0101101100000100" => data_out <= rom_array(23300);
		when "0101101100000101" => data_out <= rom_array(23301);
		when "0101101100000110" => data_out <= rom_array(23302);
		when "0101101100000111" => data_out <= rom_array(23303);
		when "0101101100001000" => data_out <= rom_array(23304);
		when "0101101100001001" => data_out <= rom_array(23305);
		when "0101101100001010" => data_out <= rom_array(23306);
		when "0101101100001011" => data_out <= rom_array(23307);
		when "0101101100001100" => data_out <= rom_array(23308);
		when "0101101100001101" => data_out <= rom_array(23309);
		when "0101101100001110" => data_out <= rom_array(23310);
		when "0101101100001111" => data_out <= rom_array(23311);
		when "0101101100010000" => data_out <= rom_array(23312);
		when "0101101100010001" => data_out <= rom_array(23313);
		when "0101101100010010" => data_out <= rom_array(23314);
		when "0101101100010011" => data_out <= rom_array(23315);
		when "0101101100010100" => data_out <= rom_array(23316);
		when "0101101100010101" => data_out <= rom_array(23317);
		when "0101101100010110" => data_out <= rom_array(23318);
		when "0101101100010111" => data_out <= rom_array(23319);
		when "0101101100011000" => data_out <= rom_array(23320);
		when "0101101100011001" => data_out <= rom_array(23321);
		when "0101101100011010" => data_out <= rom_array(23322);
		when "0101101100011011" => data_out <= rom_array(23323);
		when "0101101100011100" => data_out <= rom_array(23324);
		when "0101101100011101" => data_out <= rom_array(23325);
		when "0101101100011110" => data_out <= rom_array(23326);
		when "0101101100011111" => data_out <= rom_array(23327);
		when "0101101100100000" => data_out <= rom_array(23328);
		when "0101101100100001" => data_out <= rom_array(23329);
		when "0101101100100010" => data_out <= rom_array(23330);
		when "0101101100100011" => data_out <= rom_array(23331);
		when "0101101100100100" => data_out <= rom_array(23332);
		when "0101101100100101" => data_out <= rom_array(23333);
		when "0101101100100110" => data_out <= rom_array(23334);
		when "0101101100100111" => data_out <= rom_array(23335);
		when "0101101100101000" => data_out <= rom_array(23336);
		when "0101101100101001" => data_out <= rom_array(23337);
		when "0101101100101010" => data_out <= rom_array(23338);
		when "0101101100101011" => data_out <= rom_array(23339);
		when "0101101100101100" => data_out <= rom_array(23340);
		when "0101101100101101" => data_out <= rom_array(23341);
		when "0101101100101110" => data_out <= rom_array(23342);
		when "0101101100101111" => data_out <= rom_array(23343);
		when "0101101100110000" => data_out <= rom_array(23344);
		when "0101101100110001" => data_out <= rom_array(23345);
		when "0101101100110010" => data_out <= rom_array(23346);
		when "0101101100110011" => data_out <= rom_array(23347);
		when "0101101100110100" => data_out <= rom_array(23348);
		when "0101101100110101" => data_out <= rom_array(23349);
		when "0101101100110110" => data_out <= rom_array(23350);
		when "0101101100110111" => data_out <= rom_array(23351);
		when "0101101100111000" => data_out <= rom_array(23352);
		when "0101101100111001" => data_out <= rom_array(23353);
		when "0101101100111010" => data_out <= rom_array(23354);
		when "0101101100111011" => data_out <= rom_array(23355);
		when "0101101100111100" => data_out <= rom_array(23356);
		when "0101101100111101" => data_out <= rom_array(23357);
		when "0101101100111110" => data_out <= rom_array(23358);
		when "0101101100111111" => data_out <= rom_array(23359);
		when "0101101101000000" => data_out <= rom_array(23360);
		when "0101101101000001" => data_out <= rom_array(23361);
		when "0101101101000010" => data_out <= rom_array(23362);
		when "0101101101000011" => data_out <= rom_array(23363);
		when "0101101101000100" => data_out <= rom_array(23364);
		when "0101101101000101" => data_out <= rom_array(23365);
		when "0101101101000110" => data_out <= rom_array(23366);
		when "0101101101000111" => data_out <= rom_array(23367);
		when "0101101101001000" => data_out <= rom_array(23368);
		when "0101101101001001" => data_out <= rom_array(23369);
		when "0101101101001010" => data_out <= rom_array(23370);
		when "0101101101001011" => data_out <= rom_array(23371);
		when "0101101101001100" => data_out <= rom_array(23372);
		when "0101101101001101" => data_out <= rom_array(23373);
		when "0101101101001110" => data_out <= rom_array(23374);
		when "0101101101001111" => data_out <= rom_array(23375);
		when "0101101101010000" => data_out <= rom_array(23376);
		when "0101101101010001" => data_out <= rom_array(23377);
		when "0101101101010010" => data_out <= rom_array(23378);
		when "0101101101010011" => data_out <= rom_array(23379);
		when "0101101101010100" => data_out <= rom_array(23380);
		when "0101101101010101" => data_out <= rom_array(23381);
		when "0101101101010110" => data_out <= rom_array(23382);
		when "0101101101010111" => data_out <= rom_array(23383);
		when "0101101101011000" => data_out <= rom_array(23384);
		when "0101101101011001" => data_out <= rom_array(23385);
		when "0101101101011010" => data_out <= rom_array(23386);
		when "0101101101011011" => data_out <= rom_array(23387);
		when "0101101101011100" => data_out <= rom_array(23388);
		when "0101101101011101" => data_out <= rom_array(23389);
		when "0101101101011110" => data_out <= rom_array(23390);
		when "0101101101011111" => data_out <= rom_array(23391);
		when "0101101101100000" => data_out <= rom_array(23392);
		when "0101101101100001" => data_out <= rom_array(23393);
		when "0101101101100010" => data_out <= rom_array(23394);
		when "0101101101100011" => data_out <= rom_array(23395);
		when "0101101101100100" => data_out <= rom_array(23396);
		when "0101101101100101" => data_out <= rom_array(23397);
		when "0101101101100110" => data_out <= rom_array(23398);
		when "0101101101100111" => data_out <= rom_array(23399);
		when "0101101101101000" => data_out <= rom_array(23400);
		when "0101101101101001" => data_out <= rom_array(23401);
		when "0101101101101010" => data_out <= rom_array(23402);
		when "0101101101101011" => data_out <= rom_array(23403);
		when "0101101101101100" => data_out <= rom_array(23404);
		when "0101101101101101" => data_out <= rom_array(23405);
		when "0101101101101110" => data_out <= rom_array(23406);
		when "0101101101101111" => data_out <= rom_array(23407);
		when "0101101101110000" => data_out <= rom_array(23408);
		when "0101101101110001" => data_out <= rom_array(23409);
		when "0101101101110010" => data_out <= rom_array(23410);
		when "0101101101110011" => data_out <= rom_array(23411);
		when "0101101101110100" => data_out <= rom_array(23412);
		when "0101101101110101" => data_out <= rom_array(23413);
		when "0101101101110110" => data_out <= rom_array(23414);
		when "0101101101110111" => data_out <= rom_array(23415);
		when "0101101101111000" => data_out <= rom_array(23416);
		when "0101101101111001" => data_out <= rom_array(23417);
		when "0101101101111010" => data_out <= rom_array(23418);
		when "0101101101111011" => data_out <= rom_array(23419);
		when "0101101101111100" => data_out <= rom_array(23420);
		when "0101101101111101" => data_out <= rom_array(23421);
		when "0101101101111110" => data_out <= rom_array(23422);
		when "0101101101111111" => data_out <= rom_array(23423);
		when "0101101110000000" => data_out <= rom_array(23424);
		when "0101101110000001" => data_out <= rom_array(23425);
		when "0101101110000010" => data_out <= rom_array(23426);
		when "0101101110000011" => data_out <= rom_array(23427);
		when "0101101110000100" => data_out <= rom_array(23428);
		when "0101101110000101" => data_out <= rom_array(23429);
		when "0101101110000110" => data_out <= rom_array(23430);
		when "0101101110000111" => data_out <= rom_array(23431);
		when "0101101110001000" => data_out <= rom_array(23432);
		when "0101101110001001" => data_out <= rom_array(23433);
		when "0101101110001010" => data_out <= rom_array(23434);
		when "0101101110001011" => data_out <= rom_array(23435);
		when "0101101110001100" => data_out <= rom_array(23436);
		when "0101101110001101" => data_out <= rom_array(23437);
		when "0101101110001110" => data_out <= rom_array(23438);
		when "0101101110001111" => data_out <= rom_array(23439);
		when "0101101110010000" => data_out <= rom_array(23440);
		when "0101101110010001" => data_out <= rom_array(23441);
		when "0101101110010010" => data_out <= rom_array(23442);
		when "0101101110010011" => data_out <= rom_array(23443);
		when "0101101110010100" => data_out <= rom_array(23444);
		when "0101101110010101" => data_out <= rom_array(23445);
		when "0101101110010110" => data_out <= rom_array(23446);
		when "0101101110010111" => data_out <= rom_array(23447);
		when "0101101110011000" => data_out <= rom_array(23448);
		when "0101101110011001" => data_out <= rom_array(23449);
		when "0101101110011010" => data_out <= rom_array(23450);
		when "0101101110011011" => data_out <= rom_array(23451);
		when "0101101110011100" => data_out <= rom_array(23452);
		when "0101101110011101" => data_out <= rom_array(23453);
		when "0101101110011110" => data_out <= rom_array(23454);
		when "0101101110011111" => data_out <= rom_array(23455);
		when "0101101110100000" => data_out <= rom_array(23456);
		when "0101101110100001" => data_out <= rom_array(23457);
		when "0101101110100010" => data_out <= rom_array(23458);
		when "0101101110100011" => data_out <= rom_array(23459);
		when "0101101110100100" => data_out <= rom_array(23460);
		when "0101101110100101" => data_out <= rom_array(23461);
		when "0101101110100110" => data_out <= rom_array(23462);
		when "0101101110100111" => data_out <= rom_array(23463);
		when "0101101110101000" => data_out <= rom_array(23464);
		when "0101101110101001" => data_out <= rom_array(23465);
		when "0101101110101010" => data_out <= rom_array(23466);
		when "0101101110101011" => data_out <= rom_array(23467);
		when "0101101110101100" => data_out <= rom_array(23468);
		when "0101101110101101" => data_out <= rom_array(23469);
		when "0101101110101110" => data_out <= rom_array(23470);
		when "0101101110101111" => data_out <= rom_array(23471);
		when "0101101110110000" => data_out <= rom_array(23472);
		when "0101101110110001" => data_out <= rom_array(23473);
		when "0101101110110010" => data_out <= rom_array(23474);
		when "0101101110110011" => data_out <= rom_array(23475);
		when "0101101110110100" => data_out <= rom_array(23476);
		when "0101101110110101" => data_out <= rom_array(23477);
		when "0101101110110110" => data_out <= rom_array(23478);
		when "0101101110110111" => data_out <= rom_array(23479);
		when "0101101110111000" => data_out <= rom_array(23480);
		when "0101101110111001" => data_out <= rom_array(23481);
		when "0101101110111010" => data_out <= rom_array(23482);
		when "0101101110111011" => data_out <= rom_array(23483);
		when "0101101110111100" => data_out <= rom_array(23484);
		when "0101101110111101" => data_out <= rom_array(23485);
		when "0101101110111110" => data_out <= rom_array(23486);
		when "0101101110111111" => data_out <= rom_array(23487);
		when "0101101111000000" => data_out <= rom_array(23488);
		when "0101101111000001" => data_out <= rom_array(23489);
		when "0101101111000010" => data_out <= rom_array(23490);
		when "0101101111000011" => data_out <= rom_array(23491);
		when "0101101111000100" => data_out <= rom_array(23492);
		when "0101101111000101" => data_out <= rom_array(23493);
		when "0101101111000110" => data_out <= rom_array(23494);
		when "0101101111000111" => data_out <= rom_array(23495);
		when "0101101111001000" => data_out <= rom_array(23496);
		when "0101101111001001" => data_out <= rom_array(23497);
		when "0101101111001010" => data_out <= rom_array(23498);
		when "0101101111001011" => data_out <= rom_array(23499);
		when "0101101111001100" => data_out <= rom_array(23500);
		when "0101101111001101" => data_out <= rom_array(23501);
		when "0101101111001110" => data_out <= rom_array(23502);
		when "0101101111001111" => data_out <= rom_array(23503);
		when "0101101111010000" => data_out <= rom_array(23504);
		when "0101101111010001" => data_out <= rom_array(23505);
		when "0101101111010010" => data_out <= rom_array(23506);
		when "0101101111010011" => data_out <= rom_array(23507);
		when "0101101111010100" => data_out <= rom_array(23508);
		when "0101101111010101" => data_out <= rom_array(23509);
		when "0101101111010110" => data_out <= rom_array(23510);
		when "0101101111010111" => data_out <= rom_array(23511);
		when "0101101111011000" => data_out <= rom_array(23512);
		when "0101101111011001" => data_out <= rom_array(23513);
		when "0101101111011010" => data_out <= rom_array(23514);
		when "0101101111011011" => data_out <= rom_array(23515);
		when "0101101111011100" => data_out <= rom_array(23516);
		when "0101101111011101" => data_out <= rom_array(23517);
		when "0101101111011110" => data_out <= rom_array(23518);
		when "0101101111011111" => data_out <= rom_array(23519);
		when "0101101111100000" => data_out <= rom_array(23520);
		when "0101101111100001" => data_out <= rom_array(23521);
		when "0101101111100010" => data_out <= rom_array(23522);
		when "0101101111100011" => data_out <= rom_array(23523);
		when "0101101111100100" => data_out <= rom_array(23524);
		when "0101101111100101" => data_out <= rom_array(23525);
		when "0101101111100110" => data_out <= rom_array(23526);
		when "0101101111100111" => data_out <= rom_array(23527);
		when "0101101111101000" => data_out <= rom_array(23528);
		when "0101101111101001" => data_out <= rom_array(23529);
		when "0101101111101010" => data_out <= rom_array(23530);
		when "0101101111101011" => data_out <= rom_array(23531);
		when "0101101111101100" => data_out <= rom_array(23532);
		when "0101101111101101" => data_out <= rom_array(23533);
		when "0101101111101110" => data_out <= rom_array(23534);
		when "0101101111101111" => data_out <= rom_array(23535);
		when "0101101111110000" => data_out <= rom_array(23536);
		when "0101101111110001" => data_out <= rom_array(23537);
		when "0101101111110010" => data_out <= rom_array(23538);
		when "0101101111110011" => data_out <= rom_array(23539);
		when "0101101111110100" => data_out <= rom_array(23540);
		when "0101101111110101" => data_out <= rom_array(23541);
		when "0101101111110110" => data_out <= rom_array(23542);
		when "0101101111110111" => data_out <= rom_array(23543);
		when "0101101111111000" => data_out <= rom_array(23544);
		when "0101101111111001" => data_out <= rom_array(23545);
		when "0101101111111010" => data_out <= rom_array(23546);
		when "0101101111111011" => data_out <= rom_array(23547);
		when "0101101111111100" => data_out <= rom_array(23548);
		when "0101101111111101" => data_out <= rom_array(23549);
		when "0101101111111110" => data_out <= rom_array(23550);
		when "0101101111111111" => data_out <= rom_array(23551);
		when "0101110000000000" => data_out <= rom_array(23552);
		when "0101110000000001" => data_out <= rom_array(23553);
		when "0101110000000010" => data_out <= rom_array(23554);
		when "0101110000000011" => data_out <= rom_array(23555);
		when "0101110000000100" => data_out <= rom_array(23556);
		when "0101110000000101" => data_out <= rom_array(23557);
		when "0101110000000110" => data_out <= rom_array(23558);
		when "0101110000000111" => data_out <= rom_array(23559);
		when "0101110000001000" => data_out <= rom_array(23560);
		when "0101110000001001" => data_out <= rom_array(23561);
		when "0101110000001010" => data_out <= rom_array(23562);
		when "0101110000001011" => data_out <= rom_array(23563);
		when "0101110000001100" => data_out <= rom_array(23564);
		when "0101110000001101" => data_out <= rom_array(23565);
		when "0101110000001110" => data_out <= rom_array(23566);
		when "0101110000001111" => data_out <= rom_array(23567);
		when "0101110000010000" => data_out <= rom_array(23568);
		when "0101110000010001" => data_out <= rom_array(23569);
		when "0101110000010010" => data_out <= rom_array(23570);
		when "0101110000010011" => data_out <= rom_array(23571);
		when "0101110000010100" => data_out <= rom_array(23572);
		when "0101110000010101" => data_out <= rom_array(23573);
		when "0101110000010110" => data_out <= rom_array(23574);
		when "0101110000010111" => data_out <= rom_array(23575);
		when "0101110000011000" => data_out <= rom_array(23576);
		when "0101110000011001" => data_out <= rom_array(23577);
		when "0101110000011010" => data_out <= rom_array(23578);
		when "0101110000011011" => data_out <= rom_array(23579);
		when "0101110000011100" => data_out <= rom_array(23580);
		when "0101110000011101" => data_out <= rom_array(23581);
		when "0101110000011110" => data_out <= rom_array(23582);
		when "0101110000011111" => data_out <= rom_array(23583);
		when "0101110000100000" => data_out <= rom_array(23584);
		when "0101110000100001" => data_out <= rom_array(23585);
		when "0101110000100010" => data_out <= rom_array(23586);
		when "0101110000100011" => data_out <= rom_array(23587);
		when "0101110000100100" => data_out <= rom_array(23588);
		when "0101110000100101" => data_out <= rom_array(23589);
		when "0101110000100110" => data_out <= rom_array(23590);
		when "0101110000100111" => data_out <= rom_array(23591);
		when "0101110000101000" => data_out <= rom_array(23592);
		when "0101110000101001" => data_out <= rom_array(23593);
		when "0101110000101010" => data_out <= rom_array(23594);
		when "0101110000101011" => data_out <= rom_array(23595);
		when "0101110000101100" => data_out <= rom_array(23596);
		when "0101110000101101" => data_out <= rom_array(23597);
		when "0101110000101110" => data_out <= rom_array(23598);
		when "0101110000101111" => data_out <= rom_array(23599);
		when "0101110000110000" => data_out <= rom_array(23600);
		when "0101110000110001" => data_out <= rom_array(23601);
		when "0101110000110010" => data_out <= rom_array(23602);
		when "0101110000110011" => data_out <= rom_array(23603);
		when "0101110000110100" => data_out <= rom_array(23604);
		when "0101110000110101" => data_out <= rom_array(23605);
		when "0101110000110110" => data_out <= rom_array(23606);
		when "0101110000110111" => data_out <= rom_array(23607);
		when "0101110000111000" => data_out <= rom_array(23608);
		when "0101110000111001" => data_out <= rom_array(23609);
		when "0101110000111010" => data_out <= rom_array(23610);
		when "0101110000111011" => data_out <= rom_array(23611);
		when "0101110000111100" => data_out <= rom_array(23612);
		when "0101110000111101" => data_out <= rom_array(23613);
		when "0101110000111110" => data_out <= rom_array(23614);
		when "0101110000111111" => data_out <= rom_array(23615);
		when "0101110001000000" => data_out <= rom_array(23616);
		when "0101110001000001" => data_out <= rom_array(23617);
		when "0101110001000010" => data_out <= rom_array(23618);
		when "0101110001000011" => data_out <= rom_array(23619);
		when "0101110001000100" => data_out <= rom_array(23620);
		when "0101110001000101" => data_out <= rom_array(23621);
		when "0101110001000110" => data_out <= rom_array(23622);
		when "0101110001000111" => data_out <= rom_array(23623);
		when "0101110001001000" => data_out <= rom_array(23624);
		when "0101110001001001" => data_out <= rom_array(23625);
		when "0101110001001010" => data_out <= rom_array(23626);
		when "0101110001001011" => data_out <= rom_array(23627);
		when "0101110001001100" => data_out <= rom_array(23628);
		when "0101110001001101" => data_out <= rom_array(23629);
		when "0101110001001110" => data_out <= rom_array(23630);
		when "0101110001001111" => data_out <= rom_array(23631);
		when "0101110001010000" => data_out <= rom_array(23632);
		when "0101110001010001" => data_out <= rom_array(23633);
		when "0101110001010010" => data_out <= rom_array(23634);
		when "0101110001010011" => data_out <= rom_array(23635);
		when "0101110001010100" => data_out <= rom_array(23636);
		when "0101110001010101" => data_out <= rom_array(23637);
		when "0101110001010110" => data_out <= rom_array(23638);
		when "0101110001010111" => data_out <= rom_array(23639);
		when "0101110001011000" => data_out <= rom_array(23640);
		when "0101110001011001" => data_out <= rom_array(23641);
		when "0101110001011010" => data_out <= rom_array(23642);
		when "0101110001011011" => data_out <= rom_array(23643);
		when "0101110001011100" => data_out <= rom_array(23644);
		when "0101110001011101" => data_out <= rom_array(23645);
		when "0101110001011110" => data_out <= rom_array(23646);
		when "0101110001011111" => data_out <= rom_array(23647);
		when "0101110001100000" => data_out <= rom_array(23648);
		when "0101110001100001" => data_out <= rom_array(23649);
		when "0101110001100010" => data_out <= rom_array(23650);
		when "0101110001100011" => data_out <= rom_array(23651);
		when "0101110001100100" => data_out <= rom_array(23652);
		when "0101110001100101" => data_out <= rom_array(23653);
		when "0101110001100110" => data_out <= rom_array(23654);
		when "0101110001100111" => data_out <= rom_array(23655);
		when "0101110001101000" => data_out <= rom_array(23656);
		when "0101110001101001" => data_out <= rom_array(23657);
		when "0101110001101010" => data_out <= rom_array(23658);
		when "0101110001101011" => data_out <= rom_array(23659);
		when "0101110001101100" => data_out <= rom_array(23660);
		when "0101110001101101" => data_out <= rom_array(23661);
		when "0101110001101110" => data_out <= rom_array(23662);
		when "0101110001101111" => data_out <= rom_array(23663);
		when "0101110001110000" => data_out <= rom_array(23664);
		when "0101110001110001" => data_out <= rom_array(23665);
		when "0101110001110010" => data_out <= rom_array(23666);
		when "0101110001110011" => data_out <= rom_array(23667);
		when "0101110001110100" => data_out <= rom_array(23668);
		when "0101110001110101" => data_out <= rom_array(23669);
		when "0101110001110110" => data_out <= rom_array(23670);
		when "0101110001110111" => data_out <= rom_array(23671);
		when "0101110001111000" => data_out <= rom_array(23672);
		when "0101110001111001" => data_out <= rom_array(23673);
		when "0101110001111010" => data_out <= rom_array(23674);
		when "0101110001111011" => data_out <= rom_array(23675);
		when "0101110001111100" => data_out <= rom_array(23676);
		when "0101110001111101" => data_out <= rom_array(23677);
		when "0101110001111110" => data_out <= rom_array(23678);
		when "0101110001111111" => data_out <= rom_array(23679);
		when "0101110010000000" => data_out <= rom_array(23680);
		when "0101110010000001" => data_out <= rom_array(23681);
		when "0101110010000010" => data_out <= rom_array(23682);
		when "0101110010000011" => data_out <= rom_array(23683);
		when "0101110010000100" => data_out <= rom_array(23684);
		when "0101110010000101" => data_out <= rom_array(23685);
		when "0101110010000110" => data_out <= rom_array(23686);
		when "0101110010000111" => data_out <= rom_array(23687);
		when "0101110010001000" => data_out <= rom_array(23688);
		when "0101110010001001" => data_out <= rom_array(23689);
		when "0101110010001010" => data_out <= rom_array(23690);
		when "0101110010001011" => data_out <= rom_array(23691);
		when "0101110010001100" => data_out <= rom_array(23692);
		when "0101110010001101" => data_out <= rom_array(23693);
		when "0101110010001110" => data_out <= rom_array(23694);
		when "0101110010001111" => data_out <= rom_array(23695);
		when "0101110010010000" => data_out <= rom_array(23696);
		when "0101110010010001" => data_out <= rom_array(23697);
		when "0101110010010010" => data_out <= rom_array(23698);
		when "0101110010010011" => data_out <= rom_array(23699);
		when "0101110010010100" => data_out <= rom_array(23700);
		when "0101110010010101" => data_out <= rom_array(23701);
		when "0101110010010110" => data_out <= rom_array(23702);
		when "0101110010010111" => data_out <= rom_array(23703);
		when "0101110010011000" => data_out <= rom_array(23704);
		when "0101110010011001" => data_out <= rom_array(23705);
		when "0101110010011010" => data_out <= rom_array(23706);
		when "0101110010011011" => data_out <= rom_array(23707);
		when "0101110010011100" => data_out <= rom_array(23708);
		when "0101110010011101" => data_out <= rom_array(23709);
		when "0101110010011110" => data_out <= rom_array(23710);
		when "0101110010011111" => data_out <= rom_array(23711);
		when "0101110010100000" => data_out <= rom_array(23712);
		when "0101110010100001" => data_out <= rom_array(23713);
		when "0101110010100010" => data_out <= rom_array(23714);
		when "0101110010100011" => data_out <= rom_array(23715);
		when "0101110010100100" => data_out <= rom_array(23716);
		when "0101110010100101" => data_out <= rom_array(23717);
		when "0101110010100110" => data_out <= rom_array(23718);
		when "0101110010100111" => data_out <= rom_array(23719);
		when "0101110010101000" => data_out <= rom_array(23720);
		when "0101110010101001" => data_out <= rom_array(23721);
		when "0101110010101010" => data_out <= rom_array(23722);
		when "0101110010101011" => data_out <= rom_array(23723);
		when "0101110010101100" => data_out <= rom_array(23724);
		when "0101110010101101" => data_out <= rom_array(23725);
		when "0101110010101110" => data_out <= rom_array(23726);
		when "0101110010101111" => data_out <= rom_array(23727);
		when "0101110010110000" => data_out <= rom_array(23728);
		when "0101110010110001" => data_out <= rom_array(23729);
		when "0101110010110010" => data_out <= rom_array(23730);
		when "0101110010110011" => data_out <= rom_array(23731);
		when "0101110010110100" => data_out <= rom_array(23732);
		when "0101110010110101" => data_out <= rom_array(23733);
		when "0101110010110110" => data_out <= rom_array(23734);
		when "0101110010110111" => data_out <= rom_array(23735);
		when "0101110010111000" => data_out <= rom_array(23736);
		when "0101110010111001" => data_out <= rom_array(23737);
		when "0101110010111010" => data_out <= rom_array(23738);
		when "0101110010111011" => data_out <= rom_array(23739);
		when "0101110010111100" => data_out <= rom_array(23740);
		when "0101110010111101" => data_out <= rom_array(23741);
		when "0101110010111110" => data_out <= rom_array(23742);
		when "0101110010111111" => data_out <= rom_array(23743);
		when "0101110011000000" => data_out <= rom_array(23744);
		when "0101110011000001" => data_out <= rom_array(23745);
		when "0101110011000010" => data_out <= rom_array(23746);
		when "0101110011000011" => data_out <= rom_array(23747);
		when "0101110011000100" => data_out <= rom_array(23748);
		when "0101110011000101" => data_out <= rom_array(23749);
		when "0101110011000110" => data_out <= rom_array(23750);
		when "0101110011000111" => data_out <= rom_array(23751);
		when "0101110011001000" => data_out <= rom_array(23752);
		when "0101110011001001" => data_out <= rom_array(23753);
		when "0101110011001010" => data_out <= rom_array(23754);
		when "0101110011001011" => data_out <= rom_array(23755);
		when "0101110011001100" => data_out <= rom_array(23756);
		when "0101110011001101" => data_out <= rom_array(23757);
		when "0101110011001110" => data_out <= rom_array(23758);
		when "0101110011001111" => data_out <= rom_array(23759);
		when "0101110011010000" => data_out <= rom_array(23760);
		when "0101110011010001" => data_out <= rom_array(23761);
		when "0101110011010010" => data_out <= rom_array(23762);
		when "0101110011010011" => data_out <= rom_array(23763);
		when "0101110011010100" => data_out <= rom_array(23764);
		when "0101110011010101" => data_out <= rom_array(23765);
		when "0101110011010110" => data_out <= rom_array(23766);
		when "0101110011010111" => data_out <= rom_array(23767);
		when "0101110011011000" => data_out <= rom_array(23768);
		when "0101110011011001" => data_out <= rom_array(23769);
		when "0101110011011010" => data_out <= rom_array(23770);
		when "0101110011011011" => data_out <= rom_array(23771);
		when "0101110011011100" => data_out <= rom_array(23772);
		when "0101110011011101" => data_out <= rom_array(23773);
		when "0101110011011110" => data_out <= rom_array(23774);
		when "0101110011011111" => data_out <= rom_array(23775);
		when "0101110011100000" => data_out <= rom_array(23776);
		when "0101110011100001" => data_out <= rom_array(23777);
		when "0101110011100010" => data_out <= rom_array(23778);
		when "0101110011100011" => data_out <= rom_array(23779);
		when "0101110011100100" => data_out <= rom_array(23780);
		when "0101110011100101" => data_out <= rom_array(23781);
		when "0101110011100110" => data_out <= rom_array(23782);
		when "0101110011100111" => data_out <= rom_array(23783);
		when "0101110011101000" => data_out <= rom_array(23784);
		when "0101110011101001" => data_out <= rom_array(23785);
		when "0101110011101010" => data_out <= rom_array(23786);
		when "0101110011101011" => data_out <= rom_array(23787);
		when "0101110011101100" => data_out <= rom_array(23788);
		when "0101110011101101" => data_out <= rom_array(23789);
		when "0101110011101110" => data_out <= rom_array(23790);
		when "0101110011101111" => data_out <= rom_array(23791);
		when "0101110011110000" => data_out <= rom_array(23792);
		when "0101110011110001" => data_out <= rom_array(23793);
		when "0101110011110010" => data_out <= rom_array(23794);
		when "0101110011110011" => data_out <= rom_array(23795);
		when "0101110011110100" => data_out <= rom_array(23796);
		when "0101110011110101" => data_out <= rom_array(23797);
		when "0101110011110110" => data_out <= rom_array(23798);
		when "0101110011110111" => data_out <= rom_array(23799);
		when "0101110011111000" => data_out <= rom_array(23800);
		when "0101110011111001" => data_out <= rom_array(23801);
		when "0101110011111010" => data_out <= rom_array(23802);
		when "0101110011111011" => data_out <= rom_array(23803);
		when "0101110011111100" => data_out <= rom_array(23804);
		when "0101110011111101" => data_out <= rom_array(23805);
		when "0101110011111110" => data_out <= rom_array(23806);
		when "0101110011111111" => data_out <= rom_array(23807);
		when "0101110100000000" => data_out <= rom_array(23808);
		when "0101110100000001" => data_out <= rom_array(23809);
		when "0101110100000010" => data_out <= rom_array(23810);
		when "0101110100000011" => data_out <= rom_array(23811);
		when "0101110100000100" => data_out <= rom_array(23812);
		when "0101110100000101" => data_out <= rom_array(23813);
		when "0101110100000110" => data_out <= rom_array(23814);
		when "0101110100000111" => data_out <= rom_array(23815);
		when "0101110100001000" => data_out <= rom_array(23816);
		when "0101110100001001" => data_out <= rom_array(23817);
		when "0101110100001010" => data_out <= rom_array(23818);
		when "0101110100001011" => data_out <= rom_array(23819);
		when "0101110100001100" => data_out <= rom_array(23820);
		when "0101110100001101" => data_out <= rom_array(23821);
		when "0101110100001110" => data_out <= rom_array(23822);
		when "0101110100001111" => data_out <= rom_array(23823);
		when "0101110100010000" => data_out <= rom_array(23824);
		when "0101110100010001" => data_out <= rom_array(23825);
		when "0101110100010010" => data_out <= rom_array(23826);
		when "0101110100010011" => data_out <= rom_array(23827);
		when "0101110100010100" => data_out <= rom_array(23828);
		when "0101110100010101" => data_out <= rom_array(23829);
		when "0101110100010110" => data_out <= rom_array(23830);
		when "0101110100010111" => data_out <= rom_array(23831);
		when "0101110100011000" => data_out <= rom_array(23832);
		when "0101110100011001" => data_out <= rom_array(23833);
		when "0101110100011010" => data_out <= rom_array(23834);
		when "0101110100011011" => data_out <= rom_array(23835);
		when "0101110100011100" => data_out <= rom_array(23836);
		when "0101110100011101" => data_out <= rom_array(23837);
		when "0101110100011110" => data_out <= rom_array(23838);
		when "0101110100011111" => data_out <= rom_array(23839);
		when "0101110100100000" => data_out <= rom_array(23840);
		when "0101110100100001" => data_out <= rom_array(23841);
		when "0101110100100010" => data_out <= rom_array(23842);
		when "0101110100100011" => data_out <= rom_array(23843);
		when "0101110100100100" => data_out <= rom_array(23844);
		when "0101110100100101" => data_out <= rom_array(23845);
		when "0101110100100110" => data_out <= rom_array(23846);
		when "0101110100100111" => data_out <= rom_array(23847);
		when "0101110100101000" => data_out <= rom_array(23848);
		when "0101110100101001" => data_out <= rom_array(23849);
		when "0101110100101010" => data_out <= rom_array(23850);
		when "0101110100101011" => data_out <= rom_array(23851);
		when "0101110100101100" => data_out <= rom_array(23852);
		when "0101110100101101" => data_out <= rom_array(23853);
		when "0101110100101110" => data_out <= rom_array(23854);
		when "0101110100101111" => data_out <= rom_array(23855);
		when "0101110100110000" => data_out <= rom_array(23856);
		when "0101110100110001" => data_out <= rom_array(23857);
		when "0101110100110010" => data_out <= rom_array(23858);
		when "0101110100110011" => data_out <= rom_array(23859);
		when "0101110100110100" => data_out <= rom_array(23860);
		when "0101110100110101" => data_out <= rom_array(23861);
		when "0101110100110110" => data_out <= rom_array(23862);
		when "0101110100110111" => data_out <= rom_array(23863);
		when "0101110100111000" => data_out <= rom_array(23864);
		when "0101110100111001" => data_out <= rom_array(23865);
		when "0101110100111010" => data_out <= rom_array(23866);
		when "0101110100111011" => data_out <= rom_array(23867);
		when "0101110100111100" => data_out <= rom_array(23868);
		when "0101110100111101" => data_out <= rom_array(23869);
		when "0101110100111110" => data_out <= rom_array(23870);
		when "0101110100111111" => data_out <= rom_array(23871);
		when "0101110101000000" => data_out <= rom_array(23872);
		when "0101110101000001" => data_out <= rom_array(23873);
		when "0101110101000010" => data_out <= rom_array(23874);
		when "0101110101000011" => data_out <= rom_array(23875);
		when "0101110101000100" => data_out <= rom_array(23876);
		when "0101110101000101" => data_out <= rom_array(23877);
		when "0101110101000110" => data_out <= rom_array(23878);
		when "0101110101000111" => data_out <= rom_array(23879);
		when "0101110101001000" => data_out <= rom_array(23880);
		when "0101110101001001" => data_out <= rom_array(23881);
		when "0101110101001010" => data_out <= rom_array(23882);
		when "0101110101001011" => data_out <= rom_array(23883);
		when "0101110101001100" => data_out <= rom_array(23884);
		when "0101110101001101" => data_out <= rom_array(23885);
		when "0101110101001110" => data_out <= rom_array(23886);
		when "0101110101001111" => data_out <= rom_array(23887);
		when "0101110101010000" => data_out <= rom_array(23888);
		when "0101110101010001" => data_out <= rom_array(23889);
		when "0101110101010010" => data_out <= rom_array(23890);
		when "0101110101010011" => data_out <= rom_array(23891);
		when "0101110101010100" => data_out <= rom_array(23892);
		when "0101110101010101" => data_out <= rom_array(23893);
		when "0101110101010110" => data_out <= rom_array(23894);
		when "0101110101010111" => data_out <= rom_array(23895);
		when "0101110101011000" => data_out <= rom_array(23896);
		when "0101110101011001" => data_out <= rom_array(23897);
		when "0101110101011010" => data_out <= rom_array(23898);
		when "0101110101011011" => data_out <= rom_array(23899);
		when "0101110101011100" => data_out <= rom_array(23900);
		when "0101110101011101" => data_out <= rom_array(23901);
		when "0101110101011110" => data_out <= rom_array(23902);
		when "0101110101011111" => data_out <= rom_array(23903);
		when "0101110101100000" => data_out <= rom_array(23904);
		when "0101110101100001" => data_out <= rom_array(23905);
		when "0101110101100010" => data_out <= rom_array(23906);
		when "0101110101100011" => data_out <= rom_array(23907);
		when "0101110101100100" => data_out <= rom_array(23908);
		when "0101110101100101" => data_out <= rom_array(23909);
		when "0101110101100110" => data_out <= rom_array(23910);
		when "0101110101100111" => data_out <= rom_array(23911);
		when "0101110101101000" => data_out <= rom_array(23912);
		when "0101110101101001" => data_out <= rom_array(23913);
		when "0101110101101010" => data_out <= rom_array(23914);
		when "0101110101101011" => data_out <= rom_array(23915);
		when "0101110101101100" => data_out <= rom_array(23916);
		when "0101110101101101" => data_out <= rom_array(23917);
		when "0101110101101110" => data_out <= rom_array(23918);
		when "0101110101101111" => data_out <= rom_array(23919);
		when "0101110101110000" => data_out <= rom_array(23920);
		when "0101110101110001" => data_out <= rom_array(23921);
		when "0101110101110010" => data_out <= rom_array(23922);
		when "0101110101110011" => data_out <= rom_array(23923);
		when "0101110101110100" => data_out <= rom_array(23924);
		when "0101110101110101" => data_out <= rom_array(23925);
		when "0101110101110110" => data_out <= rom_array(23926);
		when "0101110101110111" => data_out <= rom_array(23927);
		when "0101110101111000" => data_out <= rom_array(23928);
		when "0101110101111001" => data_out <= rom_array(23929);
		when "0101110101111010" => data_out <= rom_array(23930);
		when "0101110101111011" => data_out <= rom_array(23931);
		when "0101110101111100" => data_out <= rom_array(23932);
		when "0101110101111101" => data_out <= rom_array(23933);
		when "0101110101111110" => data_out <= rom_array(23934);
		when "0101110101111111" => data_out <= rom_array(23935);
		when "0101110110000000" => data_out <= rom_array(23936);
		when "0101110110000001" => data_out <= rom_array(23937);
		when "0101110110000010" => data_out <= rom_array(23938);
		when "0101110110000011" => data_out <= rom_array(23939);
		when "0101110110000100" => data_out <= rom_array(23940);
		when "0101110110000101" => data_out <= rom_array(23941);
		when "0101110110000110" => data_out <= rom_array(23942);
		when "0101110110000111" => data_out <= rom_array(23943);
		when "0101110110001000" => data_out <= rom_array(23944);
		when "0101110110001001" => data_out <= rom_array(23945);
		when "0101110110001010" => data_out <= rom_array(23946);
		when "0101110110001011" => data_out <= rom_array(23947);
		when "0101110110001100" => data_out <= rom_array(23948);
		when "0101110110001101" => data_out <= rom_array(23949);
		when "0101110110001110" => data_out <= rom_array(23950);
		when "0101110110001111" => data_out <= rom_array(23951);
		when "0101110110010000" => data_out <= rom_array(23952);
		when "0101110110010001" => data_out <= rom_array(23953);
		when "0101110110010010" => data_out <= rom_array(23954);
		when "0101110110010011" => data_out <= rom_array(23955);
		when "0101110110010100" => data_out <= rom_array(23956);
		when "0101110110010101" => data_out <= rom_array(23957);
		when "0101110110010110" => data_out <= rom_array(23958);
		when "0101110110010111" => data_out <= rom_array(23959);
		when "0101110110011000" => data_out <= rom_array(23960);
		when "0101110110011001" => data_out <= rom_array(23961);
		when "0101110110011010" => data_out <= rom_array(23962);
		when "0101110110011011" => data_out <= rom_array(23963);
		when "0101110110011100" => data_out <= rom_array(23964);
		when "0101110110011101" => data_out <= rom_array(23965);
		when "0101110110011110" => data_out <= rom_array(23966);
		when "0101110110011111" => data_out <= rom_array(23967);
		when "0101110110100000" => data_out <= rom_array(23968);
		when "0101110110100001" => data_out <= rom_array(23969);
		when "0101110110100010" => data_out <= rom_array(23970);
		when "0101110110100011" => data_out <= rom_array(23971);
		when "0101110110100100" => data_out <= rom_array(23972);
		when "0101110110100101" => data_out <= rom_array(23973);
		when "0101110110100110" => data_out <= rom_array(23974);
		when "0101110110100111" => data_out <= rom_array(23975);
		when "0101110110101000" => data_out <= rom_array(23976);
		when "0101110110101001" => data_out <= rom_array(23977);
		when "0101110110101010" => data_out <= rom_array(23978);
		when "0101110110101011" => data_out <= rom_array(23979);
		when "0101110110101100" => data_out <= rom_array(23980);
		when "0101110110101101" => data_out <= rom_array(23981);
		when "0101110110101110" => data_out <= rom_array(23982);
		when "0101110110101111" => data_out <= rom_array(23983);
		when "0101110110110000" => data_out <= rom_array(23984);
		when "0101110110110001" => data_out <= rom_array(23985);
		when "0101110110110010" => data_out <= rom_array(23986);
		when "0101110110110011" => data_out <= rom_array(23987);
		when "0101110110110100" => data_out <= rom_array(23988);
		when "0101110110110101" => data_out <= rom_array(23989);
		when "0101110110110110" => data_out <= rom_array(23990);
		when "0101110110110111" => data_out <= rom_array(23991);
		when "0101110110111000" => data_out <= rom_array(23992);
		when "0101110110111001" => data_out <= rom_array(23993);
		when "0101110110111010" => data_out <= rom_array(23994);
		when "0101110110111011" => data_out <= rom_array(23995);
		when "0101110110111100" => data_out <= rom_array(23996);
		when "0101110110111101" => data_out <= rom_array(23997);
		when "0101110110111110" => data_out <= rom_array(23998);
		when "0101110110111111" => data_out <= rom_array(23999);
		when "0101110111000000" => data_out <= rom_array(24000);
		when "0101110111000001" => data_out <= rom_array(24001);
		when "0101110111000010" => data_out <= rom_array(24002);
		when "0101110111000011" => data_out <= rom_array(24003);
		when "0101110111000100" => data_out <= rom_array(24004);
		when "0101110111000101" => data_out <= rom_array(24005);
		when "0101110111000110" => data_out <= rom_array(24006);
		when "0101110111000111" => data_out <= rom_array(24007);
		when "0101110111001000" => data_out <= rom_array(24008);
		when "0101110111001001" => data_out <= rom_array(24009);
		when "0101110111001010" => data_out <= rom_array(24010);
		when "0101110111001011" => data_out <= rom_array(24011);
		when "0101110111001100" => data_out <= rom_array(24012);
		when "0101110111001101" => data_out <= rom_array(24013);
		when "0101110111001110" => data_out <= rom_array(24014);
		when "0101110111001111" => data_out <= rom_array(24015);
		when "0101110111010000" => data_out <= rom_array(24016);
		when "0101110111010001" => data_out <= rom_array(24017);
		when "0101110111010010" => data_out <= rom_array(24018);
		when "0101110111010011" => data_out <= rom_array(24019);
		when "0101110111010100" => data_out <= rom_array(24020);
		when "0101110111010101" => data_out <= rom_array(24021);
		when "0101110111010110" => data_out <= rom_array(24022);
		when "0101110111010111" => data_out <= rom_array(24023);
		when "0101110111011000" => data_out <= rom_array(24024);
		when "0101110111011001" => data_out <= rom_array(24025);
		when "0101110111011010" => data_out <= rom_array(24026);
		when "0101110111011011" => data_out <= rom_array(24027);
		when "0101110111011100" => data_out <= rom_array(24028);
		when "0101110111011101" => data_out <= rom_array(24029);
		when "0101110111011110" => data_out <= rom_array(24030);
		when "0101110111011111" => data_out <= rom_array(24031);
		when "0101110111100000" => data_out <= rom_array(24032);
		when "0101110111100001" => data_out <= rom_array(24033);
		when "0101110111100010" => data_out <= rom_array(24034);
		when "0101110111100011" => data_out <= rom_array(24035);
		when "0101110111100100" => data_out <= rom_array(24036);
		when "0101110111100101" => data_out <= rom_array(24037);
		when "0101110111100110" => data_out <= rom_array(24038);
		when "0101110111100111" => data_out <= rom_array(24039);
		when "0101110111101000" => data_out <= rom_array(24040);
		when "0101110111101001" => data_out <= rom_array(24041);
		when "0101110111101010" => data_out <= rom_array(24042);
		when "0101110111101011" => data_out <= rom_array(24043);
		when "0101110111101100" => data_out <= rom_array(24044);
		when "0101110111101101" => data_out <= rom_array(24045);
		when "0101110111101110" => data_out <= rom_array(24046);
		when "0101110111101111" => data_out <= rom_array(24047);
		when "0101110111110000" => data_out <= rom_array(24048);
		when "0101110111110001" => data_out <= rom_array(24049);
		when "0101110111110010" => data_out <= rom_array(24050);
		when "0101110111110011" => data_out <= rom_array(24051);
		when "0101110111110100" => data_out <= rom_array(24052);
		when "0101110111110101" => data_out <= rom_array(24053);
		when "0101110111110110" => data_out <= rom_array(24054);
		when "0101110111110111" => data_out <= rom_array(24055);
		when "0101110111111000" => data_out <= rom_array(24056);
		when "0101110111111001" => data_out <= rom_array(24057);
		when "0101110111111010" => data_out <= rom_array(24058);
		when "0101110111111011" => data_out <= rom_array(24059);
		when "0101110111111100" => data_out <= rom_array(24060);
		when "0101110111111101" => data_out <= rom_array(24061);
		when "0101110111111110" => data_out <= rom_array(24062);
		when "0101110111111111" => data_out <= rom_array(24063);
		when "0101111000000000" => data_out <= rom_array(24064);
		when "0101111000000001" => data_out <= rom_array(24065);
		when "0101111000000010" => data_out <= rom_array(24066);
		when "0101111000000011" => data_out <= rom_array(24067);
		when "0101111000000100" => data_out <= rom_array(24068);
		when "0101111000000101" => data_out <= rom_array(24069);
		when "0101111000000110" => data_out <= rom_array(24070);
		when "0101111000000111" => data_out <= rom_array(24071);
		when "0101111000001000" => data_out <= rom_array(24072);
		when "0101111000001001" => data_out <= rom_array(24073);
		when "0101111000001010" => data_out <= rom_array(24074);
		when "0101111000001011" => data_out <= rom_array(24075);
		when "0101111000001100" => data_out <= rom_array(24076);
		when "0101111000001101" => data_out <= rom_array(24077);
		when "0101111000001110" => data_out <= rom_array(24078);
		when "0101111000001111" => data_out <= rom_array(24079);
		when "0101111000010000" => data_out <= rom_array(24080);
		when "0101111000010001" => data_out <= rom_array(24081);
		when "0101111000010010" => data_out <= rom_array(24082);
		when "0101111000010011" => data_out <= rom_array(24083);
		when "0101111000010100" => data_out <= rom_array(24084);
		when "0101111000010101" => data_out <= rom_array(24085);
		when "0101111000010110" => data_out <= rom_array(24086);
		when "0101111000010111" => data_out <= rom_array(24087);
		when "0101111000011000" => data_out <= rom_array(24088);
		when "0101111000011001" => data_out <= rom_array(24089);
		when "0101111000011010" => data_out <= rom_array(24090);
		when "0101111000011011" => data_out <= rom_array(24091);
		when "0101111000011100" => data_out <= rom_array(24092);
		when "0101111000011101" => data_out <= rom_array(24093);
		when "0101111000011110" => data_out <= rom_array(24094);
		when "0101111000011111" => data_out <= rom_array(24095);
		when "0101111000100000" => data_out <= rom_array(24096);
		when "0101111000100001" => data_out <= rom_array(24097);
		when "0101111000100010" => data_out <= rom_array(24098);
		when "0101111000100011" => data_out <= rom_array(24099);
		when "0101111000100100" => data_out <= rom_array(24100);
		when "0101111000100101" => data_out <= rom_array(24101);
		when "0101111000100110" => data_out <= rom_array(24102);
		when "0101111000100111" => data_out <= rom_array(24103);
		when "0101111000101000" => data_out <= rom_array(24104);
		when "0101111000101001" => data_out <= rom_array(24105);
		when "0101111000101010" => data_out <= rom_array(24106);
		when "0101111000101011" => data_out <= rom_array(24107);
		when "0101111000101100" => data_out <= rom_array(24108);
		when "0101111000101101" => data_out <= rom_array(24109);
		when "0101111000101110" => data_out <= rom_array(24110);
		when "0101111000101111" => data_out <= rom_array(24111);
		when "0101111000110000" => data_out <= rom_array(24112);
		when "0101111000110001" => data_out <= rom_array(24113);
		when "0101111000110010" => data_out <= rom_array(24114);
		when "0101111000110011" => data_out <= rom_array(24115);
		when "0101111000110100" => data_out <= rom_array(24116);
		when "0101111000110101" => data_out <= rom_array(24117);
		when "0101111000110110" => data_out <= rom_array(24118);
		when "0101111000110111" => data_out <= rom_array(24119);
		when "0101111000111000" => data_out <= rom_array(24120);
		when "0101111000111001" => data_out <= rom_array(24121);
		when "0101111000111010" => data_out <= rom_array(24122);
		when "0101111000111011" => data_out <= rom_array(24123);
		when "0101111000111100" => data_out <= rom_array(24124);
		when "0101111000111101" => data_out <= rom_array(24125);
		when "0101111000111110" => data_out <= rom_array(24126);
		when "0101111000111111" => data_out <= rom_array(24127);
		when "0101111001000000" => data_out <= rom_array(24128);
		when "0101111001000001" => data_out <= rom_array(24129);
		when "0101111001000010" => data_out <= rom_array(24130);
		when "0101111001000011" => data_out <= rom_array(24131);
		when "0101111001000100" => data_out <= rom_array(24132);
		when "0101111001000101" => data_out <= rom_array(24133);
		when "0101111001000110" => data_out <= rom_array(24134);
		when "0101111001000111" => data_out <= rom_array(24135);
		when "0101111001001000" => data_out <= rom_array(24136);
		when "0101111001001001" => data_out <= rom_array(24137);
		when "0101111001001010" => data_out <= rom_array(24138);
		when "0101111001001011" => data_out <= rom_array(24139);
		when "0101111001001100" => data_out <= rom_array(24140);
		when "0101111001001101" => data_out <= rom_array(24141);
		when "0101111001001110" => data_out <= rom_array(24142);
		when "0101111001001111" => data_out <= rom_array(24143);
		when "0101111001010000" => data_out <= rom_array(24144);
		when "0101111001010001" => data_out <= rom_array(24145);
		when "0101111001010010" => data_out <= rom_array(24146);
		when "0101111001010011" => data_out <= rom_array(24147);
		when "0101111001010100" => data_out <= rom_array(24148);
		when "0101111001010101" => data_out <= rom_array(24149);
		when "0101111001010110" => data_out <= rom_array(24150);
		when "0101111001010111" => data_out <= rom_array(24151);
		when "0101111001011000" => data_out <= rom_array(24152);
		when "0101111001011001" => data_out <= rom_array(24153);
		when "0101111001011010" => data_out <= rom_array(24154);
		when "0101111001011011" => data_out <= rom_array(24155);
		when "0101111001011100" => data_out <= rom_array(24156);
		when "0101111001011101" => data_out <= rom_array(24157);
		when "0101111001011110" => data_out <= rom_array(24158);
		when "0101111001011111" => data_out <= rom_array(24159);
		when "0101111001100000" => data_out <= rom_array(24160);
		when "0101111001100001" => data_out <= rom_array(24161);
		when "0101111001100010" => data_out <= rom_array(24162);
		when "0101111001100011" => data_out <= rom_array(24163);
		when "0101111001100100" => data_out <= rom_array(24164);
		when "0101111001100101" => data_out <= rom_array(24165);
		when "0101111001100110" => data_out <= rom_array(24166);
		when "0101111001100111" => data_out <= rom_array(24167);
		when "0101111001101000" => data_out <= rom_array(24168);
		when "0101111001101001" => data_out <= rom_array(24169);
		when "0101111001101010" => data_out <= rom_array(24170);
		when "0101111001101011" => data_out <= rom_array(24171);
		when "0101111001101100" => data_out <= rom_array(24172);
		when "0101111001101101" => data_out <= rom_array(24173);
		when "0101111001101110" => data_out <= rom_array(24174);
		when "0101111001101111" => data_out <= rom_array(24175);
		when "0101111001110000" => data_out <= rom_array(24176);
		when "0101111001110001" => data_out <= rom_array(24177);
		when "0101111001110010" => data_out <= rom_array(24178);
		when "0101111001110011" => data_out <= rom_array(24179);
		when "0101111001110100" => data_out <= rom_array(24180);
		when "0101111001110101" => data_out <= rom_array(24181);
		when "0101111001110110" => data_out <= rom_array(24182);
		when "0101111001110111" => data_out <= rom_array(24183);
		when "0101111001111000" => data_out <= rom_array(24184);
		when "0101111001111001" => data_out <= rom_array(24185);
		when "0101111001111010" => data_out <= rom_array(24186);
		when "0101111001111011" => data_out <= rom_array(24187);
		when "0101111001111100" => data_out <= rom_array(24188);
		when "0101111001111101" => data_out <= rom_array(24189);
		when "0101111001111110" => data_out <= rom_array(24190);
		when "0101111001111111" => data_out <= rom_array(24191);
		when "0101111010000000" => data_out <= rom_array(24192);
		when "0101111010000001" => data_out <= rom_array(24193);
		when "0101111010000010" => data_out <= rom_array(24194);
		when "0101111010000011" => data_out <= rom_array(24195);
		when "0101111010000100" => data_out <= rom_array(24196);
		when "0101111010000101" => data_out <= rom_array(24197);
		when "0101111010000110" => data_out <= rom_array(24198);
		when "0101111010000111" => data_out <= rom_array(24199);
		when "0101111010001000" => data_out <= rom_array(24200);
		when "0101111010001001" => data_out <= rom_array(24201);
		when "0101111010001010" => data_out <= rom_array(24202);
		when "0101111010001011" => data_out <= rom_array(24203);
		when "0101111010001100" => data_out <= rom_array(24204);
		when "0101111010001101" => data_out <= rom_array(24205);
		when "0101111010001110" => data_out <= rom_array(24206);
		when "0101111010001111" => data_out <= rom_array(24207);
		when "0101111010010000" => data_out <= rom_array(24208);
		when "0101111010010001" => data_out <= rom_array(24209);
		when "0101111010010010" => data_out <= rom_array(24210);
		when "0101111010010011" => data_out <= rom_array(24211);
		when "0101111010010100" => data_out <= rom_array(24212);
		when "0101111010010101" => data_out <= rom_array(24213);
		when "0101111010010110" => data_out <= rom_array(24214);
		when "0101111010010111" => data_out <= rom_array(24215);
		when "0101111010011000" => data_out <= rom_array(24216);
		when "0101111010011001" => data_out <= rom_array(24217);
		when "0101111010011010" => data_out <= rom_array(24218);
		when "0101111010011011" => data_out <= rom_array(24219);
		when "0101111010011100" => data_out <= rom_array(24220);
		when "0101111010011101" => data_out <= rom_array(24221);
		when "0101111010011110" => data_out <= rom_array(24222);
		when "0101111010011111" => data_out <= rom_array(24223);
		when "0101111010100000" => data_out <= rom_array(24224);
		when "0101111010100001" => data_out <= rom_array(24225);
		when "0101111010100010" => data_out <= rom_array(24226);
		when "0101111010100011" => data_out <= rom_array(24227);
		when "0101111010100100" => data_out <= rom_array(24228);
		when "0101111010100101" => data_out <= rom_array(24229);
		when "0101111010100110" => data_out <= rom_array(24230);
		when "0101111010100111" => data_out <= rom_array(24231);
		when "0101111010101000" => data_out <= rom_array(24232);
		when "0101111010101001" => data_out <= rom_array(24233);
		when "0101111010101010" => data_out <= rom_array(24234);
		when "0101111010101011" => data_out <= rom_array(24235);
		when "0101111010101100" => data_out <= rom_array(24236);
		when "0101111010101101" => data_out <= rom_array(24237);
		when "0101111010101110" => data_out <= rom_array(24238);
		when "0101111010101111" => data_out <= rom_array(24239);
		when "0101111010110000" => data_out <= rom_array(24240);
		when "0101111010110001" => data_out <= rom_array(24241);
		when "0101111010110010" => data_out <= rom_array(24242);
		when "0101111010110011" => data_out <= rom_array(24243);
		when "0101111010110100" => data_out <= rom_array(24244);
		when "0101111010110101" => data_out <= rom_array(24245);
		when "0101111010110110" => data_out <= rom_array(24246);
		when "0101111010110111" => data_out <= rom_array(24247);
		when "0101111010111000" => data_out <= rom_array(24248);
		when "0101111010111001" => data_out <= rom_array(24249);
		when "0101111010111010" => data_out <= rom_array(24250);
		when "0101111010111011" => data_out <= rom_array(24251);
		when "0101111010111100" => data_out <= rom_array(24252);
		when "0101111010111101" => data_out <= rom_array(24253);
		when "0101111010111110" => data_out <= rom_array(24254);
		when "0101111010111111" => data_out <= rom_array(24255);
		when "0101111011000000" => data_out <= rom_array(24256);
		when "0101111011000001" => data_out <= rom_array(24257);
		when "0101111011000010" => data_out <= rom_array(24258);
		when "0101111011000011" => data_out <= rom_array(24259);
		when "0101111011000100" => data_out <= rom_array(24260);
		when "0101111011000101" => data_out <= rom_array(24261);
		when "0101111011000110" => data_out <= rom_array(24262);
		when "0101111011000111" => data_out <= rom_array(24263);
		when "0101111011001000" => data_out <= rom_array(24264);
		when "0101111011001001" => data_out <= rom_array(24265);
		when "0101111011001010" => data_out <= rom_array(24266);
		when "0101111011001011" => data_out <= rom_array(24267);
		when "0101111011001100" => data_out <= rom_array(24268);
		when "0101111011001101" => data_out <= rom_array(24269);
		when "0101111011001110" => data_out <= rom_array(24270);
		when "0101111011001111" => data_out <= rom_array(24271);
		when "0101111011010000" => data_out <= rom_array(24272);
		when "0101111011010001" => data_out <= rom_array(24273);
		when "0101111011010010" => data_out <= rom_array(24274);
		when "0101111011010011" => data_out <= rom_array(24275);
		when "0101111011010100" => data_out <= rom_array(24276);
		when "0101111011010101" => data_out <= rom_array(24277);
		when "0101111011010110" => data_out <= rom_array(24278);
		when "0101111011010111" => data_out <= rom_array(24279);
		when "0101111011011000" => data_out <= rom_array(24280);
		when "0101111011011001" => data_out <= rom_array(24281);
		when "0101111011011010" => data_out <= rom_array(24282);
		when "0101111011011011" => data_out <= rom_array(24283);
		when "0101111011011100" => data_out <= rom_array(24284);
		when "0101111011011101" => data_out <= rom_array(24285);
		when "0101111011011110" => data_out <= rom_array(24286);
		when "0101111011011111" => data_out <= rom_array(24287);
		when "0101111011100000" => data_out <= rom_array(24288);
		when "0101111011100001" => data_out <= rom_array(24289);
		when "0101111011100010" => data_out <= rom_array(24290);
		when "0101111011100011" => data_out <= rom_array(24291);
		when "0101111011100100" => data_out <= rom_array(24292);
		when "0101111011100101" => data_out <= rom_array(24293);
		when "0101111011100110" => data_out <= rom_array(24294);
		when "0101111011100111" => data_out <= rom_array(24295);
		when "0101111011101000" => data_out <= rom_array(24296);
		when "0101111011101001" => data_out <= rom_array(24297);
		when "0101111011101010" => data_out <= rom_array(24298);
		when "0101111011101011" => data_out <= rom_array(24299);
		when "0101111011101100" => data_out <= rom_array(24300);
		when "0101111011101101" => data_out <= rom_array(24301);
		when "0101111011101110" => data_out <= rom_array(24302);
		when "0101111011101111" => data_out <= rom_array(24303);
		when "0101111011110000" => data_out <= rom_array(24304);
		when "0101111011110001" => data_out <= rom_array(24305);
		when "0101111011110010" => data_out <= rom_array(24306);
		when "0101111011110011" => data_out <= rom_array(24307);
		when "0101111011110100" => data_out <= rom_array(24308);
		when "0101111011110101" => data_out <= rom_array(24309);
		when "0101111011110110" => data_out <= rom_array(24310);
		when "0101111011110111" => data_out <= rom_array(24311);
		when "0101111011111000" => data_out <= rom_array(24312);
		when "0101111011111001" => data_out <= rom_array(24313);
		when "0101111011111010" => data_out <= rom_array(24314);
		when "0101111011111011" => data_out <= rom_array(24315);
		when "0101111011111100" => data_out <= rom_array(24316);
		when "0101111011111101" => data_out <= rom_array(24317);
		when "0101111011111110" => data_out <= rom_array(24318);
		when "0101111011111111" => data_out <= rom_array(24319);
		when "0101111100000000" => data_out <= rom_array(24320);
		when "0101111100000001" => data_out <= rom_array(24321);
		when "0101111100000010" => data_out <= rom_array(24322);
		when "0101111100000011" => data_out <= rom_array(24323);
		when "0101111100000100" => data_out <= rom_array(24324);
		when "0101111100000101" => data_out <= rom_array(24325);
		when "0101111100000110" => data_out <= rom_array(24326);
		when "0101111100000111" => data_out <= rom_array(24327);
		when "0101111100001000" => data_out <= rom_array(24328);
		when "0101111100001001" => data_out <= rom_array(24329);
		when "0101111100001010" => data_out <= rom_array(24330);
		when "0101111100001011" => data_out <= rom_array(24331);
		when "0101111100001100" => data_out <= rom_array(24332);
		when "0101111100001101" => data_out <= rom_array(24333);
		when "0101111100001110" => data_out <= rom_array(24334);
		when "0101111100001111" => data_out <= rom_array(24335);
		when "0101111100010000" => data_out <= rom_array(24336);
		when "0101111100010001" => data_out <= rom_array(24337);
		when "0101111100010010" => data_out <= rom_array(24338);
		when "0101111100010011" => data_out <= rom_array(24339);
		when "0101111100010100" => data_out <= rom_array(24340);
		when "0101111100010101" => data_out <= rom_array(24341);
		when "0101111100010110" => data_out <= rom_array(24342);
		when "0101111100010111" => data_out <= rom_array(24343);
		when "0101111100011000" => data_out <= rom_array(24344);
		when "0101111100011001" => data_out <= rom_array(24345);
		when "0101111100011010" => data_out <= rom_array(24346);
		when "0101111100011011" => data_out <= rom_array(24347);
		when "0101111100011100" => data_out <= rom_array(24348);
		when "0101111100011101" => data_out <= rom_array(24349);
		when "0101111100011110" => data_out <= rom_array(24350);
		when "0101111100011111" => data_out <= rom_array(24351);
		when "0101111100100000" => data_out <= rom_array(24352);
		when "0101111100100001" => data_out <= rom_array(24353);
		when "0101111100100010" => data_out <= rom_array(24354);
		when "0101111100100011" => data_out <= rom_array(24355);
		when "0101111100100100" => data_out <= rom_array(24356);
		when "0101111100100101" => data_out <= rom_array(24357);
		when "0101111100100110" => data_out <= rom_array(24358);
		when "0101111100100111" => data_out <= rom_array(24359);
		when "0101111100101000" => data_out <= rom_array(24360);
		when "0101111100101001" => data_out <= rom_array(24361);
		when "0101111100101010" => data_out <= rom_array(24362);
		when "0101111100101011" => data_out <= rom_array(24363);
		when "0101111100101100" => data_out <= rom_array(24364);
		when "0101111100101101" => data_out <= rom_array(24365);
		when "0101111100101110" => data_out <= rom_array(24366);
		when "0101111100101111" => data_out <= rom_array(24367);
		when "0101111100110000" => data_out <= rom_array(24368);
		when "0101111100110001" => data_out <= rom_array(24369);
		when "0101111100110010" => data_out <= rom_array(24370);
		when "0101111100110011" => data_out <= rom_array(24371);
		when "0101111100110100" => data_out <= rom_array(24372);
		when "0101111100110101" => data_out <= rom_array(24373);
		when "0101111100110110" => data_out <= rom_array(24374);
		when "0101111100110111" => data_out <= rom_array(24375);
		when "0101111100111000" => data_out <= rom_array(24376);
		when "0101111100111001" => data_out <= rom_array(24377);
		when "0101111100111010" => data_out <= rom_array(24378);
		when "0101111100111011" => data_out <= rom_array(24379);
		when "0101111100111100" => data_out <= rom_array(24380);
		when "0101111100111101" => data_out <= rom_array(24381);
		when "0101111100111110" => data_out <= rom_array(24382);
		when "0101111100111111" => data_out <= rom_array(24383);
		when "0101111101000000" => data_out <= rom_array(24384);
		when "0101111101000001" => data_out <= rom_array(24385);
		when "0101111101000010" => data_out <= rom_array(24386);
		when "0101111101000011" => data_out <= rom_array(24387);
		when "0101111101000100" => data_out <= rom_array(24388);
		when "0101111101000101" => data_out <= rom_array(24389);
		when "0101111101000110" => data_out <= rom_array(24390);
		when "0101111101000111" => data_out <= rom_array(24391);
		when "0101111101001000" => data_out <= rom_array(24392);
		when "0101111101001001" => data_out <= rom_array(24393);
		when "0101111101001010" => data_out <= rom_array(24394);
		when "0101111101001011" => data_out <= rom_array(24395);
		when "0101111101001100" => data_out <= rom_array(24396);
		when "0101111101001101" => data_out <= rom_array(24397);
		when "0101111101001110" => data_out <= rom_array(24398);
		when "0101111101001111" => data_out <= rom_array(24399);
		when "0101111101010000" => data_out <= rom_array(24400);
		when "0101111101010001" => data_out <= rom_array(24401);
		when "0101111101010010" => data_out <= rom_array(24402);
		when "0101111101010011" => data_out <= rom_array(24403);
		when "0101111101010100" => data_out <= rom_array(24404);
		when "0101111101010101" => data_out <= rom_array(24405);
		when "0101111101010110" => data_out <= rom_array(24406);
		when "0101111101010111" => data_out <= rom_array(24407);
		when "0101111101011000" => data_out <= rom_array(24408);
		when "0101111101011001" => data_out <= rom_array(24409);
		when "0101111101011010" => data_out <= rom_array(24410);
		when "0101111101011011" => data_out <= rom_array(24411);
		when "0101111101011100" => data_out <= rom_array(24412);
		when "0101111101011101" => data_out <= rom_array(24413);
		when "0101111101011110" => data_out <= rom_array(24414);
		when "0101111101011111" => data_out <= rom_array(24415);
		when "0101111101100000" => data_out <= rom_array(24416);
		when "0101111101100001" => data_out <= rom_array(24417);
		when "0101111101100010" => data_out <= rom_array(24418);
		when "0101111101100011" => data_out <= rom_array(24419);
		when "0101111101100100" => data_out <= rom_array(24420);
		when "0101111101100101" => data_out <= rom_array(24421);
		when "0101111101100110" => data_out <= rom_array(24422);
		when "0101111101100111" => data_out <= rom_array(24423);
		when "0101111101101000" => data_out <= rom_array(24424);
		when "0101111101101001" => data_out <= rom_array(24425);
		when "0101111101101010" => data_out <= rom_array(24426);
		when "0101111101101011" => data_out <= rom_array(24427);
		when "0101111101101100" => data_out <= rom_array(24428);
		when "0101111101101101" => data_out <= rom_array(24429);
		when "0101111101101110" => data_out <= rom_array(24430);
		when "0101111101101111" => data_out <= rom_array(24431);
		when "0101111101110000" => data_out <= rom_array(24432);
		when "0101111101110001" => data_out <= rom_array(24433);
		when "0101111101110010" => data_out <= rom_array(24434);
		when "0101111101110011" => data_out <= rom_array(24435);
		when "0101111101110100" => data_out <= rom_array(24436);
		when "0101111101110101" => data_out <= rom_array(24437);
		when "0101111101110110" => data_out <= rom_array(24438);
		when "0101111101110111" => data_out <= rom_array(24439);
		when "0101111101111000" => data_out <= rom_array(24440);
		when "0101111101111001" => data_out <= rom_array(24441);
		when "0101111101111010" => data_out <= rom_array(24442);
		when "0101111101111011" => data_out <= rom_array(24443);
		when "0101111101111100" => data_out <= rom_array(24444);
		when "0101111101111101" => data_out <= rom_array(24445);
		when "0101111101111110" => data_out <= rom_array(24446);
		when "0101111101111111" => data_out <= rom_array(24447);
		when "0101111110000000" => data_out <= rom_array(24448);
		when "0101111110000001" => data_out <= rom_array(24449);
		when "0101111110000010" => data_out <= rom_array(24450);
		when "0101111110000011" => data_out <= rom_array(24451);
		when "0101111110000100" => data_out <= rom_array(24452);
		when "0101111110000101" => data_out <= rom_array(24453);
		when "0101111110000110" => data_out <= rom_array(24454);
		when "0101111110000111" => data_out <= rom_array(24455);
		when "0101111110001000" => data_out <= rom_array(24456);
		when "0101111110001001" => data_out <= rom_array(24457);
		when "0101111110001010" => data_out <= rom_array(24458);
		when "0101111110001011" => data_out <= rom_array(24459);
		when "0101111110001100" => data_out <= rom_array(24460);
		when "0101111110001101" => data_out <= rom_array(24461);
		when "0101111110001110" => data_out <= rom_array(24462);
		when "0101111110001111" => data_out <= rom_array(24463);
		when "0101111110010000" => data_out <= rom_array(24464);
		when "0101111110010001" => data_out <= rom_array(24465);
		when "0101111110010010" => data_out <= rom_array(24466);
		when "0101111110010011" => data_out <= rom_array(24467);
		when "0101111110010100" => data_out <= rom_array(24468);
		when "0101111110010101" => data_out <= rom_array(24469);
		when "0101111110010110" => data_out <= rom_array(24470);
		when "0101111110010111" => data_out <= rom_array(24471);
		when "0101111110011000" => data_out <= rom_array(24472);
		when "0101111110011001" => data_out <= rom_array(24473);
		when "0101111110011010" => data_out <= rom_array(24474);
		when "0101111110011011" => data_out <= rom_array(24475);
		when "0101111110011100" => data_out <= rom_array(24476);
		when "0101111110011101" => data_out <= rom_array(24477);
		when "0101111110011110" => data_out <= rom_array(24478);
		when "0101111110011111" => data_out <= rom_array(24479);
		when "0101111110100000" => data_out <= rom_array(24480);
		when "0101111110100001" => data_out <= rom_array(24481);
		when "0101111110100010" => data_out <= rom_array(24482);
		when "0101111110100011" => data_out <= rom_array(24483);
		when "0101111110100100" => data_out <= rom_array(24484);
		when "0101111110100101" => data_out <= rom_array(24485);
		when "0101111110100110" => data_out <= rom_array(24486);
		when "0101111110100111" => data_out <= rom_array(24487);
		when "0101111110101000" => data_out <= rom_array(24488);
		when "0101111110101001" => data_out <= rom_array(24489);
		when "0101111110101010" => data_out <= rom_array(24490);
		when "0101111110101011" => data_out <= rom_array(24491);
		when "0101111110101100" => data_out <= rom_array(24492);
		when "0101111110101101" => data_out <= rom_array(24493);
		when "0101111110101110" => data_out <= rom_array(24494);
		when "0101111110101111" => data_out <= rom_array(24495);
		when "0101111110110000" => data_out <= rom_array(24496);
		when "0101111110110001" => data_out <= rom_array(24497);
		when "0101111110110010" => data_out <= rom_array(24498);
		when "0101111110110011" => data_out <= rom_array(24499);
		when "0101111110110100" => data_out <= rom_array(24500);
		when "0101111110110101" => data_out <= rom_array(24501);
		when "0101111110110110" => data_out <= rom_array(24502);
		when "0101111110110111" => data_out <= rom_array(24503);
		when "0101111110111000" => data_out <= rom_array(24504);
		when "0101111110111001" => data_out <= rom_array(24505);
		when "0101111110111010" => data_out <= rom_array(24506);
		when "0101111110111011" => data_out <= rom_array(24507);
		when "0101111110111100" => data_out <= rom_array(24508);
		when "0101111110111101" => data_out <= rom_array(24509);
		when "0101111110111110" => data_out <= rom_array(24510);
		when "0101111110111111" => data_out <= rom_array(24511);
		when "0101111111000000" => data_out <= rom_array(24512);
		when "0101111111000001" => data_out <= rom_array(24513);
		when "0101111111000010" => data_out <= rom_array(24514);
		when "0101111111000011" => data_out <= rom_array(24515);
		when "0101111111000100" => data_out <= rom_array(24516);
		when "0101111111000101" => data_out <= rom_array(24517);
		when "0101111111000110" => data_out <= rom_array(24518);
		when "0101111111000111" => data_out <= rom_array(24519);
		when "0101111111001000" => data_out <= rom_array(24520);
		when "0101111111001001" => data_out <= rom_array(24521);
		when "0101111111001010" => data_out <= rom_array(24522);
		when "0101111111001011" => data_out <= rom_array(24523);
		when "0101111111001100" => data_out <= rom_array(24524);
		when "0101111111001101" => data_out <= rom_array(24525);
		when "0101111111001110" => data_out <= rom_array(24526);
		when "0101111111001111" => data_out <= rom_array(24527);
		when "0101111111010000" => data_out <= rom_array(24528);
		when "0101111111010001" => data_out <= rom_array(24529);
		when "0101111111010010" => data_out <= rom_array(24530);
		when "0101111111010011" => data_out <= rom_array(24531);
		when "0101111111010100" => data_out <= rom_array(24532);
		when "0101111111010101" => data_out <= rom_array(24533);
		when "0101111111010110" => data_out <= rom_array(24534);
		when "0101111111010111" => data_out <= rom_array(24535);
		when "0101111111011000" => data_out <= rom_array(24536);
		when "0101111111011001" => data_out <= rom_array(24537);
		when "0101111111011010" => data_out <= rom_array(24538);
		when "0101111111011011" => data_out <= rom_array(24539);
		when "0101111111011100" => data_out <= rom_array(24540);
		when "0101111111011101" => data_out <= rom_array(24541);
		when "0101111111011110" => data_out <= rom_array(24542);
		when "0101111111011111" => data_out <= rom_array(24543);
		when "0101111111100000" => data_out <= rom_array(24544);
		when "0101111111100001" => data_out <= rom_array(24545);
		when "0101111111100010" => data_out <= rom_array(24546);
		when "0101111111100011" => data_out <= rom_array(24547);
		when "0101111111100100" => data_out <= rom_array(24548);
		when "0101111111100101" => data_out <= rom_array(24549);
		when "0101111111100110" => data_out <= rom_array(24550);
		when "0101111111100111" => data_out <= rom_array(24551);
		when "0101111111101000" => data_out <= rom_array(24552);
		when "0101111111101001" => data_out <= rom_array(24553);
		when "0101111111101010" => data_out <= rom_array(24554);
		when "0101111111101011" => data_out <= rom_array(24555);
		when "0101111111101100" => data_out <= rom_array(24556);
		when "0101111111101101" => data_out <= rom_array(24557);
		when "0101111111101110" => data_out <= rom_array(24558);
		when "0101111111101111" => data_out <= rom_array(24559);
		when "0101111111110000" => data_out <= rom_array(24560);
		when "0101111111110001" => data_out <= rom_array(24561);
		when "0101111111110010" => data_out <= rom_array(24562);
		when "0101111111110011" => data_out <= rom_array(24563);
		when "0101111111110100" => data_out <= rom_array(24564);
		when "0101111111110101" => data_out <= rom_array(24565);
		when "0101111111110110" => data_out <= rom_array(24566);
		when "0101111111110111" => data_out <= rom_array(24567);
		when "0101111111111000" => data_out <= rom_array(24568);
		when "0101111111111001" => data_out <= rom_array(24569);
		when "0101111111111010" => data_out <= rom_array(24570);
		when "0101111111111011" => data_out <= rom_array(24571);
		when "0101111111111100" => data_out <= rom_array(24572);
		when "0101111111111101" => data_out <= rom_array(24573);
		when "0101111111111110" => data_out <= rom_array(24574);
		when "0101111111111111" => data_out <= rom_array(24575);
		when "0110000000000000" => data_out <= rom_array(24576);
		when "0110000000000001" => data_out <= rom_array(24577);
		when "0110000000000010" => data_out <= rom_array(24578);
		when "0110000000000011" => data_out <= rom_array(24579);
		when "0110000000000100" => data_out <= rom_array(24580);
		when "0110000000000101" => data_out <= rom_array(24581);
		when "0110000000000110" => data_out <= rom_array(24582);
		when "0110000000000111" => data_out <= rom_array(24583);
		when "0110000000001000" => data_out <= rom_array(24584);
		when "0110000000001001" => data_out <= rom_array(24585);
		when "0110000000001010" => data_out <= rom_array(24586);
		when "0110000000001011" => data_out <= rom_array(24587);
		when "0110000000001100" => data_out <= rom_array(24588);
		when "0110000000001101" => data_out <= rom_array(24589);
		when "0110000000001110" => data_out <= rom_array(24590);
		when "0110000000001111" => data_out <= rom_array(24591);
		when "0110000000010000" => data_out <= rom_array(24592);
		when "0110000000010001" => data_out <= rom_array(24593);
		when "0110000000010010" => data_out <= rom_array(24594);
		when "0110000000010011" => data_out <= rom_array(24595);
		when "0110000000010100" => data_out <= rom_array(24596);
		when "0110000000010101" => data_out <= rom_array(24597);
		when "0110000000010110" => data_out <= rom_array(24598);
		when "0110000000010111" => data_out <= rom_array(24599);
		when "0110000000011000" => data_out <= rom_array(24600);
		when "0110000000011001" => data_out <= rom_array(24601);
		when "0110000000011010" => data_out <= rom_array(24602);
		when "0110000000011011" => data_out <= rom_array(24603);
		when "0110000000011100" => data_out <= rom_array(24604);
		when "0110000000011101" => data_out <= rom_array(24605);
		when "0110000000011110" => data_out <= rom_array(24606);
		when "0110000000011111" => data_out <= rom_array(24607);
		when "0110000000100000" => data_out <= rom_array(24608);
		when "0110000000100001" => data_out <= rom_array(24609);
		when "0110000000100010" => data_out <= rom_array(24610);
		when "0110000000100011" => data_out <= rom_array(24611);
		when "0110000000100100" => data_out <= rom_array(24612);
		when "0110000000100101" => data_out <= rom_array(24613);
		when "0110000000100110" => data_out <= rom_array(24614);
		when "0110000000100111" => data_out <= rom_array(24615);
		when "0110000000101000" => data_out <= rom_array(24616);
		when "0110000000101001" => data_out <= rom_array(24617);
		when "0110000000101010" => data_out <= rom_array(24618);
		when "0110000000101011" => data_out <= rom_array(24619);
		when "0110000000101100" => data_out <= rom_array(24620);
		when "0110000000101101" => data_out <= rom_array(24621);
		when "0110000000101110" => data_out <= rom_array(24622);
		when "0110000000101111" => data_out <= rom_array(24623);
		when "0110000000110000" => data_out <= rom_array(24624);
		when "0110000000110001" => data_out <= rom_array(24625);
		when "0110000000110010" => data_out <= rom_array(24626);
		when "0110000000110011" => data_out <= rom_array(24627);
		when "0110000000110100" => data_out <= rom_array(24628);
		when "0110000000110101" => data_out <= rom_array(24629);
		when "0110000000110110" => data_out <= rom_array(24630);
		when "0110000000110111" => data_out <= rom_array(24631);
		when "0110000000111000" => data_out <= rom_array(24632);
		when "0110000000111001" => data_out <= rom_array(24633);
		when "0110000000111010" => data_out <= rom_array(24634);
		when "0110000000111011" => data_out <= rom_array(24635);
		when "0110000000111100" => data_out <= rom_array(24636);
		when "0110000000111101" => data_out <= rom_array(24637);
		when "0110000000111110" => data_out <= rom_array(24638);
		when "0110000000111111" => data_out <= rom_array(24639);
		when "0110000001000000" => data_out <= rom_array(24640);
		when "0110000001000001" => data_out <= rom_array(24641);
		when "0110000001000010" => data_out <= rom_array(24642);
		when "0110000001000011" => data_out <= rom_array(24643);
		when "0110000001000100" => data_out <= rom_array(24644);
		when "0110000001000101" => data_out <= rom_array(24645);
		when "0110000001000110" => data_out <= rom_array(24646);
		when "0110000001000111" => data_out <= rom_array(24647);
		when "0110000001001000" => data_out <= rom_array(24648);
		when "0110000001001001" => data_out <= rom_array(24649);
		when "0110000001001010" => data_out <= rom_array(24650);
		when "0110000001001011" => data_out <= rom_array(24651);
		when "0110000001001100" => data_out <= rom_array(24652);
		when "0110000001001101" => data_out <= rom_array(24653);
		when "0110000001001110" => data_out <= rom_array(24654);
		when "0110000001001111" => data_out <= rom_array(24655);
		when "0110000001010000" => data_out <= rom_array(24656);
		when "0110000001010001" => data_out <= rom_array(24657);
		when "0110000001010010" => data_out <= rom_array(24658);
		when "0110000001010011" => data_out <= rom_array(24659);
		when "0110000001010100" => data_out <= rom_array(24660);
		when "0110000001010101" => data_out <= rom_array(24661);
		when "0110000001010110" => data_out <= rom_array(24662);
		when "0110000001010111" => data_out <= rom_array(24663);
		when "0110000001011000" => data_out <= rom_array(24664);
		when "0110000001011001" => data_out <= rom_array(24665);
		when "0110000001011010" => data_out <= rom_array(24666);
		when "0110000001011011" => data_out <= rom_array(24667);
		when "0110000001011100" => data_out <= rom_array(24668);
		when "0110000001011101" => data_out <= rom_array(24669);
		when "0110000001011110" => data_out <= rom_array(24670);
		when "0110000001011111" => data_out <= rom_array(24671);
		when "0110000001100000" => data_out <= rom_array(24672);
		when "0110000001100001" => data_out <= rom_array(24673);
		when "0110000001100010" => data_out <= rom_array(24674);
		when "0110000001100011" => data_out <= rom_array(24675);
		when "0110000001100100" => data_out <= rom_array(24676);
		when "0110000001100101" => data_out <= rom_array(24677);
		when "0110000001100110" => data_out <= rom_array(24678);
		when "0110000001100111" => data_out <= rom_array(24679);
		when "0110000001101000" => data_out <= rom_array(24680);
		when "0110000001101001" => data_out <= rom_array(24681);
		when "0110000001101010" => data_out <= rom_array(24682);
		when "0110000001101011" => data_out <= rom_array(24683);
		when "0110000001101100" => data_out <= rom_array(24684);
		when "0110000001101101" => data_out <= rom_array(24685);
		when "0110000001101110" => data_out <= rom_array(24686);
		when "0110000001101111" => data_out <= rom_array(24687);
		when "0110000001110000" => data_out <= rom_array(24688);
		when "0110000001110001" => data_out <= rom_array(24689);
		when "0110000001110010" => data_out <= rom_array(24690);
		when "0110000001110011" => data_out <= rom_array(24691);
		when "0110000001110100" => data_out <= rom_array(24692);
		when "0110000001110101" => data_out <= rom_array(24693);
		when "0110000001110110" => data_out <= rom_array(24694);
		when "0110000001110111" => data_out <= rom_array(24695);
		when "0110000001111000" => data_out <= rom_array(24696);
		when "0110000001111001" => data_out <= rom_array(24697);
		when "0110000001111010" => data_out <= rom_array(24698);
		when "0110000001111011" => data_out <= rom_array(24699);
		when "0110000001111100" => data_out <= rom_array(24700);
		when "0110000001111101" => data_out <= rom_array(24701);
		when "0110000001111110" => data_out <= rom_array(24702);
		when "0110000001111111" => data_out <= rom_array(24703);
		when "0110000010000000" => data_out <= rom_array(24704);
		when "0110000010000001" => data_out <= rom_array(24705);
		when "0110000010000010" => data_out <= rom_array(24706);
		when "0110000010000011" => data_out <= rom_array(24707);
		when "0110000010000100" => data_out <= rom_array(24708);
		when "0110000010000101" => data_out <= rom_array(24709);
		when "0110000010000110" => data_out <= rom_array(24710);
		when "0110000010000111" => data_out <= rom_array(24711);
		when "0110000010001000" => data_out <= rom_array(24712);
		when "0110000010001001" => data_out <= rom_array(24713);
		when "0110000010001010" => data_out <= rom_array(24714);
		when "0110000010001011" => data_out <= rom_array(24715);
		when "0110000010001100" => data_out <= rom_array(24716);
		when "0110000010001101" => data_out <= rom_array(24717);
		when "0110000010001110" => data_out <= rom_array(24718);
		when "0110000010001111" => data_out <= rom_array(24719);
		when "0110000010010000" => data_out <= rom_array(24720);
		when "0110000010010001" => data_out <= rom_array(24721);
		when "0110000010010010" => data_out <= rom_array(24722);
		when "0110000010010011" => data_out <= rom_array(24723);
		when "0110000010010100" => data_out <= rom_array(24724);
		when "0110000010010101" => data_out <= rom_array(24725);
		when "0110000010010110" => data_out <= rom_array(24726);
		when "0110000010010111" => data_out <= rom_array(24727);
		when "0110000010011000" => data_out <= rom_array(24728);
		when "0110000010011001" => data_out <= rom_array(24729);
		when "0110000010011010" => data_out <= rom_array(24730);
		when "0110000010011011" => data_out <= rom_array(24731);
		when "0110000010011100" => data_out <= rom_array(24732);
		when "0110000010011101" => data_out <= rom_array(24733);
		when "0110000010011110" => data_out <= rom_array(24734);
		when "0110000010011111" => data_out <= rom_array(24735);
		when "0110000010100000" => data_out <= rom_array(24736);
		when "0110000010100001" => data_out <= rom_array(24737);
		when "0110000010100010" => data_out <= rom_array(24738);
		when "0110000010100011" => data_out <= rom_array(24739);
		when "0110000010100100" => data_out <= rom_array(24740);
		when "0110000010100101" => data_out <= rom_array(24741);
		when "0110000010100110" => data_out <= rom_array(24742);
		when "0110000010100111" => data_out <= rom_array(24743);
		when "0110000010101000" => data_out <= rom_array(24744);
		when "0110000010101001" => data_out <= rom_array(24745);
		when "0110000010101010" => data_out <= rom_array(24746);
		when "0110000010101011" => data_out <= rom_array(24747);
		when "0110000010101100" => data_out <= rom_array(24748);
		when "0110000010101101" => data_out <= rom_array(24749);
		when "0110000010101110" => data_out <= rom_array(24750);
		when "0110000010101111" => data_out <= rom_array(24751);
		when "0110000010110000" => data_out <= rom_array(24752);
		when "0110000010110001" => data_out <= rom_array(24753);
		when "0110000010110010" => data_out <= rom_array(24754);
		when "0110000010110011" => data_out <= rom_array(24755);
		when "0110000010110100" => data_out <= rom_array(24756);
		when "0110000010110101" => data_out <= rom_array(24757);
		when "0110000010110110" => data_out <= rom_array(24758);
		when "0110000010110111" => data_out <= rom_array(24759);
		when "0110000010111000" => data_out <= rom_array(24760);
		when "0110000010111001" => data_out <= rom_array(24761);
		when "0110000010111010" => data_out <= rom_array(24762);
		when "0110000010111011" => data_out <= rom_array(24763);
		when "0110000010111100" => data_out <= rom_array(24764);
		when "0110000010111101" => data_out <= rom_array(24765);
		when "0110000010111110" => data_out <= rom_array(24766);
		when "0110000010111111" => data_out <= rom_array(24767);
		when "0110000011000000" => data_out <= rom_array(24768);
		when "0110000011000001" => data_out <= rom_array(24769);
		when "0110000011000010" => data_out <= rom_array(24770);
		when "0110000011000011" => data_out <= rom_array(24771);
		when "0110000011000100" => data_out <= rom_array(24772);
		when "0110000011000101" => data_out <= rom_array(24773);
		when "0110000011000110" => data_out <= rom_array(24774);
		when "0110000011000111" => data_out <= rom_array(24775);
		when "0110000011001000" => data_out <= rom_array(24776);
		when "0110000011001001" => data_out <= rom_array(24777);
		when "0110000011001010" => data_out <= rom_array(24778);
		when "0110000011001011" => data_out <= rom_array(24779);
		when "0110000011001100" => data_out <= rom_array(24780);
		when "0110000011001101" => data_out <= rom_array(24781);
		when "0110000011001110" => data_out <= rom_array(24782);
		when "0110000011001111" => data_out <= rom_array(24783);
		when "0110000011010000" => data_out <= rom_array(24784);
		when "0110000011010001" => data_out <= rom_array(24785);
		when "0110000011010010" => data_out <= rom_array(24786);
		when "0110000011010011" => data_out <= rom_array(24787);
		when "0110000011010100" => data_out <= rom_array(24788);
		when "0110000011010101" => data_out <= rom_array(24789);
		when "0110000011010110" => data_out <= rom_array(24790);
		when "0110000011010111" => data_out <= rom_array(24791);
		when "0110000011011000" => data_out <= rom_array(24792);
		when "0110000011011001" => data_out <= rom_array(24793);
		when "0110000011011010" => data_out <= rom_array(24794);
		when "0110000011011011" => data_out <= rom_array(24795);
		when "0110000011011100" => data_out <= rom_array(24796);
		when "0110000011011101" => data_out <= rom_array(24797);
		when "0110000011011110" => data_out <= rom_array(24798);
		when "0110000011011111" => data_out <= rom_array(24799);
		when "0110000011100000" => data_out <= rom_array(24800);
		when "0110000011100001" => data_out <= rom_array(24801);
		when "0110000011100010" => data_out <= rom_array(24802);
		when "0110000011100011" => data_out <= rom_array(24803);
		when "0110000011100100" => data_out <= rom_array(24804);
		when "0110000011100101" => data_out <= rom_array(24805);
		when "0110000011100110" => data_out <= rom_array(24806);
		when "0110000011100111" => data_out <= rom_array(24807);
		when "0110000011101000" => data_out <= rom_array(24808);
		when "0110000011101001" => data_out <= rom_array(24809);
		when "0110000011101010" => data_out <= rom_array(24810);
		when "0110000011101011" => data_out <= rom_array(24811);
		when "0110000011101100" => data_out <= rom_array(24812);
		when "0110000011101101" => data_out <= rom_array(24813);
		when "0110000011101110" => data_out <= rom_array(24814);
		when "0110000011101111" => data_out <= rom_array(24815);
		when "0110000011110000" => data_out <= rom_array(24816);
		when "0110000011110001" => data_out <= rom_array(24817);
		when "0110000011110010" => data_out <= rom_array(24818);
		when "0110000011110011" => data_out <= rom_array(24819);
		when "0110000011110100" => data_out <= rom_array(24820);
		when "0110000011110101" => data_out <= rom_array(24821);
		when "0110000011110110" => data_out <= rom_array(24822);
		when "0110000011110111" => data_out <= rom_array(24823);
		when "0110000011111000" => data_out <= rom_array(24824);
		when "0110000011111001" => data_out <= rom_array(24825);
		when "0110000011111010" => data_out <= rom_array(24826);
		when "0110000011111011" => data_out <= rom_array(24827);
		when "0110000011111100" => data_out <= rom_array(24828);
		when "0110000011111101" => data_out <= rom_array(24829);
		when "0110000011111110" => data_out <= rom_array(24830);
		when "0110000011111111" => data_out <= rom_array(24831);
		when "0110000100000000" => data_out <= rom_array(24832);
		when "0110000100000001" => data_out <= rom_array(24833);
		when "0110000100000010" => data_out <= rom_array(24834);
		when "0110000100000011" => data_out <= rom_array(24835);
		when "0110000100000100" => data_out <= rom_array(24836);
		when "0110000100000101" => data_out <= rom_array(24837);
		when "0110000100000110" => data_out <= rom_array(24838);
		when "0110000100000111" => data_out <= rom_array(24839);
		when "0110000100001000" => data_out <= rom_array(24840);
		when "0110000100001001" => data_out <= rom_array(24841);
		when "0110000100001010" => data_out <= rom_array(24842);
		when "0110000100001011" => data_out <= rom_array(24843);
		when "0110000100001100" => data_out <= rom_array(24844);
		when "0110000100001101" => data_out <= rom_array(24845);
		when "0110000100001110" => data_out <= rom_array(24846);
		when "0110000100001111" => data_out <= rom_array(24847);
		when "0110000100010000" => data_out <= rom_array(24848);
		when "0110000100010001" => data_out <= rom_array(24849);
		when "0110000100010010" => data_out <= rom_array(24850);
		when "0110000100010011" => data_out <= rom_array(24851);
		when "0110000100010100" => data_out <= rom_array(24852);
		when "0110000100010101" => data_out <= rom_array(24853);
		when "0110000100010110" => data_out <= rom_array(24854);
		when "0110000100010111" => data_out <= rom_array(24855);
		when "0110000100011000" => data_out <= rom_array(24856);
		when "0110000100011001" => data_out <= rom_array(24857);
		when "0110000100011010" => data_out <= rom_array(24858);
		when "0110000100011011" => data_out <= rom_array(24859);
		when "0110000100011100" => data_out <= rom_array(24860);
		when "0110000100011101" => data_out <= rom_array(24861);
		when "0110000100011110" => data_out <= rom_array(24862);
		when "0110000100011111" => data_out <= rom_array(24863);
		when "0110000100100000" => data_out <= rom_array(24864);
		when "0110000100100001" => data_out <= rom_array(24865);
		when "0110000100100010" => data_out <= rom_array(24866);
		when "0110000100100011" => data_out <= rom_array(24867);
		when "0110000100100100" => data_out <= rom_array(24868);
		when "0110000100100101" => data_out <= rom_array(24869);
		when "0110000100100110" => data_out <= rom_array(24870);
		when "0110000100100111" => data_out <= rom_array(24871);
		when "0110000100101000" => data_out <= rom_array(24872);
		when "0110000100101001" => data_out <= rom_array(24873);
		when "0110000100101010" => data_out <= rom_array(24874);
		when "0110000100101011" => data_out <= rom_array(24875);
		when "0110000100101100" => data_out <= rom_array(24876);
		when "0110000100101101" => data_out <= rom_array(24877);
		when "0110000100101110" => data_out <= rom_array(24878);
		when "0110000100101111" => data_out <= rom_array(24879);
		when "0110000100110000" => data_out <= rom_array(24880);
		when "0110000100110001" => data_out <= rom_array(24881);
		when "0110000100110010" => data_out <= rom_array(24882);
		when "0110000100110011" => data_out <= rom_array(24883);
		when "0110000100110100" => data_out <= rom_array(24884);
		when "0110000100110101" => data_out <= rom_array(24885);
		when "0110000100110110" => data_out <= rom_array(24886);
		when "0110000100110111" => data_out <= rom_array(24887);
		when "0110000100111000" => data_out <= rom_array(24888);
		when "0110000100111001" => data_out <= rom_array(24889);
		when "0110000100111010" => data_out <= rom_array(24890);
		when "0110000100111011" => data_out <= rom_array(24891);
		when "0110000100111100" => data_out <= rom_array(24892);
		when "0110000100111101" => data_out <= rom_array(24893);
		when "0110000100111110" => data_out <= rom_array(24894);
		when "0110000100111111" => data_out <= rom_array(24895);
		when "0110000101000000" => data_out <= rom_array(24896);
		when "0110000101000001" => data_out <= rom_array(24897);
		when "0110000101000010" => data_out <= rom_array(24898);
		when "0110000101000011" => data_out <= rom_array(24899);
		when "0110000101000100" => data_out <= rom_array(24900);
		when "0110000101000101" => data_out <= rom_array(24901);
		when "0110000101000110" => data_out <= rom_array(24902);
		when "0110000101000111" => data_out <= rom_array(24903);
		when "0110000101001000" => data_out <= rom_array(24904);
		when "0110000101001001" => data_out <= rom_array(24905);
		when "0110000101001010" => data_out <= rom_array(24906);
		when "0110000101001011" => data_out <= rom_array(24907);
		when "0110000101001100" => data_out <= rom_array(24908);
		when "0110000101001101" => data_out <= rom_array(24909);
		when "0110000101001110" => data_out <= rom_array(24910);
		when "0110000101001111" => data_out <= rom_array(24911);
		when "0110000101010000" => data_out <= rom_array(24912);
		when "0110000101010001" => data_out <= rom_array(24913);
		when "0110000101010010" => data_out <= rom_array(24914);
		when "0110000101010011" => data_out <= rom_array(24915);
		when "0110000101010100" => data_out <= rom_array(24916);
		when "0110000101010101" => data_out <= rom_array(24917);
		when "0110000101010110" => data_out <= rom_array(24918);
		when "0110000101010111" => data_out <= rom_array(24919);
		when "0110000101011000" => data_out <= rom_array(24920);
		when "0110000101011001" => data_out <= rom_array(24921);
		when "0110000101011010" => data_out <= rom_array(24922);
		when "0110000101011011" => data_out <= rom_array(24923);
		when "0110000101011100" => data_out <= rom_array(24924);
		when "0110000101011101" => data_out <= rom_array(24925);
		when "0110000101011110" => data_out <= rom_array(24926);
		when "0110000101011111" => data_out <= rom_array(24927);
		when "0110000101100000" => data_out <= rom_array(24928);
		when "0110000101100001" => data_out <= rom_array(24929);
		when "0110000101100010" => data_out <= rom_array(24930);
		when "0110000101100011" => data_out <= rom_array(24931);
		when "0110000101100100" => data_out <= rom_array(24932);
		when "0110000101100101" => data_out <= rom_array(24933);
		when "0110000101100110" => data_out <= rom_array(24934);
		when "0110000101100111" => data_out <= rom_array(24935);
		when "0110000101101000" => data_out <= rom_array(24936);
		when "0110000101101001" => data_out <= rom_array(24937);
		when "0110000101101010" => data_out <= rom_array(24938);
		when "0110000101101011" => data_out <= rom_array(24939);
		when "0110000101101100" => data_out <= rom_array(24940);
		when "0110000101101101" => data_out <= rom_array(24941);
		when "0110000101101110" => data_out <= rom_array(24942);
		when "0110000101101111" => data_out <= rom_array(24943);
		when "0110000101110000" => data_out <= rom_array(24944);
		when "0110000101110001" => data_out <= rom_array(24945);
		when "0110000101110010" => data_out <= rom_array(24946);
		when "0110000101110011" => data_out <= rom_array(24947);
		when "0110000101110100" => data_out <= rom_array(24948);
		when "0110000101110101" => data_out <= rom_array(24949);
		when "0110000101110110" => data_out <= rom_array(24950);
		when "0110000101110111" => data_out <= rom_array(24951);
		when "0110000101111000" => data_out <= rom_array(24952);
		when "0110000101111001" => data_out <= rom_array(24953);
		when "0110000101111010" => data_out <= rom_array(24954);
		when "0110000101111011" => data_out <= rom_array(24955);
		when "0110000101111100" => data_out <= rom_array(24956);
		when "0110000101111101" => data_out <= rom_array(24957);
		when "0110000101111110" => data_out <= rom_array(24958);
		when "0110000101111111" => data_out <= rom_array(24959);
		when "0110000110000000" => data_out <= rom_array(24960);
		when "0110000110000001" => data_out <= rom_array(24961);
		when "0110000110000010" => data_out <= rom_array(24962);
		when "0110000110000011" => data_out <= rom_array(24963);
		when "0110000110000100" => data_out <= rom_array(24964);
		when "0110000110000101" => data_out <= rom_array(24965);
		when "0110000110000110" => data_out <= rom_array(24966);
		when "0110000110000111" => data_out <= rom_array(24967);
		when "0110000110001000" => data_out <= rom_array(24968);
		when "0110000110001001" => data_out <= rom_array(24969);
		when "0110000110001010" => data_out <= rom_array(24970);
		when "0110000110001011" => data_out <= rom_array(24971);
		when "0110000110001100" => data_out <= rom_array(24972);
		when "0110000110001101" => data_out <= rom_array(24973);
		when "0110000110001110" => data_out <= rom_array(24974);
		when "0110000110001111" => data_out <= rom_array(24975);
		when "0110000110010000" => data_out <= rom_array(24976);
		when "0110000110010001" => data_out <= rom_array(24977);
		when "0110000110010010" => data_out <= rom_array(24978);
		when "0110000110010011" => data_out <= rom_array(24979);
		when "0110000110010100" => data_out <= rom_array(24980);
		when "0110000110010101" => data_out <= rom_array(24981);
		when "0110000110010110" => data_out <= rom_array(24982);
		when "0110000110010111" => data_out <= rom_array(24983);
		when "0110000110011000" => data_out <= rom_array(24984);
		when "0110000110011001" => data_out <= rom_array(24985);
		when "0110000110011010" => data_out <= rom_array(24986);
		when "0110000110011011" => data_out <= rom_array(24987);
		when "0110000110011100" => data_out <= rom_array(24988);
		when "0110000110011101" => data_out <= rom_array(24989);
		when "0110000110011110" => data_out <= rom_array(24990);
		when "0110000110011111" => data_out <= rom_array(24991);
		when "0110000110100000" => data_out <= rom_array(24992);
		when "0110000110100001" => data_out <= rom_array(24993);
		when "0110000110100010" => data_out <= rom_array(24994);
		when "0110000110100011" => data_out <= rom_array(24995);
		when "0110000110100100" => data_out <= rom_array(24996);
		when "0110000110100101" => data_out <= rom_array(24997);
		when "0110000110100110" => data_out <= rom_array(24998);
		when "0110000110100111" => data_out <= rom_array(24999);
		when "0110000110101000" => data_out <= rom_array(25000);
		when "0110000110101001" => data_out <= rom_array(25001);
		when "0110000110101010" => data_out <= rom_array(25002);
		when "0110000110101011" => data_out <= rom_array(25003);
		when "0110000110101100" => data_out <= rom_array(25004);
		when "0110000110101101" => data_out <= rom_array(25005);
		when "0110000110101110" => data_out <= rom_array(25006);
		when "0110000110101111" => data_out <= rom_array(25007);
		when "0110000110110000" => data_out <= rom_array(25008);
		when "0110000110110001" => data_out <= rom_array(25009);
		when "0110000110110010" => data_out <= rom_array(25010);
		when "0110000110110011" => data_out <= rom_array(25011);
		when "0110000110110100" => data_out <= rom_array(25012);
		when "0110000110110101" => data_out <= rom_array(25013);
		when "0110000110110110" => data_out <= rom_array(25014);
		when "0110000110110111" => data_out <= rom_array(25015);
		when "0110000110111000" => data_out <= rom_array(25016);
		when "0110000110111001" => data_out <= rom_array(25017);
		when "0110000110111010" => data_out <= rom_array(25018);
		when "0110000110111011" => data_out <= rom_array(25019);
		when "0110000110111100" => data_out <= rom_array(25020);
		when "0110000110111101" => data_out <= rom_array(25021);
		when "0110000110111110" => data_out <= rom_array(25022);
		when "0110000110111111" => data_out <= rom_array(25023);
		when "0110000111000000" => data_out <= rom_array(25024);
		when "0110000111000001" => data_out <= rom_array(25025);
		when "0110000111000010" => data_out <= rom_array(25026);
		when "0110000111000011" => data_out <= rom_array(25027);
		when "0110000111000100" => data_out <= rom_array(25028);
		when "0110000111000101" => data_out <= rom_array(25029);
		when "0110000111000110" => data_out <= rom_array(25030);
		when "0110000111000111" => data_out <= rom_array(25031);
		when "0110000111001000" => data_out <= rom_array(25032);
		when "0110000111001001" => data_out <= rom_array(25033);
		when "0110000111001010" => data_out <= rom_array(25034);
		when "0110000111001011" => data_out <= rom_array(25035);
		when "0110000111001100" => data_out <= rom_array(25036);
		when "0110000111001101" => data_out <= rom_array(25037);
		when "0110000111001110" => data_out <= rom_array(25038);
		when "0110000111001111" => data_out <= rom_array(25039);
		when "0110000111010000" => data_out <= rom_array(25040);
		when "0110000111010001" => data_out <= rom_array(25041);
		when "0110000111010010" => data_out <= rom_array(25042);
		when "0110000111010011" => data_out <= rom_array(25043);
		when "0110000111010100" => data_out <= rom_array(25044);
		when "0110000111010101" => data_out <= rom_array(25045);
		when "0110000111010110" => data_out <= rom_array(25046);
		when "0110000111010111" => data_out <= rom_array(25047);
		when "0110000111011000" => data_out <= rom_array(25048);
		when "0110000111011001" => data_out <= rom_array(25049);
		when "0110000111011010" => data_out <= rom_array(25050);
		when "0110000111011011" => data_out <= rom_array(25051);
		when "0110000111011100" => data_out <= rom_array(25052);
		when "0110000111011101" => data_out <= rom_array(25053);
		when "0110000111011110" => data_out <= rom_array(25054);
		when "0110000111011111" => data_out <= rom_array(25055);
		when "0110000111100000" => data_out <= rom_array(25056);
		when "0110000111100001" => data_out <= rom_array(25057);
		when "0110000111100010" => data_out <= rom_array(25058);
		when "0110000111100011" => data_out <= rom_array(25059);
		when "0110000111100100" => data_out <= rom_array(25060);
		when "0110000111100101" => data_out <= rom_array(25061);
		when "0110000111100110" => data_out <= rom_array(25062);
		when "0110000111100111" => data_out <= rom_array(25063);
		when "0110000111101000" => data_out <= rom_array(25064);
		when "0110000111101001" => data_out <= rom_array(25065);
		when "0110000111101010" => data_out <= rom_array(25066);
		when "0110000111101011" => data_out <= rom_array(25067);
		when "0110000111101100" => data_out <= rom_array(25068);
		when "0110000111101101" => data_out <= rom_array(25069);
		when "0110000111101110" => data_out <= rom_array(25070);
		when "0110000111101111" => data_out <= rom_array(25071);
		when "0110000111110000" => data_out <= rom_array(25072);
		when "0110000111110001" => data_out <= rom_array(25073);
		when "0110000111110010" => data_out <= rom_array(25074);
		when "0110000111110011" => data_out <= rom_array(25075);
		when "0110000111110100" => data_out <= rom_array(25076);
		when "0110000111110101" => data_out <= rom_array(25077);
		when "0110000111110110" => data_out <= rom_array(25078);
		when "0110000111110111" => data_out <= rom_array(25079);
		when "0110000111111000" => data_out <= rom_array(25080);
		when "0110000111111001" => data_out <= rom_array(25081);
		when "0110000111111010" => data_out <= rom_array(25082);
		when "0110000111111011" => data_out <= rom_array(25083);
		when "0110000111111100" => data_out <= rom_array(25084);
		when "0110000111111101" => data_out <= rom_array(25085);
		when "0110000111111110" => data_out <= rom_array(25086);
		when "0110000111111111" => data_out <= rom_array(25087);
		when "0110001000000000" => data_out <= rom_array(25088);
		when "0110001000000001" => data_out <= rom_array(25089);
		when "0110001000000010" => data_out <= rom_array(25090);
		when "0110001000000011" => data_out <= rom_array(25091);
		when "0110001000000100" => data_out <= rom_array(25092);
		when "0110001000000101" => data_out <= rom_array(25093);
		when "0110001000000110" => data_out <= rom_array(25094);
		when "0110001000000111" => data_out <= rom_array(25095);
		when "0110001000001000" => data_out <= rom_array(25096);
		when "0110001000001001" => data_out <= rom_array(25097);
		when "0110001000001010" => data_out <= rom_array(25098);
		when "0110001000001011" => data_out <= rom_array(25099);
		when "0110001000001100" => data_out <= rom_array(25100);
		when "0110001000001101" => data_out <= rom_array(25101);
		when "0110001000001110" => data_out <= rom_array(25102);
		when "0110001000001111" => data_out <= rom_array(25103);
		when "0110001000010000" => data_out <= rom_array(25104);
		when "0110001000010001" => data_out <= rom_array(25105);
		when "0110001000010010" => data_out <= rom_array(25106);
		when "0110001000010011" => data_out <= rom_array(25107);
		when "0110001000010100" => data_out <= rom_array(25108);
		when "0110001000010101" => data_out <= rom_array(25109);
		when "0110001000010110" => data_out <= rom_array(25110);
		when "0110001000010111" => data_out <= rom_array(25111);
		when "0110001000011000" => data_out <= rom_array(25112);
		when "0110001000011001" => data_out <= rom_array(25113);
		when "0110001000011010" => data_out <= rom_array(25114);
		when "0110001000011011" => data_out <= rom_array(25115);
		when "0110001000011100" => data_out <= rom_array(25116);
		when "0110001000011101" => data_out <= rom_array(25117);
		when "0110001000011110" => data_out <= rom_array(25118);
		when "0110001000011111" => data_out <= rom_array(25119);
		when "0110001000100000" => data_out <= rom_array(25120);
		when "0110001000100001" => data_out <= rom_array(25121);
		when "0110001000100010" => data_out <= rom_array(25122);
		when "0110001000100011" => data_out <= rom_array(25123);
		when "0110001000100100" => data_out <= rom_array(25124);
		when "0110001000100101" => data_out <= rom_array(25125);
		when "0110001000100110" => data_out <= rom_array(25126);
		when "0110001000100111" => data_out <= rom_array(25127);
		when "0110001000101000" => data_out <= rom_array(25128);
		when "0110001000101001" => data_out <= rom_array(25129);
		when "0110001000101010" => data_out <= rom_array(25130);
		when "0110001000101011" => data_out <= rom_array(25131);
		when "0110001000101100" => data_out <= rom_array(25132);
		when "0110001000101101" => data_out <= rom_array(25133);
		when "0110001000101110" => data_out <= rom_array(25134);
		when "0110001000101111" => data_out <= rom_array(25135);
		when "0110001000110000" => data_out <= rom_array(25136);
		when "0110001000110001" => data_out <= rom_array(25137);
		when "0110001000110010" => data_out <= rom_array(25138);
		when "0110001000110011" => data_out <= rom_array(25139);
		when "0110001000110100" => data_out <= rom_array(25140);
		when "0110001000110101" => data_out <= rom_array(25141);
		when "0110001000110110" => data_out <= rom_array(25142);
		when "0110001000110111" => data_out <= rom_array(25143);
		when "0110001000111000" => data_out <= rom_array(25144);
		when "0110001000111001" => data_out <= rom_array(25145);
		when "0110001000111010" => data_out <= rom_array(25146);
		when "0110001000111011" => data_out <= rom_array(25147);
		when "0110001000111100" => data_out <= rom_array(25148);
		when "0110001000111101" => data_out <= rom_array(25149);
		when "0110001000111110" => data_out <= rom_array(25150);
		when "0110001000111111" => data_out <= rom_array(25151);
		when "0110001001000000" => data_out <= rom_array(25152);
		when "0110001001000001" => data_out <= rom_array(25153);
		when "0110001001000010" => data_out <= rom_array(25154);
		when "0110001001000011" => data_out <= rom_array(25155);
		when "0110001001000100" => data_out <= rom_array(25156);
		when "0110001001000101" => data_out <= rom_array(25157);
		when "0110001001000110" => data_out <= rom_array(25158);
		when "0110001001000111" => data_out <= rom_array(25159);
		when "0110001001001000" => data_out <= rom_array(25160);
		when "0110001001001001" => data_out <= rom_array(25161);
		when "0110001001001010" => data_out <= rom_array(25162);
		when "0110001001001011" => data_out <= rom_array(25163);
		when "0110001001001100" => data_out <= rom_array(25164);
		when "0110001001001101" => data_out <= rom_array(25165);
		when "0110001001001110" => data_out <= rom_array(25166);
		when "0110001001001111" => data_out <= rom_array(25167);
		when "0110001001010000" => data_out <= rom_array(25168);
		when "0110001001010001" => data_out <= rom_array(25169);
		when "0110001001010010" => data_out <= rom_array(25170);
		when "0110001001010011" => data_out <= rom_array(25171);
		when "0110001001010100" => data_out <= rom_array(25172);
		when "0110001001010101" => data_out <= rom_array(25173);
		when "0110001001010110" => data_out <= rom_array(25174);
		when "0110001001010111" => data_out <= rom_array(25175);
		when "0110001001011000" => data_out <= rom_array(25176);
		when "0110001001011001" => data_out <= rom_array(25177);
		when "0110001001011010" => data_out <= rom_array(25178);
		when "0110001001011011" => data_out <= rom_array(25179);
		when "0110001001011100" => data_out <= rom_array(25180);
		when "0110001001011101" => data_out <= rom_array(25181);
		when "0110001001011110" => data_out <= rom_array(25182);
		when "0110001001011111" => data_out <= rom_array(25183);
		when "0110001001100000" => data_out <= rom_array(25184);
		when "0110001001100001" => data_out <= rom_array(25185);
		when "0110001001100010" => data_out <= rom_array(25186);
		when "0110001001100011" => data_out <= rom_array(25187);
		when "0110001001100100" => data_out <= rom_array(25188);
		when "0110001001100101" => data_out <= rom_array(25189);
		when "0110001001100110" => data_out <= rom_array(25190);
		when "0110001001100111" => data_out <= rom_array(25191);
		when "0110001001101000" => data_out <= rom_array(25192);
		when "0110001001101001" => data_out <= rom_array(25193);
		when "0110001001101010" => data_out <= rom_array(25194);
		when "0110001001101011" => data_out <= rom_array(25195);
		when "0110001001101100" => data_out <= rom_array(25196);
		when "0110001001101101" => data_out <= rom_array(25197);
		when "0110001001101110" => data_out <= rom_array(25198);
		when "0110001001101111" => data_out <= rom_array(25199);
		when "0110001001110000" => data_out <= rom_array(25200);
		when "0110001001110001" => data_out <= rom_array(25201);
		when "0110001001110010" => data_out <= rom_array(25202);
		when "0110001001110011" => data_out <= rom_array(25203);
		when "0110001001110100" => data_out <= rom_array(25204);
		when "0110001001110101" => data_out <= rom_array(25205);
		when "0110001001110110" => data_out <= rom_array(25206);
		when "0110001001110111" => data_out <= rom_array(25207);
		when "0110001001111000" => data_out <= rom_array(25208);
		when "0110001001111001" => data_out <= rom_array(25209);
		when "0110001001111010" => data_out <= rom_array(25210);
		when "0110001001111011" => data_out <= rom_array(25211);
		when "0110001001111100" => data_out <= rom_array(25212);
		when "0110001001111101" => data_out <= rom_array(25213);
		when "0110001001111110" => data_out <= rom_array(25214);
		when "0110001001111111" => data_out <= rom_array(25215);
		when "0110001010000000" => data_out <= rom_array(25216);
		when "0110001010000001" => data_out <= rom_array(25217);
		when "0110001010000010" => data_out <= rom_array(25218);
		when "0110001010000011" => data_out <= rom_array(25219);
		when "0110001010000100" => data_out <= rom_array(25220);
		when "0110001010000101" => data_out <= rom_array(25221);
		when "0110001010000110" => data_out <= rom_array(25222);
		when "0110001010000111" => data_out <= rom_array(25223);
		when "0110001010001000" => data_out <= rom_array(25224);
		when "0110001010001001" => data_out <= rom_array(25225);
		when "0110001010001010" => data_out <= rom_array(25226);
		when "0110001010001011" => data_out <= rom_array(25227);
		when "0110001010001100" => data_out <= rom_array(25228);
		when "0110001010001101" => data_out <= rom_array(25229);
		when "0110001010001110" => data_out <= rom_array(25230);
		when "0110001010001111" => data_out <= rom_array(25231);
		when "0110001010010000" => data_out <= rom_array(25232);
		when "0110001010010001" => data_out <= rom_array(25233);
		when "0110001010010010" => data_out <= rom_array(25234);
		when "0110001010010011" => data_out <= rom_array(25235);
		when "0110001010010100" => data_out <= rom_array(25236);
		when "0110001010010101" => data_out <= rom_array(25237);
		when "0110001010010110" => data_out <= rom_array(25238);
		when "0110001010010111" => data_out <= rom_array(25239);
		when "0110001010011000" => data_out <= rom_array(25240);
		when "0110001010011001" => data_out <= rom_array(25241);
		when "0110001010011010" => data_out <= rom_array(25242);
		when "0110001010011011" => data_out <= rom_array(25243);
		when "0110001010011100" => data_out <= rom_array(25244);
		when "0110001010011101" => data_out <= rom_array(25245);
		when "0110001010011110" => data_out <= rom_array(25246);
		when "0110001010011111" => data_out <= rom_array(25247);
		when "0110001010100000" => data_out <= rom_array(25248);
		when "0110001010100001" => data_out <= rom_array(25249);
		when "0110001010100010" => data_out <= rom_array(25250);
		when "0110001010100011" => data_out <= rom_array(25251);
		when "0110001010100100" => data_out <= rom_array(25252);
		when "0110001010100101" => data_out <= rom_array(25253);
		when "0110001010100110" => data_out <= rom_array(25254);
		when "0110001010100111" => data_out <= rom_array(25255);
		when "0110001010101000" => data_out <= rom_array(25256);
		when "0110001010101001" => data_out <= rom_array(25257);
		when "0110001010101010" => data_out <= rom_array(25258);
		when "0110001010101011" => data_out <= rom_array(25259);
		when "0110001010101100" => data_out <= rom_array(25260);
		when "0110001010101101" => data_out <= rom_array(25261);
		when "0110001010101110" => data_out <= rom_array(25262);
		when "0110001010101111" => data_out <= rom_array(25263);
		when "0110001010110000" => data_out <= rom_array(25264);
		when "0110001010110001" => data_out <= rom_array(25265);
		when "0110001010110010" => data_out <= rom_array(25266);
		when "0110001010110011" => data_out <= rom_array(25267);
		when "0110001010110100" => data_out <= rom_array(25268);
		when "0110001010110101" => data_out <= rom_array(25269);
		when "0110001010110110" => data_out <= rom_array(25270);
		when "0110001010110111" => data_out <= rom_array(25271);
		when "0110001010111000" => data_out <= rom_array(25272);
		when "0110001010111001" => data_out <= rom_array(25273);
		when "0110001010111010" => data_out <= rom_array(25274);
		when "0110001010111011" => data_out <= rom_array(25275);
		when "0110001010111100" => data_out <= rom_array(25276);
		when "0110001010111101" => data_out <= rom_array(25277);
		when "0110001010111110" => data_out <= rom_array(25278);
		when "0110001010111111" => data_out <= rom_array(25279);
		when "0110001011000000" => data_out <= rom_array(25280);
		when "0110001011000001" => data_out <= rom_array(25281);
		when "0110001011000010" => data_out <= rom_array(25282);
		when "0110001011000011" => data_out <= rom_array(25283);
		when "0110001011000100" => data_out <= rom_array(25284);
		when "0110001011000101" => data_out <= rom_array(25285);
		when "0110001011000110" => data_out <= rom_array(25286);
		when "0110001011000111" => data_out <= rom_array(25287);
		when "0110001011001000" => data_out <= rom_array(25288);
		when "0110001011001001" => data_out <= rom_array(25289);
		when "0110001011001010" => data_out <= rom_array(25290);
		when "0110001011001011" => data_out <= rom_array(25291);
		when "0110001011001100" => data_out <= rom_array(25292);
		when "0110001011001101" => data_out <= rom_array(25293);
		when "0110001011001110" => data_out <= rom_array(25294);
		when "0110001011001111" => data_out <= rom_array(25295);
		when "0110001011010000" => data_out <= rom_array(25296);
		when "0110001011010001" => data_out <= rom_array(25297);
		when "0110001011010010" => data_out <= rom_array(25298);
		when "0110001011010011" => data_out <= rom_array(25299);
		when "0110001011010100" => data_out <= rom_array(25300);
		when "0110001011010101" => data_out <= rom_array(25301);
		when "0110001011010110" => data_out <= rom_array(25302);
		when "0110001011010111" => data_out <= rom_array(25303);
		when "0110001011011000" => data_out <= rom_array(25304);
		when "0110001011011001" => data_out <= rom_array(25305);
		when "0110001011011010" => data_out <= rom_array(25306);
		when "0110001011011011" => data_out <= rom_array(25307);
		when "0110001011011100" => data_out <= rom_array(25308);
		when "0110001011011101" => data_out <= rom_array(25309);
		when "0110001011011110" => data_out <= rom_array(25310);
		when "0110001011011111" => data_out <= rom_array(25311);
		when "0110001011100000" => data_out <= rom_array(25312);
		when "0110001011100001" => data_out <= rom_array(25313);
		when "0110001011100010" => data_out <= rom_array(25314);
		when "0110001011100011" => data_out <= rom_array(25315);
		when "0110001011100100" => data_out <= rom_array(25316);
		when "0110001011100101" => data_out <= rom_array(25317);
		when "0110001011100110" => data_out <= rom_array(25318);
		when "0110001011100111" => data_out <= rom_array(25319);
		when "0110001011101000" => data_out <= rom_array(25320);
		when "0110001011101001" => data_out <= rom_array(25321);
		when "0110001011101010" => data_out <= rom_array(25322);
		when "0110001011101011" => data_out <= rom_array(25323);
		when "0110001011101100" => data_out <= rom_array(25324);
		when "0110001011101101" => data_out <= rom_array(25325);
		when "0110001011101110" => data_out <= rom_array(25326);
		when "0110001011101111" => data_out <= rom_array(25327);
		when "0110001011110000" => data_out <= rom_array(25328);
		when "0110001011110001" => data_out <= rom_array(25329);
		when "0110001011110010" => data_out <= rom_array(25330);
		when "0110001011110011" => data_out <= rom_array(25331);
		when "0110001011110100" => data_out <= rom_array(25332);
		when "0110001011110101" => data_out <= rom_array(25333);
		when "0110001011110110" => data_out <= rom_array(25334);
		when "0110001011110111" => data_out <= rom_array(25335);
		when "0110001011111000" => data_out <= rom_array(25336);
		when "0110001011111001" => data_out <= rom_array(25337);
		when "0110001011111010" => data_out <= rom_array(25338);
		when "0110001011111011" => data_out <= rom_array(25339);
		when "0110001011111100" => data_out <= rom_array(25340);
		when "0110001011111101" => data_out <= rom_array(25341);
		when "0110001011111110" => data_out <= rom_array(25342);
		when "0110001011111111" => data_out <= rom_array(25343);
		when "0110001100000000" => data_out <= rom_array(25344);
		when "0110001100000001" => data_out <= rom_array(25345);
		when "0110001100000010" => data_out <= rom_array(25346);
		when "0110001100000011" => data_out <= rom_array(25347);
		when "0110001100000100" => data_out <= rom_array(25348);
		when "0110001100000101" => data_out <= rom_array(25349);
		when "0110001100000110" => data_out <= rom_array(25350);
		when "0110001100000111" => data_out <= rom_array(25351);
		when "0110001100001000" => data_out <= rom_array(25352);
		when "0110001100001001" => data_out <= rom_array(25353);
		when "0110001100001010" => data_out <= rom_array(25354);
		when "0110001100001011" => data_out <= rom_array(25355);
		when "0110001100001100" => data_out <= rom_array(25356);
		when "0110001100001101" => data_out <= rom_array(25357);
		when "0110001100001110" => data_out <= rom_array(25358);
		when "0110001100001111" => data_out <= rom_array(25359);
		when "0110001100010000" => data_out <= rom_array(25360);
		when "0110001100010001" => data_out <= rom_array(25361);
		when "0110001100010010" => data_out <= rom_array(25362);
		when "0110001100010011" => data_out <= rom_array(25363);
		when "0110001100010100" => data_out <= rom_array(25364);
		when "0110001100010101" => data_out <= rom_array(25365);
		when "0110001100010110" => data_out <= rom_array(25366);
		when "0110001100010111" => data_out <= rom_array(25367);
		when "0110001100011000" => data_out <= rom_array(25368);
		when "0110001100011001" => data_out <= rom_array(25369);
		when "0110001100011010" => data_out <= rom_array(25370);
		when "0110001100011011" => data_out <= rom_array(25371);
		when "0110001100011100" => data_out <= rom_array(25372);
		when "0110001100011101" => data_out <= rom_array(25373);
		when "0110001100011110" => data_out <= rom_array(25374);
		when "0110001100011111" => data_out <= rom_array(25375);
		when "0110001100100000" => data_out <= rom_array(25376);
		when "0110001100100001" => data_out <= rom_array(25377);
		when "0110001100100010" => data_out <= rom_array(25378);
		when "0110001100100011" => data_out <= rom_array(25379);
		when "0110001100100100" => data_out <= rom_array(25380);
		when "0110001100100101" => data_out <= rom_array(25381);
		when "0110001100100110" => data_out <= rom_array(25382);
		when "0110001100100111" => data_out <= rom_array(25383);
		when "0110001100101000" => data_out <= rom_array(25384);
		when "0110001100101001" => data_out <= rom_array(25385);
		when "0110001100101010" => data_out <= rom_array(25386);
		when "0110001100101011" => data_out <= rom_array(25387);
		when "0110001100101100" => data_out <= rom_array(25388);
		when "0110001100101101" => data_out <= rom_array(25389);
		when "0110001100101110" => data_out <= rom_array(25390);
		when "0110001100101111" => data_out <= rom_array(25391);
		when "0110001100110000" => data_out <= rom_array(25392);
		when "0110001100110001" => data_out <= rom_array(25393);
		when "0110001100110010" => data_out <= rom_array(25394);
		when "0110001100110011" => data_out <= rom_array(25395);
		when "0110001100110100" => data_out <= rom_array(25396);
		when "0110001100110101" => data_out <= rom_array(25397);
		when "0110001100110110" => data_out <= rom_array(25398);
		when "0110001100110111" => data_out <= rom_array(25399);
		when "0110001100111000" => data_out <= rom_array(25400);
		when "0110001100111001" => data_out <= rom_array(25401);
		when "0110001100111010" => data_out <= rom_array(25402);
		when "0110001100111011" => data_out <= rom_array(25403);
		when "0110001100111100" => data_out <= rom_array(25404);
		when "0110001100111101" => data_out <= rom_array(25405);
		when "0110001100111110" => data_out <= rom_array(25406);
		when "0110001100111111" => data_out <= rom_array(25407);
		when "0110001101000000" => data_out <= rom_array(25408);
		when "0110001101000001" => data_out <= rom_array(25409);
		when "0110001101000010" => data_out <= rom_array(25410);
		when "0110001101000011" => data_out <= rom_array(25411);
		when "0110001101000100" => data_out <= rom_array(25412);
		when "0110001101000101" => data_out <= rom_array(25413);
		when "0110001101000110" => data_out <= rom_array(25414);
		when "0110001101000111" => data_out <= rom_array(25415);
		when "0110001101001000" => data_out <= rom_array(25416);
		when "0110001101001001" => data_out <= rom_array(25417);
		when "0110001101001010" => data_out <= rom_array(25418);
		when "0110001101001011" => data_out <= rom_array(25419);
		when "0110001101001100" => data_out <= rom_array(25420);
		when "0110001101001101" => data_out <= rom_array(25421);
		when "0110001101001110" => data_out <= rom_array(25422);
		when "0110001101001111" => data_out <= rom_array(25423);
		when "0110001101010000" => data_out <= rom_array(25424);
		when "0110001101010001" => data_out <= rom_array(25425);
		when "0110001101010010" => data_out <= rom_array(25426);
		when "0110001101010011" => data_out <= rom_array(25427);
		when "0110001101010100" => data_out <= rom_array(25428);
		when "0110001101010101" => data_out <= rom_array(25429);
		when "0110001101010110" => data_out <= rom_array(25430);
		when "0110001101010111" => data_out <= rom_array(25431);
		when "0110001101011000" => data_out <= rom_array(25432);
		when "0110001101011001" => data_out <= rom_array(25433);
		when "0110001101011010" => data_out <= rom_array(25434);
		when "0110001101011011" => data_out <= rom_array(25435);
		when "0110001101011100" => data_out <= rom_array(25436);
		when "0110001101011101" => data_out <= rom_array(25437);
		when "0110001101011110" => data_out <= rom_array(25438);
		when "0110001101011111" => data_out <= rom_array(25439);
		when "0110001101100000" => data_out <= rom_array(25440);
		when "0110001101100001" => data_out <= rom_array(25441);
		when "0110001101100010" => data_out <= rom_array(25442);
		when "0110001101100011" => data_out <= rom_array(25443);
		when "0110001101100100" => data_out <= rom_array(25444);
		when "0110001101100101" => data_out <= rom_array(25445);
		when "0110001101100110" => data_out <= rom_array(25446);
		when "0110001101100111" => data_out <= rom_array(25447);
		when "0110001101101000" => data_out <= rom_array(25448);
		when "0110001101101001" => data_out <= rom_array(25449);
		when "0110001101101010" => data_out <= rom_array(25450);
		when "0110001101101011" => data_out <= rom_array(25451);
		when "0110001101101100" => data_out <= rom_array(25452);
		when "0110001101101101" => data_out <= rom_array(25453);
		when "0110001101101110" => data_out <= rom_array(25454);
		when "0110001101101111" => data_out <= rom_array(25455);
		when "0110001101110000" => data_out <= rom_array(25456);
		when "0110001101110001" => data_out <= rom_array(25457);
		when "0110001101110010" => data_out <= rom_array(25458);
		when "0110001101110011" => data_out <= rom_array(25459);
		when "0110001101110100" => data_out <= rom_array(25460);
		when "0110001101110101" => data_out <= rom_array(25461);
		when "0110001101110110" => data_out <= rom_array(25462);
		when "0110001101110111" => data_out <= rom_array(25463);
		when "0110001101111000" => data_out <= rom_array(25464);
		when "0110001101111001" => data_out <= rom_array(25465);
		when "0110001101111010" => data_out <= rom_array(25466);
		when "0110001101111011" => data_out <= rom_array(25467);
		when "0110001101111100" => data_out <= rom_array(25468);
		when "0110001101111101" => data_out <= rom_array(25469);
		when "0110001101111110" => data_out <= rom_array(25470);
		when "0110001101111111" => data_out <= rom_array(25471);
		when "0110001110000000" => data_out <= rom_array(25472);
		when "0110001110000001" => data_out <= rom_array(25473);
		when "0110001110000010" => data_out <= rom_array(25474);
		when "0110001110000011" => data_out <= rom_array(25475);
		when "0110001110000100" => data_out <= rom_array(25476);
		when "0110001110000101" => data_out <= rom_array(25477);
		when "0110001110000110" => data_out <= rom_array(25478);
		when "0110001110000111" => data_out <= rom_array(25479);
		when "0110001110001000" => data_out <= rom_array(25480);
		when "0110001110001001" => data_out <= rom_array(25481);
		when "0110001110001010" => data_out <= rom_array(25482);
		when "0110001110001011" => data_out <= rom_array(25483);
		when "0110001110001100" => data_out <= rom_array(25484);
		when "0110001110001101" => data_out <= rom_array(25485);
		when "0110001110001110" => data_out <= rom_array(25486);
		when "0110001110001111" => data_out <= rom_array(25487);
		when "0110001110010000" => data_out <= rom_array(25488);
		when "0110001110010001" => data_out <= rom_array(25489);
		when "0110001110010010" => data_out <= rom_array(25490);
		when "0110001110010011" => data_out <= rom_array(25491);
		when "0110001110010100" => data_out <= rom_array(25492);
		when "0110001110010101" => data_out <= rom_array(25493);
		when "0110001110010110" => data_out <= rom_array(25494);
		when "0110001110010111" => data_out <= rom_array(25495);
		when "0110001110011000" => data_out <= rom_array(25496);
		when "0110001110011001" => data_out <= rom_array(25497);
		when "0110001110011010" => data_out <= rom_array(25498);
		when "0110001110011011" => data_out <= rom_array(25499);
		when "0110001110011100" => data_out <= rom_array(25500);
		when "0110001110011101" => data_out <= rom_array(25501);
		when "0110001110011110" => data_out <= rom_array(25502);
		when "0110001110011111" => data_out <= rom_array(25503);
		when "0110001110100000" => data_out <= rom_array(25504);
		when "0110001110100001" => data_out <= rom_array(25505);
		when "0110001110100010" => data_out <= rom_array(25506);
		when "0110001110100011" => data_out <= rom_array(25507);
		when "0110001110100100" => data_out <= rom_array(25508);
		when "0110001110100101" => data_out <= rom_array(25509);
		when "0110001110100110" => data_out <= rom_array(25510);
		when "0110001110100111" => data_out <= rom_array(25511);
		when "0110001110101000" => data_out <= rom_array(25512);
		when "0110001110101001" => data_out <= rom_array(25513);
		when "0110001110101010" => data_out <= rom_array(25514);
		when "0110001110101011" => data_out <= rom_array(25515);
		when "0110001110101100" => data_out <= rom_array(25516);
		when "0110001110101101" => data_out <= rom_array(25517);
		when "0110001110101110" => data_out <= rom_array(25518);
		when "0110001110101111" => data_out <= rom_array(25519);
		when "0110001110110000" => data_out <= rom_array(25520);
		when "0110001110110001" => data_out <= rom_array(25521);
		when "0110001110110010" => data_out <= rom_array(25522);
		when "0110001110110011" => data_out <= rom_array(25523);
		when "0110001110110100" => data_out <= rom_array(25524);
		when "0110001110110101" => data_out <= rom_array(25525);
		when "0110001110110110" => data_out <= rom_array(25526);
		when "0110001110110111" => data_out <= rom_array(25527);
		when "0110001110111000" => data_out <= rom_array(25528);
		when "0110001110111001" => data_out <= rom_array(25529);
		when "0110001110111010" => data_out <= rom_array(25530);
		when "0110001110111011" => data_out <= rom_array(25531);
		when "0110001110111100" => data_out <= rom_array(25532);
		when "0110001110111101" => data_out <= rom_array(25533);
		when "0110001110111110" => data_out <= rom_array(25534);
		when "0110001110111111" => data_out <= rom_array(25535);
		when "0110001111000000" => data_out <= rom_array(25536);
		when "0110001111000001" => data_out <= rom_array(25537);
		when "0110001111000010" => data_out <= rom_array(25538);
		when "0110001111000011" => data_out <= rom_array(25539);
		when "0110001111000100" => data_out <= rom_array(25540);
		when "0110001111000101" => data_out <= rom_array(25541);
		when "0110001111000110" => data_out <= rom_array(25542);
		when "0110001111000111" => data_out <= rom_array(25543);
		when "0110001111001000" => data_out <= rom_array(25544);
		when "0110001111001001" => data_out <= rom_array(25545);
		when "0110001111001010" => data_out <= rom_array(25546);
		when "0110001111001011" => data_out <= rom_array(25547);
		when "0110001111001100" => data_out <= rom_array(25548);
		when "0110001111001101" => data_out <= rom_array(25549);
		when "0110001111001110" => data_out <= rom_array(25550);
		when "0110001111001111" => data_out <= rom_array(25551);
		when "0110001111010000" => data_out <= rom_array(25552);
		when "0110001111010001" => data_out <= rom_array(25553);
		when "0110001111010010" => data_out <= rom_array(25554);
		when "0110001111010011" => data_out <= rom_array(25555);
		when "0110001111010100" => data_out <= rom_array(25556);
		when "0110001111010101" => data_out <= rom_array(25557);
		when "0110001111010110" => data_out <= rom_array(25558);
		when "0110001111010111" => data_out <= rom_array(25559);
		when "0110001111011000" => data_out <= rom_array(25560);
		when "0110001111011001" => data_out <= rom_array(25561);
		when "0110001111011010" => data_out <= rom_array(25562);
		when "0110001111011011" => data_out <= rom_array(25563);
		when "0110001111011100" => data_out <= rom_array(25564);
		when "0110001111011101" => data_out <= rom_array(25565);
		when "0110001111011110" => data_out <= rom_array(25566);
		when "0110001111011111" => data_out <= rom_array(25567);
		when "0110001111100000" => data_out <= rom_array(25568);
		when "0110001111100001" => data_out <= rom_array(25569);
		when "0110001111100010" => data_out <= rom_array(25570);
		when "0110001111100011" => data_out <= rom_array(25571);
		when "0110001111100100" => data_out <= rom_array(25572);
		when "0110001111100101" => data_out <= rom_array(25573);
		when "0110001111100110" => data_out <= rom_array(25574);
		when "0110001111100111" => data_out <= rom_array(25575);
		when "0110001111101000" => data_out <= rom_array(25576);
		when "0110001111101001" => data_out <= rom_array(25577);
		when "0110001111101010" => data_out <= rom_array(25578);
		when "0110001111101011" => data_out <= rom_array(25579);
		when "0110001111101100" => data_out <= rom_array(25580);
		when "0110001111101101" => data_out <= rom_array(25581);
		when "0110001111101110" => data_out <= rom_array(25582);
		when "0110001111101111" => data_out <= rom_array(25583);
		when "0110001111110000" => data_out <= rom_array(25584);
		when "0110001111110001" => data_out <= rom_array(25585);
		when "0110001111110010" => data_out <= rom_array(25586);
		when "0110001111110011" => data_out <= rom_array(25587);
		when "0110001111110100" => data_out <= rom_array(25588);
		when "0110001111110101" => data_out <= rom_array(25589);
		when "0110001111110110" => data_out <= rom_array(25590);
		when "0110001111110111" => data_out <= rom_array(25591);
		when "0110001111111000" => data_out <= rom_array(25592);
		when "0110001111111001" => data_out <= rom_array(25593);
		when "0110001111111010" => data_out <= rom_array(25594);
		when "0110001111111011" => data_out <= rom_array(25595);
		when "0110001111111100" => data_out <= rom_array(25596);
		when "0110001111111101" => data_out <= rom_array(25597);
		when "0110001111111110" => data_out <= rom_array(25598);
		when "0110001111111111" => data_out <= rom_array(25599);
		when "0110010000000000" => data_out <= rom_array(25600);
		when "0110010000000001" => data_out <= rom_array(25601);
		when "0110010000000010" => data_out <= rom_array(25602);
		when "0110010000000011" => data_out <= rom_array(25603);
		when "0110010000000100" => data_out <= rom_array(25604);
		when "0110010000000101" => data_out <= rom_array(25605);
		when "0110010000000110" => data_out <= rom_array(25606);
		when "0110010000000111" => data_out <= rom_array(25607);
		when "0110010000001000" => data_out <= rom_array(25608);
		when "0110010000001001" => data_out <= rom_array(25609);
		when "0110010000001010" => data_out <= rom_array(25610);
		when "0110010000001011" => data_out <= rom_array(25611);
		when "0110010000001100" => data_out <= rom_array(25612);
		when "0110010000001101" => data_out <= rom_array(25613);
		when "0110010000001110" => data_out <= rom_array(25614);
		when "0110010000001111" => data_out <= rom_array(25615);
		when "0110010000010000" => data_out <= rom_array(25616);
		when "0110010000010001" => data_out <= rom_array(25617);
		when "0110010000010010" => data_out <= rom_array(25618);
		when "0110010000010011" => data_out <= rom_array(25619);
		when "0110010000010100" => data_out <= rom_array(25620);
		when "0110010000010101" => data_out <= rom_array(25621);
		when "0110010000010110" => data_out <= rom_array(25622);
		when "0110010000010111" => data_out <= rom_array(25623);
		when "0110010000011000" => data_out <= rom_array(25624);
		when "0110010000011001" => data_out <= rom_array(25625);
		when "0110010000011010" => data_out <= rom_array(25626);
		when "0110010000011011" => data_out <= rom_array(25627);
		when "0110010000011100" => data_out <= rom_array(25628);
		when "0110010000011101" => data_out <= rom_array(25629);
		when "0110010000011110" => data_out <= rom_array(25630);
		when "0110010000011111" => data_out <= rom_array(25631);
		when "0110010000100000" => data_out <= rom_array(25632);
		when "0110010000100001" => data_out <= rom_array(25633);
		when "0110010000100010" => data_out <= rom_array(25634);
		when "0110010000100011" => data_out <= rom_array(25635);
		when "0110010000100100" => data_out <= rom_array(25636);
		when "0110010000100101" => data_out <= rom_array(25637);
		when "0110010000100110" => data_out <= rom_array(25638);
		when "0110010000100111" => data_out <= rom_array(25639);
		when "0110010000101000" => data_out <= rom_array(25640);
		when "0110010000101001" => data_out <= rom_array(25641);
		when "0110010000101010" => data_out <= rom_array(25642);
		when "0110010000101011" => data_out <= rom_array(25643);
		when "0110010000101100" => data_out <= rom_array(25644);
		when "0110010000101101" => data_out <= rom_array(25645);
		when "0110010000101110" => data_out <= rom_array(25646);
		when "0110010000101111" => data_out <= rom_array(25647);
		when "0110010000110000" => data_out <= rom_array(25648);
		when "0110010000110001" => data_out <= rom_array(25649);
		when "0110010000110010" => data_out <= rom_array(25650);
		when "0110010000110011" => data_out <= rom_array(25651);
		when "0110010000110100" => data_out <= rom_array(25652);
		when "0110010000110101" => data_out <= rom_array(25653);
		when "0110010000110110" => data_out <= rom_array(25654);
		when "0110010000110111" => data_out <= rom_array(25655);
		when "0110010000111000" => data_out <= rom_array(25656);
		when "0110010000111001" => data_out <= rom_array(25657);
		when "0110010000111010" => data_out <= rom_array(25658);
		when "0110010000111011" => data_out <= rom_array(25659);
		when "0110010000111100" => data_out <= rom_array(25660);
		when "0110010000111101" => data_out <= rom_array(25661);
		when "0110010000111110" => data_out <= rom_array(25662);
		when "0110010000111111" => data_out <= rom_array(25663);
		when "0110010001000000" => data_out <= rom_array(25664);
		when "0110010001000001" => data_out <= rom_array(25665);
		when "0110010001000010" => data_out <= rom_array(25666);
		when "0110010001000011" => data_out <= rom_array(25667);
		when "0110010001000100" => data_out <= rom_array(25668);
		when "0110010001000101" => data_out <= rom_array(25669);
		when "0110010001000110" => data_out <= rom_array(25670);
		when "0110010001000111" => data_out <= rom_array(25671);
		when "0110010001001000" => data_out <= rom_array(25672);
		when "0110010001001001" => data_out <= rom_array(25673);
		when "0110010001001010" => data_out <= rom_array(25674);
		when "0110010001001011" => data_out <= rom_array(25675);
		when "0110010001001100" => data_out <= rom_array(25676);
		when "0110010001001101" => data_out <= rom_array(25677);
		when "0110010001001110" => data_out <= rom_array(25678);
		when "0110010001001111" => data_out <= rom_array(25679);
		when "0110010001010000" => data_out <= rom_array(25680);
		when "0110010001010001" => data_out <= rom_array(25681);
		when "0110010001010010" => data_out <= rom_array(25682);
		when "0110010001010011" => data_out <= rom_array(25683);
		when "0110010001010100" => data_out <= rom_array(25684);
		when "0110010001010101" => data_out <= rom_array(25685);
		when "0110010001010110" => data_out <= rom_array(25686);
		when "0110010001010111" => data_out <= rom_array(25687);
		when "0110010001011000" => data_out <= rom_array(25688);
		when "0110010001011001" => data_out <= rom_array(25689);
		when "0110010001011010" => data_out <= rom_array(25690);
		when "0110010001011011" => data_out <= rom_array(25691);
		when "0110010001011100" => data_out <= rom_array(25692);
		when "0110010001011101" => data_out <= rom_array(25693);
		when "0110010001011110" => data_out <= rom_array(25694);
		when "0110010001011111" => data_out <= rom_array(25695);
		when "0110010001100000" => data_out <= rom_array(25696);
		when "0110010001100001" => data_out <= rom_array(25697);
		when "0110010001100010" => data_out <= rom_array(25698);
		when "0110010001100011" => data_out <= rom_array(25699);
		when "0110010001100100" => data_out <= rom_array(25700);
		when "0110010001100101" => data_out <= rom_array(25701);
		when "0110010001100110" => data_out <= rom_array(25702);
		when "0110010001100111" => data_out <= rom_array(25703);
		when "0110010001101000" => data_out <= rom_array(25704);
		when "0110010001101001" => data_out <= rom_array(25705);
		when "0110010001101010" => data_out <= rom_array(25706);
		when "0110010001101011" => data_out <= rom_array(25707);
		when "0110010001101100" => data_out <= rom_array(25708);
		when "0110010001101101" => data_out <= rom_array(25709);
		when "0110010001101110" => data_out <= rom_array(25710);
		when "0110010001101111" => data_out <= rom_array(25711);
		when "0110010001110000" => data_out <= rom_array(25712);
		when "0110010001110001" => data_out <= rom_array(25713);
		when "0110010001110010" => data_out <= rom_array(25714);
		when "0110010001110011" => data_out <= rom_array(25715);
		when "0110010001110100" => data_out <= rom_array(25716);
		when "0110010001110101" => data_out <= rom_array(25717);
		when "0110010001110110" => data_out <= rom_array(25718);
		when "0110010001110111" => data_out <= rom_array(25719);
		when "0110010001111000" => data_out <= rom_array(25720);
		when "0110010001111001" => data_out <= rom_array(25721);
		when "0110010001111010" => data_out <= rom_array(25722);
		when "0110010001111011" => data_out <= rom_array(25723);
		when "0110010001111100" => data_out <= rom_array(25724);
		when "0110010001111101" => data_out <= rom_array(25725);
		when "0110010001111110" => data_out <= rom_array(25726);
		when "0110010001111111" => data_out <= rom_array(25727);
		when "0110010010000000" => data_out <= rom_array(25728);
		when "0110010010000001" => data_out <= rom_array(25729);
		when "0110010010000010" => data_out <= rom_array(25730);
		when "0110010010000011" => data_out <= rom_array(25731);
		when "0110010010000100" => data_out <= rom_array(25732);
		when "0110010010000101" => data_out <= rom_array(25733);
		when "0110010010000110" => data_out <= rom_array(25734);
		when "0110010010000111" => data_out <= rom_array(25735);
		when "0110010010001000" => data_out <= rom_array(25736);
		when "0110010010001001" => data_out <= rom_array(25737);
		when "0110010010001010" => data_out <= rom_array(25738);
		when "0110010010001011" => data_out <= rom_array(25739);
		when "0110010010001100" => data_out <= rom_array(25740);
		when "0110010010001101" => data_out <= rom_array(25741);
		when "0110010010001110" => data_out <= rom_array(25742);
		when "0110010010001111" => data_out <= rom_array(25743);
		when "0110010010010000" => data_out <= rom_array(25744);
		when "0110010010010001" => data_out <= rom_array(25745);
		when "0110010010010010" => data_out <= rom_array(25746);
		when "0110010010010011" => data_out <= rom_array(25747);
		when "0110010010010100" => data_out <= rom_array(25748);
		when "0110010010010101" => data_out <= rom_array(25749);
		when "0110010010010110" => data_out <= rom_array(25750);
		when "0110010010010111" => data_out <= rom_array(25751);
		when "0110010010011000" => data_out <= rom_array(25752);
		when "0110010010011001" => data_out <= rom_array(25753);
		when "0110010010011010" => data_out <= rom_array(25754);
		when "0110010010011011" => data_out <= rom_array(25755);
		when "0110010010011100" => data_out <= rom_array(25756);
		when "0110010010011101" => data_out <= rom_array(25757);
		when "0110010010011110" => data_out <= rom_array(25758);
		when "0110010010011111" => data_out <= rom_array(25759);
		when "0110010010100000" => data_out <= rom_array(25760);
		when "0110010010100001" => data_out <= rom_array(25761);
		when "0110010010100010" => data_out <= rom_array(25762);
		when "0110010010100011" => data_out <= rom_array(25763);
		when "0110010010100100" => data_out <= rom_array(25764);
		when "0110010010100101" => data_out <= rom_array(25765);
		when "0110010010100110" => data_out <= rom_array(25766);
		when "0110010010100111" => data_out <= rom_array(25767);
		when "0110010010101000" => data_out <= rom_array(25768);
		when "0110010010101001" => data_out <= rom_array(25769);
		when "0110010010101010" => data_out <= rom_array(25770);
		when "0110010010101011" => data_out <= rom_array(25771);
		when "0110010010101100" => data_out <= rom_array(25772);
		when "0110010010101101" => data_out <= rom_array(25773);
		when "0110010010101110" => data_out <= rom_array(25774);
		when "0110010010101111" => data_out <= rom_array(25775);
		when "0110010010110000" => data_out <= rom_array(25776);
		when "0110010010110001" => data_out <= rom_array(25777);
		when "0110010010110010" => data_out <= rom_array(25778);
		when "0110010010110011" => data_out <= rom_array(25779);
		when "0110010010110100" => data_out <= rom_array(25780);
		when "0110010010110101" => data_out <= rom_array(25781);
		when "0110010010110110" => data_out <= rom_array(25782);
		when "0110010010110111" => data_out <= rom_array(25783);
		when "0110010010111000" => data_out <= rom_array(25784);
		when "0110010010111001" => data_out <= rom_array(25785);
		when "0110010010111010" => data_out <= rom_array(25786);
		when "0110010010111011" => data_out <= rom_array(25787);
		when "0110010010111100" => data_out <= rom_array(25788);
		when "0110010010111101" => data_out <= rom_array(25789);
		when "0110010010111110" => data_out <= rom_array(25790);
		when "0110010010111111" => data_out <= rom_array(25791);
		when "0110010011000000" => data_out <= rom_array(25792);
		when "0110010011000001" => data_out <= rom_array(25793);
		when "0110010011000010" => data_out <= rom_array(25794);
		when "0110010011000011" => data_out <= rom_array(25795);
		when "0110010011000100" => data_out <= rom_array(25796);
		when "0110010011000101" => data_out <= rom_array(25797);
		when "0110010011000110" => data_out <= rom_array(25798);
		when "0110010011000111" => data_out <= rom_array(25799);
		when "0110010011001000" => data_out <= rom_array(25800);
		when "0110010011001001" => data_out <= rom_array(25801);
		when "0110010011001010" => data_out <= rom_array(25802);
		when "0110010011001011" => data_out <= rom_array(25803);
		when "0110010011001100" => data_out <= rom_array(25804);
		when "0110010011001101" => data_out <= rom_array(25805);
		when "0110010011001110" => data_out <= rom_array(25806);
		when "0110010011001111" => data_out <= rom_array(25807);
		when "0110010011010000" => data_out <= rom_array(25808);
		when "0110010011010001" => data_out <= rom_array(25809);
		when "0110010011010010" => data_out <= rom_array(25810);
		when "0110010011010011" => data_out <= rom_array(25811);
		when "0110010011010100" => data_out <= rom_array(25812);
		when "0110010011010101" => data_out <= rom_array(25813);
		when "0110010011010110" => data_out <= rom_array(25814);
		when "0110010011010111" => data_out <= rom_array(25815);
		when "0110010011011000" => data_out <= rom_array(25816);
		when "0110010011011001" => data_out <= rom_array(25817);
		when "0110010011011010" => data_out <= rom_array(25818);
		when "0110010011011011" => data_out <= rom_array(25819);
		when "0110010011011100" => data_out <= rom_array(25820);
		when "0110010011011101" => data_out <= rom_array(25821);
		when "0110010011011110" => data_out <= rom_array(25822);
		when "0110010011011111" => data_out <= rom_array(25823);
		when "0110010011100000" => data_out <= rom_array(25824);
		when "0110010011100001" => data_out <= rom_array(25825);
		when "0110010011100010" => data_out <= rom_array(25826);
		when "0110010011100011" => data_out <= rom_array(25827);
		when "0110010011100100" => data_out <= rom_array(25828);
		when "0110010011100101" => data_out <= rom_array(25829);
		when "0110010011100110" => data_out <= rom_array(25830);
		when "0110010011100111" => data_out <= rom_array(25831);
		when "0110010011101000" => data_out <= rom_array(25832);
		when "0110010011101001" => data_out <= rom_array(25833);
		when "0110010011101010" => data_out <= rom_array(25834);
		when "0110010011101011" => data_out <= rom_array(25835);
		when "0110010011101100" => data_out <= rom_array(25836);
		when "0110010011101101" => data_out <= rom_array(25837);
		when "0110010011101110" => data_out <= rom_array(25838);
		when "0110010011101111" => data_out <= rom_array(25839);
		when "0110010011110000" => data_out <= rom_array(25840);
		when "0110010011110001" => data_out <= rom_array(25841);
		when "0110010011110010" => data_out <= rom_array(25842);
		when "0110010011110011" => data_out <= rom_array(25843);
		when "0110010011110100" => data_out <= rom_array(25844);
		when "0110010011110101" => data_out <= rom_array(25845);
		when "0110010011110110" => data_out <= rom_array(25846);
		when "0110010011110111" => data_out <= rom_array(25847);
		when "0110010011111000" => data_out <= rom_array(25848);
		when "0110010011111001" => data_out <= rom_array(25849);
		when "0110010011111010" => data_out <= rom_array(25850);
		when "0110010011111011" => data_out <= rom_array(25851);
		when "0110010011111100" => data_out <= rom_array(25852);
		when "0110010011111101" => data_out <= rom_array(25853);
		when "0110010011111110" => data_out <= rom_array(25854);
		when "0110010011111111" => data_out <= rom_array(25855);
		when "0110010100000000" => data_out <= rom_array(25856);
		when "0110010100000001" => data_out <= rom_array(25857);
		when "0110010100000010" => data_out <= rom_array(25858);
		when "0110010100000011" => data_out <= rom_array(25859);
		when "0110010100000100" => data_out <= rom_array(25860);
		when "0110010100000101" => data_out <= rom_array(25861);
		when "0110010100000110" => data_out <= rom_array(25862);
		when "0110010100000111" => data_out <= rom_array(25863);
		when "0110010100001000" => data_out <= rom_array(25864);
		when "0110010100001001" => data_out <= rom_array(25865);
		when "0110010100001010" => data_out <= rom_array(25866);
		when "0110010100001011" => data_out <= rom_array(25867);
		when "0110010100001100" => data_out <= rom_array(25868);
		when "0110010100001101" => data_out <= rom_array(25869);
		when "0110010100001110" => data_out <= rom_array(25870);
		when "0110010100001111" => data_out <= rom_array(25871);
		when "0110010100010000" => data_out <= rom_array(25872);
		when "0110010100010001" => data_out <= rom_array(25873);
		when "0110010100010010" => data_out <= rom_array(25874);
		when "0110010100010011" => data_out <= rom_array(25875);
		when "0110010100010100" => data_out <= rom_array(25876);
		when "0110010100010101" => data_out <= rom_array(25877);
		when "0110010100010110" => data_out <= rom_array(25878);
		when "0110010100010111" => data_out <= rom_array(25879);
		when "0110010100011000" => data_out <= rom_array(25880);
		when "0110010100011001" => data_out <= rom_array(25881);
		when "0110010100011010" => data_out <= rom_array(25882);
		when "0110010100011011" => data_out <= rom_array(25883);
		when "0110010100011100" => data_out <= rom_array(25884);
		when "0110010100011101" => data_out <= rom_array(25885);
		when "0110010100011110" => data_out <= rom_array(25886);
		when "0110010100011111" => data_out <= rom_array(25887);
		when "0110010100100000" => data_out <= rom_array(25888);
		when "0110010100100001" => data_out <= rom_array(25889);
		when "0110010100100010" => data_out <= rom_array(25890);
		when "0110010100100011" => data_out <= rom_array(25891);
		when "0110010100100100" => data_out <= rom_array(25892);
		when "0110010100100101" => data_out <= rom_array(25893);
		when "0110010100100110" => data_out <= rom_array(25894);
		when "0110010100100111" => data_out <= rom_array(25895);
		when "0110010100101000" => data_out <= rom_array(25896);
		when "0110010100101001" => data_out <= rom_array(25897);
		when "0110010100101010" => data_out <= rom_array(25898);
		when "0110010100101011" => data_out <= rom_array(25899);
		when "0110010100101100" => data_out <= rom_array(25900);
		when "0110010100101101" => data_out <= rom_array(25901);
		when "0110010100101110" => data_out <= rom_array(25902);
		when "0110010100101111" => data_out <= rom_array(25903);
		when "0110010100110000" => data_out <= rom_array(25904);
		when "0110010100110001" => data_out <= rom_array(25905);
		when "0110010100110010" => data_out <= rom_array(25906);
		when "0110010100110011" => data_out <= rom_array(25907);
		when "0110010100110100" => data_out <= rom_array(25908);
		when "0110010100110101" => data_out <= rom_array(25909);
		when "0110010100110110" => data_out <= rom_array(25910);
		when "0110010100110111" => data_out <= rom_array(25911);
		when "0110010100111000" => data_out <= rom_array(25912);
		when "0110010100111001" => data_out <= rom_array(25913);
		when "0110010100111010" => data_out <= rom_array(25914);
		when "0110010100111011" => data_out <= rom_array(25915);
		when "0110010100111100" => data_out <= rom_array(25916);
		when "0110010100111101" => data_out <= rom_array(25917);
		when "0110010100111110" => data_out <= rom_array(25918);
		when "0110010100111111" => data_out <= rom_array(25919);
		when "0110010101000000" => data_out <= rom_array(25920);
		when "0110010101000001" => data_out <= rom_array(25921);
		when "0110010101000010" => data_out <= rom_array(25922);
		when "0110010101000011" => data_out <= rom_array(25923);
		when "0110010101000100" => data_out <= rom_array(25924);
		when "0110010101000101" => data_out <= rom_array(25925);
		when "0110010101000110" => data_out <= rom_array(25926);
		when "0110010101000111" => data_out <= rom_array(25927);
		when "0110010101001000" => data_out <= rom_array(25928);
		when "0110010101001001" => data_out <= rom_array(25929);
		when "0110010101001010" => data_out <= rom_array(25930);
		when "0110010101001011" => data_out <= rom_array(25931);
		when "0110010101001100" => data_out <= rom_array(25932);
		when "0110010101001101" => data_out <= rom_array(25933);
		when "0110010101001110" => data_out <= rom_array(25934);
		when "0110010101001111" => data_out <= rom_array(25935);
		when "0110010101010000" => data_out <= rom_array(25936);
		when "0110010101010001" => data_out <= rom_array(25937);
		when "0110010101010010" => data_out <= rom_array(25938);
		when "0110010101010011" => data_out <= rom_array(25939);
		when "0110010101010100" => data_out <= rom_array(25940);
		when "0110010101010101" => data_out <= rom_array(25941);
		when "0110010101010110" => data_out <= rom_array(25942);
		when "0110010101010111" => data_out <= rom_array(25943);
		when "0110010101011000" => data_out <= rom_array(25944);
		when "0110010101011001" => data_out <= rom_array(25945);
		when "0110010101011010" => data_out <= rom_array(25946);
		when "0110010101011011" => data_out <= rom_array(25947);
		when "0110010101011100" => data_out <= rom_array(25948);
		when "0110010101011101" => data_out <= rom_array(25949);
		when "0110010101011110" => data_out <= rom_array(25950);
		when "0110010101011111" => data_out <= rom_array(25951);
		when "0110010101100000" => data_out <= rom_array(25952);
		when "0110010101100001" => data_out <= rom_array(25953);
		when "0110010101100010" => data_out <= rom_array(25954);
		when "0110010101100011" => data_out <= rom_array(25955);
		when "0110010101100100" => data_out <= rom_array(25956);
		when "0110010101100101" => data_out <= rom_array(25957);
		when "0110010101100110" => data_out <= rom_array(25958);
		when "0110010101100111" => data_out <= rom_array(25959);
		when "0110010101101000" => data_out <= rom_array(25960);
		when "0110010101101001" => data_out <= rom_array(25961);
		when "0110010101101010" => data_out <= rom_array(25962);
		when "0110010101101011" => data_out <= rom_array(25963);
		when "0110010101101100" => data_out <= rom_array(25964);
		when "0110010101101101" => data_out <= rom_array(25965);
		when "0110010101101110" => data_out <= rom_array(25966);
		when "0110010101101111" => data_out <= rom_array(25967);
		when "0110010101110000" => data_out <= rom_array(25968);
		when "0110010101110001" => data_out <= rom_array(25969);
		when "0110010101110010" => data_out <= rom_array(25970);
		when "0110010101110011" => data_out <= rom_array(25971);
		when "0110010101110100" => data_out <= rom_array(25972);
		when "0110010101110101" => data_out <= rom_array(25973);
		when "0110010101110110" => data_out <= rom_array(25974);
		when "0110010101110111" => data_out <= rom_array(25975);
		when "0110010101111000" => data_out <= rom_array(25976);
		when "0110010101111001" => data_out <= rom_array(25977);
		when "0110010101111010" => data_out <= rom_array(25978);
		when "0110010101111011" => data_out <= rom_array(25979);
		when "0110010101111100" => data_out <= rom_array(25980);
		when "0110010101111101" => data_out <= rom_array(25981);
		when "0110010101111110" => data_out <= rom_array(25982);
		when "0110010101111111" => data_out <= rom_array(25983);
		when "0110010110000000" => data_out <= rom_array(25984);
		when "0110010110000001" => data_out <= rom_array(25985);
		when "0110010110000010" => data_out <= rom_array(25986);
		when "0110010110000011" => data_out <= rom_array(25987);
		when "0110010110000100" => data_out <= rom_array(25988);
		when "0110010110000101" => data_out <= rom_array(25989);
		when "0110010110000110" => data_out <= rom_array(25990);
		when "0110010110000111" => data_out <= rom_array(25991);
		when "0110010110001000" => data_out <= rom_array(25992);
		when "0110010110001001" => data_out <= rom_array(25993);
		when "0110010110001010" => data_out <= rom_array(25994);
		when "0110010110001011" => data_out <= rom_array(25995);
		when "0110010110001100" => data_out <= rom_array(25996);
		when "0110010110001101" => data_out <= rom_array(25997);
		when "0110010110001110" => data_out <= rom_array(25998);
		when "0110010110001111" => data_out <= rom_array(25999);
		when "0110010110010000" => data_out <= rom_array(26000);
		when "0110010110010001" => data_out <= rom_array(26001);
		when "0110010110010010" => data_out <= rom_array(26002);
		when "0110010110010011" => data_out <= rom_array(26003);
		when "0110010110010100" => data_out <= rom_array(26004);
		when "0110010110010101" => data_out <= rom_array(26005);
		when "0110010110010110" => data_out <= rom_array(26006);
		when "0110010110010111" => data_out <= rom_array(26007);
		when "0110010110011000" => data_out <= rom_array(26008);
		when "0110010110011001" => data_out <= rom_array(26009);
		when "0110010110011010" => data_out <= rom_array(26010);
		when "0110010110011011" => data_out <= rom_array(26011);
		when "0110010110011100" => data_out <= rom_array(26012);
		when "0110010110011101" => data_out <= rom_array(26013);
		when "0110010110011110" => data_out <= rom_array(26014);
		when "0110010110011111" => data_out <= rom_array(26015);
		when "0110010110100000" => data_out <= rom_array(26016);
		when "0110010110100001" => data_out <= rom_array(26017);
		when "0110010110100010" => data_out <= rom_array(26018);
		when "0110010110100011" => data_out <= rom_array(26019);
		when "0110010110100100" => data_out <= rom_array(26020);
		when "0110010110100101" => data_out <= rom_array(26021);
		when "0110010110100110" => data_out <= rom_array(26022);
		when "0110010110100111" => data_out <= rom_array(26023);
		when "0110010110101000" => data_out <= rom_array(26024);
		when "0110010110101001" => data_out <= rom_array(26025);
		when "0110010110101010" => data_out <= rom_array(26026);
		when "0110010110101011" => data_out <= rom_array(26027);
		when "0110010110101100" => data_out <= rom_array(26028);
		when "0110010110101101" => data_out <= rom_array(26029);
		when "0110010110101110" => data_out <= rom_array(26030);
		when "0110010110101111" => data_out <= rom_array(26031);
		when "0110010110110000" => data_out <= rom_array(26032);
		when "0110010110110001" => data_out <= rom_array(26033);
		when "0110010110110010" => data_out <= rom_array(26034);
		when "0110010110110011" => data_out <= rom_array(26035);
		when "0110010110110100" => data_out <= rom_array(26036);
		when "0110010110110101" => data_out <= rom_array(26037);
		when "0110010110110110" => data_out <= rom_array(26038);
		when "0110010110110111" => data_out <= rom_array(26039);
		when "0110010110111000" => data_out <= rom_array(26040);
		when "0110010110111001" => data_out <= rom_array(26041);
		when "0110010110111010" => data_out <= rom_array(26042);
		when "0110010110111011" => data_out <= rom_array(26043);
		when "0110010110111100" => data_out <= rom_array(26044);
		when "0110010110111101" => data_out <= rom_array(26045);
		when "0110010110111110" => data_out <= rom_array(26046);
		when "0110010110111111" => data_out <= rom_array(26047);
		when "0110010111000000" => data_out <= rom_array(26048);
		when "0110010111000001" => data_out <= rom_array(26049);
		when "0110010111000010" => data_out <= rom_array(26050);
		when "0110010111000011" => data_out <= rom_array(26051);
		when "0110010111000100" => data_out <= rom_array(26052);
		when "0110010111000101" => data_out <= rom_array(26053);
		when "0110010111000110" => data_out <= rom_array(26054);
		when "0110010111000111" => data_out <= rom_array(26055);
		when "0110010111001000" => data_out <= rom_array(26056);
		when "0110010111001001" => data_out <= rom_array(26057);
		when "0110010111001010" => data_out <= rom_array(26058);
		when "0110010111001011" => data_out <= rom_array(26059);
		when "0110010111001100" => data_out <= rom_array(26060);
		when "0110010111001101" => data_out <= rom_array(26061);
		when "0110010111001110" => data_out <= rom_array(26062);
		when "0110010111001111" => data_out <= rom_array(26063);
		when "0110010111010000" => data_out <= rom_array(26064);
		when "0110010111010001" => data_out <= rom_array(26065);
		when "0110010111010010" => data_out <= rom_array(26066);
		when "0110010111010011" => data_out <= rom_array(26067);
		when "0110010111010100" => data_out <= rom_array(26068);
		when "0110010111010101" => data_out <= rom_array(26069);
		when "0110010111010110" => data_out <= rom_array(26070);
		when "0110010111010111" => data_out <= rom_array(26071);
		when "0110010111011000" => data_out <= rom_array(26072);
		when "0110010111011001" => data_out <= rom_array(26073);
		when "0110010111011010" => data_out <= rom_array(26074);
		when "0110010111011011" => data_out <= rom_array(26075);
		when "0110010111011100" => data_out <= rom_array(26076);
		when "0110010111011101" => data_out <= rom_array(26077);
		when "0110010111011110" => data_out <= rom_array(26078);
		when "0110010111011111" => data_out <= rom_array(26079);
		when "0110010111100000" => data_out <= rom_array(26080);
		when "0110010111100001" => data_out <= rom_array(26081);
		when "0110010111100010" => data_out <= rom_array(26082);
		when "0110010111100011" => data_out <= rom_array(26083);
		when "0110010111100100" => data_out <= rom_array(26084);
		when "0110010111100101" => data_out <= rom_array(26085);
		when "0110010111100110" => data_out <= rom_array(26086);
		when "0110010111100111" => data_out <= rom_array(26087);
		when "0110010111101000" => data_out <= rom_array(26088);
		when "0110010111101001" => data_out <= rom_array(26089);
		when "0110010111101010" => data_out <= rom_array(26090);
		when "0110010111101011" => data_out <= rom_array(26091);
		when "0110010111101100" => data_out <= rom_array(26092);
		when "0110010111101101" => data_out <= rom_array(26093);
		when "0110010111101110" => data_out <= rom_array(26094);
		when "0110010111101111" => data_out <= rom_array(26095);
		when "0110010111110000" => data_out <= rom_array(26096);
		when "0110010111110001" => data_out <= rom_array(26097);
		when "0110010111110010" => data_out <= rom_array(26098);
		when "0110010111110011" => data_out <= rom_array(26099);
		when "0110010111110100" => data_out <= rom_array(26100);
		when "0110010111110101" => data_out <= rom_array(26101);
		when "0110010111110110" => data_out <= rom_array(26102);
		when "0110010111110111" => data_out <= rom_array(26103);
		when "0110010111111000" => data_out <= rom_array(26104);
		when "0110010111111001" => data_out <= rom_array(26105);
		when "0110010111111010" => data_out <= rom_array(26106);
		when "0110010111111011" => data_out <= rom_array(26107);
		when "0110010111111100" => data_out <= rom_array(26108);
		when "0110010111111101" => data_out <= rom_array(26109);
		when "0110010111111110" => data_out <= rom_array(26110);
		when "0110010111111111" => data_out <= rom_array(26111);
		when "0110011000000000" => data_out <= rom_array(26112);
		when "0110011000000001" => data_out <= rom_array(26113);
		when "0110011000000010" => data_out <= rom_array(26114);
		when "0110011000000011" => data_out <= rom_array(26115);
		when "0110011000000100" => data_out <= rom_array(26116);
		when "0110011000000101" => data_out <= rom_array(26117);
		when "0110011000000110" => data_out <= rom_array(26118);
		when "0110011000000111" => data_out <= rom_array(26119);
		when "0110011000001000" => data_out <= rom_array(26120);
		when "0110011000001001" => data_out <= rom_array(26121);
		when "0110011000001010" => data_out <= rom_array(26122);
		when "0110011000001011" => data_out <= rom_array(26123);
		when "0110011000001100" => data_out <= rom_array(26124);
		when "0110011000001101" => data_out <= rom_array(26125);
		when "0110011000001110" => data_out <= rom_array(26126);
		when "0110011000001111" => data_out <= rom_array(26127);
		when "0110011000010000" => data_out <= rom_array(26128);
		when "0110011000010001" => data_out <= rom_array(26129);
		when "0110011000010010" => data_out <= rom_array(26130);
		when "0110011000010011" => data_out <= rom_array(26131);
		when "0110011000010100" => data_out <= rom_array(26132);
		when "0110011000010101" => data_out <= rom_array(26133);
		when "0110011000010110" => data_out <= rom_array(26134);
		when "0110011000010111" => data_out <= rom_array(26135);
		when "0110011000011000" => data_out <= rom_array(26136);
		when "0110011000011001" => data_out <= rom_array(26137);
		when "0110011000011010" => data_out <= rom_array(26138);
		when "0110011000011011" => data_out <= rom_array(26139);
		when "0110011000011100" => data_out <= rom_array(26140);
		when "0110011000011101" => data_out <= rom_array(26141);
		when "0110011000011110" => data_out <= rom_array(26142);
		when "0110011000011111" => data_out <= rom_array(26143);
		when "0110011000100000" => data_out <= rom_array(26144);
		when "0110011000100001" => data_out <= rom_array(26145);
		when "0110011000100010" => data_out <= rom_array(26146);
		when "0110011000100011" => data_out <= rom_array(26147);
		when "0110011000100100" => data_out <= rom_array(26148);
		when "0110011000100101" => data_out <= rom_array(26149);
		when "0110011000100110" => data_out <= rom_array(26150);
		when "0110011000100111" => data_out <= rom_array(26151);
		when "0110011000101000" => data_out <= rom_array(26152);
		when "0110011000101001" => data_out <= rom_array(26153);
		when "0110011000101010" => data_out <= rom_array(26154);
		when "0110011000101011" => data_out <= rom_array(26155);
		when "0110011000101100" => data_out <= rom_array(26156);
		when "0110011000101101" => data_out <= rom_array(26157);
		when "0110011000101110" => data_out <= rom_array(26158);
		when "0110011000101111" => data_out <= rom_array(26159);
		when "0110011000110000" => data_out <= rom_array(26160);
		when "0110011000110001" => data_out <= rom_array(26161);
		when "0110011000110010" => data_out <= rom_array(26162);
		when "0110011000110011" => data_out <= rom_array(26163);
		when "0110011000110100" => data_out <= rom_array(26164);
		when "0110011000110101" => data_out <= rom_array(26165);
		when "0110011000110110" => data_out <= rom_array(26166);
		when "0110011000110111" => data_out <= rom_array(26167);
		when "0110011000111000" => data_out <= rom_array(26168);
		when "0110011000111001" => data_out <= rom_array(26169);
		when "0110011000111010" => data_out <= rom_array(26170);
		when "0110011000111011" => data_out <= rom_array(26171);
		when "0110011000111100" => data_out <= rom_array(26172);
		when "0110011000111101" => data_out <= rom_array(26173);
		when "0110011000111110" => data_out <= rom_array(26174);
		when "0110011000111111" => data_out <= rom_array(26175);
		when "0110011001000000" => data_out <= rom_array(26176);
		when "0110011001000001" => data_out <= rom_array(26177);
		when "0110011001000010" => data_out <= rom_array(26178);
		when "0110011001000011" => data_out <= rom_array(26179);
		when "0110011001000100" => data_out <= rom_array(26180);
		when "0110011001000101" => data_out <= rom_array(26181);
		when "0110011001000110" => data_out <= rom_array(26182);
		when "0110011001000111" => data_out <= rom_array(26183);
		when "0110011001001000" => data_out <= rom_array(26184);
		when "0110011001001001" => data_out <= rom_array(26185);
		when "0110011001001010" => data_out <= rom_array(26186);
		when "0110011001001011" => data_out <= rom_array(26187);
		when "0110011001001100" => data_out <= rom_array(26188);
		when "0110011001001101" => data_out <= rom_array(26189);
		when "0110011001001110" => data_out <= rom_array(26190);
		when "0110011001001111" => data_out <= rom_array(26191);
		when "0110011001010000" => data_out <= rom_array(26192);
		when "0110011001010001" => data_out <= rom_array(26193);
		when "0110011001010010" => data_out <= rom_array(26194);
		when "0110011001010011" => data_out <= rom_array(26195);
		when "0110011001010100" => data_out <= rom_array(26196);
		when "0110011001010101" => data_out <= rom_array(26197);
		when "0110011001010110" => data_out <= rom_array(26198);
		when "0110011001010111" => data_out <= rom_array(26199);
		when "0110011001011000" => data_out <= rom_array(26200);
		when "0110011001011001" => data_out <= rom_array(26201);
		when "0110011001011010" => data_out <= rom_array(26202);
		when "0110011001011011" => data_out <= rom_array(26203);
		when "0110011001011100" => data_out <= rom_array(26204);
		when "0110011001011101" => data_out <= rom_array(26205);
		when "0110011001011110" => data_out <= rom_array(26206);
		when "0110011001011111" => data_out <= rom_array(26207);
		when "0110011001100000" => data_out <= rom_array(26208);
		when "0110011001100001" => data_out <= rom_array(26209);
		when "0110011001100010" => data_out <= rom_array(26210);
		when "0110011001100011" => data_out <= rom_array(26211);
		when "0110011001100100" => data_out <= rom_array(26212);
		when "0110011001100101" => data_out <= rom_array(26213);
		when "0110011001100110" => data_out <= rom_array(26214);
		when "0110011001100111" => data_out <= rom_array(26215);
		when "0110011001101000" => data_out <= rom_array(26216);
		when "0110011001101001" => data_out <= rom_array(26217);
		when "0110011001101010" => data_out <= rom_array(26218);
		when "0110011001101011" => data_out <= rom_array(26219);
		when "0110011001101100" => data_out <= rom_array(26220);
		when "0110011001101101" => data_out <= rom_array(26221);
		when "0110011001101110" => data_out <= rom_array(26222);
		when "0110011001101111" => data_out <= rom_array(26223);
		when "0110011001110000" => data_out <= rom_array(26224);
		when "0110011001110001" => data_out <= rom_array(26225);
		when "0110011001110010" => data_out <= rom_array(26226);
		when "0110011001110011" => data_out <= rom_array(26227);
		when "0110011001110100" => data_out <= rom_array(26228);
		when "0110011001110101" => data_out <= rom_array(26229);
		when "0110011001110110" => data_out <= rom_array(26230);
		when "0110011001110111" => data_out <= rom_array(26231);
		when "0110011001111000" => data_out <= rom_array(26232);
		when "0110011001111001" => data_out <= rom_array(26233);
		when "0110011001111010" => data_out <= rom_array(26234);
		when "0110011001111011" => data_out <= rom_array(26235);
		when "0110011001111100" => data_out <= rom_array(26236);
		when "0110011001111101" => data_out <= rom_array(26237);
		when "0110011001111110" => data_out <= rom_array(26238);
		when "0110011001111111" => data_out <= rom_array(26239);
		when "0110011010000000" => data_out <= rom_array(26240);
		when "0110011010000001" => data_out <= rom_array(26241);
		when "0110011010000010" => data_out <= rom_array(26242);
		when "0110011010000011" => data_out <= rom_array(26243);
		when "0110011010000100" => data_out <= rom_array(26244);
		when "0110011010000101" => data_out <= rom_array(26245);
		when "0110011010000110" => data_out <= rom_array(26246);
		when "0110011010000111" => data_out <= rom_array(26247);
		when "0110011010001000" => data_out <= rom_array(26248);
		when "0110011010001001" => data_out <= rom_array(26249);
		when "0110011010001010" => data_out <= rom_array(26250);
		when "0110011010001011" => data_out <= rom_array(26251);
		when "0110011010001100" => data_out <= rom_array(26252);
		when "0110011010001101" => data_out <= rom_array(26253);
		when "0110011010001110" => data_out <= rom_array(26254);
		when "0110011010001111" => data_out <= rom_array(26255);
		when "0110011010010000" => data_out <= rom_array(26256);
		when "0110011010010001" => data_out <= rom_array(26257);
		when "0110011010010010" => data_out <= rom_array(26258);
		when "0110011010010011" => data_out <= rom_array(26259);
		when "0110011010010100" => data_out <= rom_array(26260);
		when "0110011010010101" => data_out <= rom_array(26261);
		when "0110011010010110" => data_out <= rom_array(26262);
		when "0110011010010111" => data_out <= rom_array(26263);
		when "0110011010011000" => data_out <= rom_array(26264);
		when "0110011010011001" => data_out <= rom_array(26265);
		when "0110011010011010" => data_out <= rom_array(26266);
		when "0110011010011011" => data_out <= rom_array(26267);
		when "0110011010011100" => data_out <= rom_array(26268);
		when "0110011010011101" => data_out <= rom_array(26269);
		when "0110011010011110" => data_out <= rom_array(26270);
		when "0110011010011111" => data_out <= rom_array(26271);
		when "0110011010100000" => data_out <= rom_array(26272);
		when "0110011010100001" => data_out <= rom_array(26273);
		when "0110011010100010" => data_out <= rom_array(26274);
		when "0110011010100011" => data_out <= rom_array(26275);
		when "0110011010100100" => data_out <= rom_array(26276);
		when "0110011010100101" => data_out <= rom_array(26277);
		when "0110011010100110" => data_out <= rom_array(26278);
		when "0110011010100111" => data_out <= rom_array(26279);
		when "0110011010101000" => data_out <= rom_array(26280);
		when "0110011010101001" => data_out <= rom_array(26281);
		when "0110011010101010" => data_out <= rom_array(26282);
		when "0110011010101011" => data_out <= rom_array(26283);
		when "0110011010101100" => data_out <= rom_array(26284);
		when "0110011010101101" => data_out <= rom_array(26285);
		when "0110011010101110" => data_out <= rom_array(26286);
		when "0110011010101111" => data_out <= rom_array(26287);
		when "0110011010110000" => data_out <= rom_array(26288);
		when "0110011010110001" => data_out <= rom_array(26289);
		when "0110011010110010" => data_out <= rom_array(26290);
		when "0110011010110011" => data_out <= rom_array(26291);
		when "0110011010110100" => data_out <= rom_array(26292);
		when "0110011010110101" => data_out <= rom_array(26293);
		when "0110011010110110" => data_out <= rom_array(26294);
		when "0110011010110111" => data_out <= rom_array(26295);
		when "0110011010111000" => data_out <= rom_array(26296);
		when "0110011010111001" => data_out <= rom_array(26297);
		when "0110011010111010" => data_out <= rom_array(26298);
		when "0110011010111011" => data_out <= rom_array(26299);
		when "0110011010111100" => data_out <= rom_array(26300);
		when "0110011010111101" => data_out <= rom_array(26301);
		when "0110011010111110" => data_out <= rom_array(26302);
		when "0110011010111111" => data_out <= rom_array(26303);
		when "0110011011000000" => data_out <= rom_array(26304);
		when "0110011011000001" => data_out <= rom_array(26305);
		when "0110011011000010" => data_out <= rom_array(26306);
		when "0110011011000011" => data_out <= rom_array(26307);
		when "0110011011000100" => data_out <= rom_array(26308);
		when "0110011011000101" => data_out <= rom_array(26309);
		when "0110011011000110" => data_out <= rom_array(26310);
		when "0110011011000111" => data_out <= rom_array(26311);
		when "0110011011001000" => data_out <= rom_array(26312);
		when "0110011011001001" => data_out <= rom_array(26313);
		when "0110011011001010" => data_out <= rom_array(26314);
		when "0110011011001011" => data_out <= rom_array(26315);
		when "0110011011001100" => data_out <= rom_array(26316);
		when "0110011011001101" => data_out <= rom_array(26317);
		when "0110011011001110" => data_out <= rom_array(26318);
		when "0110011011001111" => data_out <= rom_array(26319);
		when "0110011011010000" => data_out <= rom_array(26320);
		when "0110011011010001" => data_out <= rom_array(26321);
		when "0110011011010010" => data_out <= rom_array(26322);
		when "0110011011010011" => data_out <= rom_array(26323);
		when "0110011011010100" => data_out <= rom_array(26324);
		when "0110011011010101" => data_out <= rom_array(26325);
		when "0110011011010110" => data_out <= rom_array(26326);
		when "0110011011010111" => data_out <= rom_array(26327);
		when "0110011011011000" => data_out <= rom_array(26328);
		when "0110011011011001" => data_out <= rom_array(26329);
		when "0110011011011010" => data_out <= rom_array(26330);
		when "0110011011011011" => data_out <= rom_array(26331);
		when "0110011011011100" => data_out <= rom_array(26332);
		when "0110011011011101" => data_out <= rom_array(26333);
		when "0110011011011110" => data_out <= rom_array(26334);
		when "0110011011011111" => data_out <= rom_array(26335);
		when "0110011011100000" => data_out <= rom_array(26336);
		when "0110011011100001" => data_out <= rom_array(26337);
		when "0110011011100010" => data_out <= rom_array(26338);
		when "0110011011100011" => data_out <= rom_array(26339);
		when "0110011011100100" => data_out <= rom_array(26340);
		when "0110011011100101" => data_out <= rom_array(26341);
		when "0110011011100110" => data_out <= rom_array(26342);
		when "0110011011100111" => data_out <= rom_array(26343);
		when "0110011011101000" => data_out <= rom_array(26344);
		when "0110011011101001" => data_out <= rom_array(26345);
		when "0110011011101010" => data_out <= rom_array(26346);
		when "0110011011101011" => data_out <= rom_array(26347);
		when "0110011011101100" => data_out <= rom_array(26348);
		when "0110011011101101" => data_out <= rom_array(26349);
		when "0110011011101110" => data_out <= rom_array(26350);
		when "0110011011101111" => data_out <= rom_array(26351);
		when "0110011011110000" => data_out <= rom_array(26352);
		when "0110011011110001" => data_out <= rom_array(26353);
		when "0110011011110010" => data_out <= rom_array(26354);
		when "0110011011110011" => data_out <= rom_array(26355);
		when "0110011011110100" => data_out <= rom_array(26356);
		when "0110011011110101" => data_out <= rom_array(26357);
		when "0110011011110110" => data_out <= rom_array(26358);
		when "0110011011110111" => data_out <= rom_array(26359);
		when "0110011011111000" => data_out <= rom_array(26360);
		when "0110011011111001" => data_out <= rom_array(26361);
		when "0110011011111010" => data_out <= rom_array(26362);
		when "0110011011111011" => data_out <= rom_array(26363);
		when "0110011011111100" => data_out <= rom_array(26364);
		when "0110011011111101" => data_out <= rom_array(26365);
		when "0110011011111110" => data_out <= rom_array(26366);
		when "0110011011111111" => data_out <= rom_array(26367);
		when "0110011100000000" => data_out <= rom_array(26368);
		when "0110011100000001" => data_out <= rom_array(26369);
		when "0110011100000010" => data_out <= rom_array(26370);
		when "0110011100000011" => data_out <= rom_array(26371);
		when "0110011100000100" => data_out <= rom_array(26372);
		when "0110011100000101" => data_out <= rom_array(26373);
		when "0110011100000110" => data_out <= rom_array(26374);
		when "0110011100000111" => data_out <= rom_array(26375);
		when "0110011100001000" => data_out <= rom_array(26376);
		when "0110011100001001" => data_out <= rom_array(26377);
		when "0110011100001010" => data_out <= rom_array(26378);
		when "0110011100001011" => data_out <= rom_array(26379);
		when "0110011100001100" => data_out <= rom_array(26380);
		when "0110011100001101" => data_out <= rom_array(26381);
		when "0110011100001110" => data_out <= rom_array(26382);
		when "0110011100001111" => data_out <= rom_array(26383);
		when "0110011100010000" => data_out <= rom_array(26384);
		when "0110011100010001" => data_out <= rom_array(26385);
		when "0110011100010010" => data_out <= rom_array(26386);
		when "0110011100010011" => data_out <= rom_array(26387);
		when "0110011100010100" => data_out <= rom_array(26388);
		when "0110011100010101" => data_out <= rom_array(26389);
		when "0110011100010110" => data_out <= rom_array(26390);
		when "0110011100010111" => data_out <= rom_array(26391);
		when "0110011100011000" => data_out <= rom_array(26392);
		when "0110011100011001" => data_out <= rom_array(26393);
		when "0110011100011010" => data_out <= rom_array(26394);
		when "0110011100011011" => data_out <= rom_array(26395);
		when "0110011100011100" => data_out <= rom_array(26396);
		when "0110011100011101" => data_out <= rom_array(26397);
		when "0110011100011110" => data_out <= rom_array(26398);
		when "0110011100011111" => data_out <= rom_array(26399);
		when "0110011100100000" => data_out <= rom_array(26400);
		when "0110011100100001" => data_out <= rom_array(26401);
		when "0110011100100010" => data_out <= rom_array(26402);
		when "0110011100100011" => data_out <= rom_array(26403);
		when "0110011100100100" => data_out <= rom_array(26404);
		when "0110011100100101" => data_out <= rom_array(26405);
		when "0110011100100110" => data_out <= rom_array(26406);
		when "0110011100100111" => data_out <= rom_array(26407);
		when "0110011100101000" => data_out <= rom_array(26408);
		when "0110011100101001" => data_out <= rom_array(26409);
		when "0110011100101010" => data_out <= rom_array(26410);
		when "0110011100101011" => data_out <= rom_array(26411);
		when "0110011100101100" => data_out <= rom_array(26412);
		when "0110011100101101" => data_out <= rom_array(26413);
		when "0110011100101110" => data_out <= rom_array(26414);
		when "0110011100101111" => data_out <= rom_array(26415);
		when "0110011100110000" => data_out <= rom_array(26416);
		when "0110011100110001" => data_out <= rom_array(26417);
		when "0110011100110010" => data_out <= rom_array(26418);
		when "0110011100110011" => data_out <= rom_array(26419);
		when "0110011100110100" => data_out <= rom_array(26420);
		when "0110011100110101" => data_out <= rom_array(26421);
		when "0110011100110110" => data_out <= rom_array(26422);
		when "0110011100110111" => data_out <= rom_array(26423);
		when "0110011100111000" => data_out <= rom_array(26424);
		when "0110011100111001" => data_out <= rom_array(26425);
		when "0110011100111010" => data_out <= rom_array(26426);
		when "0110011100111011" => data_out <= rom_array(26427);
		when "0110011100111100" => data_out <= rom_array(26428);
		when "0110011100111101" => data_out <= rom_array(26429);
		when "0110011100111110" => data_out <= rom_array(26430);
		when "0110011100111111" => data_out <= rom_array(26431);
		when "0110011101000000" => data_out <= rom_array(26432);
		when "0110011101000001" => data_out <= rom_array(26433);
		when "0110011101000010" => data_out <= rom_array(26434);
		when "0110011101000011" => data_out <= rom_array(26435);
		when "0110011101000100" => data_out <= rom_array(26436);
		when "0110011101000101" => data_out <= rom_array(26437);
		when "0110011101000110" => data_out <= rom_array(26438);
		when "0110011101000111" => data_out <= rom_array(26439);
		when "0110011101001000" => data_out <= rom_array(26440);
		when "0110011101001001" => data_out <= rom_array(26441);
		when "0110011101001010" => data_out <= rom_array(26442);
		when "0110011101001011" => data_out <= rom_array(26443);
		when "0110011101001100" => data_out <= rom_array(26444);
		when "0110011101001101" => data_out <= rom_array(26445);
		when "0110011101001110" => data_out <= rom_array(26446);
		when "0110011101001111" => data_out <= rom_array(26447);
		when "0110011101010000" => data_out <= rom_array(26448);
		when "0110011101010001" => data_out <= rom_array(26449);
		when "0110011101010010" => data_out <= rom_array(26450);
		when "0110011101010011" => data_out <= rom_array(26451);
		when "0110011101010100" => data_out <= rom_array(26452);
		when "0110011101010101" => data_out <= rom_array(26453);
		when "0110011101010110" => data_out <= rom_array(26454);
		when "0110011101010111" => data_out <= rom_array(26455);
		when "0110011101011000" => data_out <= rom_array(26456);
		when "0110011101011001" => data_out <= rom_array(26457);
		when "0110011101011010" => data_out <= rom_array(26458);
		when "0110011101011011" => data_out <= rom_array(26459);
		when "0110011101011100" => data_out <= rom_array(26460);
		when "0110011101011101" => data_out <= rom_array(26461);
		when "0110011101011110" => data_out <= rom_array(26462);
		when "0110011101011111" => data_out <= rom_array(26463);
		when "0110011101100000" => data_out <= rom_array(26464);
		when "0110011101100001" => data_out <= rom_array(26465);
		when "0110011101100010" => data_out <= rom_array(26466);
		when "0110011101100011" => data_out <= rom_array(26467);
		when "0110011101100100" => data_out <= rom_array(26468);
		when "0110011101100101" => data_out <= rom_array(26469);
		when "0110011101100110" => data_out <= rom_array(26470);
		when "0110011101100111" => data_out <= rom_array(26471);
		when "0110011101101000" => data_out <= rom_array(26472);
		when "0110011101101001" => data_out <= rom_array(26473);
		when "0110011101101010" => data_out <= rom_array(26474);
		when "0110011101101011" => data_out <= rom_array(26475);
		when "0110011101101100" => data_out <= rom_array(26476);
		when "0110011101101101" => data_out <= rom_array(26477);
		when "0110011101101110" => data_out <= rom_array(26478);
		when "0110011101101111" => data_out <= rom_array(26479);
		when "0110011101110000" => data_out <= rom_array(26480);
		when "0110011101110001" => data_out <= rom_array(26481);
		when "0110011101110010" => data_out <= rom_array(26482);
		when "0110011101110011" => data_out <= rom_array(26483);
		when "0110011101110100" => data_out <= rom_array(26484);
		when "0110011101110101" => data_out <= rom_array(26485);
		when "0110011101110110" => data_out <= rom_array(26486);
		when "0110011101110111" => data_out <= rom_array(26487);
		when "0110011101111000" => data_out <= rom_array(26488);
		when "0110011101111001" => data_out <= rom_array(26489);
		when "0110011101111010" => data_out <= rom_array(26490);
		when "0110011101111011" => data_out <= rom_array(26491);
		when "0110011101111100" => data_out <= rom_array(26492);
		when "0110011101111101" => data_out <= rom_array(26493);
		when "0110011101111110" => data_out <= rom_array(26494);
		when "0110011101111111" => data_out <= rom_array(26495);
		when "0110011110000000" => data_out <= rom_array(26496);
		when "0110011110000001" => data_out <= rom_array(26497);
		when "0110011110000010" => data_out <= rom_array(26498);
		when "0110011110000011" => data_out <= rom_array(26499);
		when "0110011110000100" => data_out <= rom_array(26500);
		when "0110011110000101" => data_out <= rom_array(26501);
		when "0110011110000110" => data_out <= rom_array(26502);
		when "0110011110000111" => data_out <= rom_array(26503);
		when "0110011110001000" => data_out <= rom_array(26504);
		when "0110011110001001" => data_out <= rom_array(26505);
		when "0110011110001010" => data_out <= rom_array(26506);
		when "0110011110001011" => data_out <= rom_array(26507);
		when "0110011110001100" => data_out <= rom_array(26508);
		when "0110011110001101" => data_out <= rom_array(26509);
		when "0110011110001110" => data_out <= rom_array(26510);
		when "0110011110001111" => data_out <= rom_array(26511);
		when "0110011110010000" => data_out <= rom_array(26512);
		when "0110011110010001" => data_out <= rom_array(26513);
		when "0110011110010010" => data_out <= rom_array(26514);
		when "0110011110010011" => data_out <= rom_array(26515);
		when "0110011110010100" => data_out <= rom_array(26516);
		when "0110011110010101" => data_out <= rom_array(26517);
		when "0110011110010110" => data_out <= rom_array(26518);
		when "0110011110010111" => data_out <= rom_array(26519);
		when "0110011110011000" => data_out <= rom_array(26520);
		when "0110011110011001" => data_out <= rom_array(26521);
		when "0110011110011010" => data_out <= rom_array(26522);
		when "0110011110011011" => data_out <= rom_array(26523);
		when "0110011110011100" => data_out <= rom_array(26524);
		when "0110011110011101" => data_out <= rom_array(26525);
		when "0110011110011110" => data_out <= rom_array(26526);
		when "0110011110011111" => data_out <= rom_array(26527);
		when "0110011110100000" => data_out <= rom_array(26528);
		when "0110011110100001" => data_out <= rom_array(26529);
		when "0110011110100010" => data_out <= rom_array(26530);
		when "0110011110100011" => data_out <= rom_array(26531);
		when "0110011110100100" => data_out <= rom_array(26532);
		when "0110011110100101" => data_out <= rom_array(26533);
		when "0110011110100110" => data_out <= rom_array(26534);
		when "0110011110100111" => data_out <= rom_array(26535);
		when "0110011110101000" => data_out <= rom_array(26536);
		when "0110011110101001" => data_out <= rom_array(26537);
		when "0110011110101010" => data_out <= rom_array(26538);
		when "0110011110101011" => data_out <= rom_array(26539);
		when "0110011110101100" => data_out <= rom_array(26540);
		when "0110011110101101" => data_out <= rom_array(26541);
		when "0110011110101110" => data_out <= rom_array(26542);
		when "0110011110101111" => data_out <= rom_array(26543);
		when "0110011110110000" => data_out <= rom_array(26544);
		when "0110011110110001" => data_out <= rom_array(26545);
		when "0110011110110010" => data_out <= rom_array(26546);
		when "0110011110110011" => data_out <= rom_array(26547);
		when "0110011110110100" => data_out <= rom_array(26548);
		when "0110011110110101" => data_out <= rom_array(26549);
		when "0110011110110110" => data_out <= rom_array(26550);
		when "0110011110110111" => data_out <= rom_array(26551);
		when "0110011110111000" => data_out <= rom_array(26552);
		when "0110011110111001" => data_out <= rom_array(26553);
		when "0110011110111010" => data_out <= rom_array(26554);
		when "0110011110111011" => data_out <= rom_array(26555);
		when "0110011110111100" => data_out <= rom_array(26556);
		when "0110011110111101" => data_out <= rom_array(26557);
		when "0110011110111110" => data_out <= rom_array(26558);
		when "0110011110111111" => data_out <= rom_array(26559);
		when "0110011111000000" => data_out <= rom_array(26560);
		when "0110011111000001" => data_out <= rom_array(26561);
		when "0110011111000010" => data_out <= rom_array(26562);
		when "0110011111000011" => data_out <= rom_array(26563);
		when "0110011111000100" => data_out <= rom_array(26564);
		when "0110011111000101" => data_out <= rom_array(26565);
		when "0110011111000110" => data_out <= rom_array(26566);
		when "0110011111000111" => data_out <= rom_array(26567);
		when "0110011111001000" => data_out <= rom_array(26568);
		when "0110011111001001" => data_out <= rom_array(26569);
		when "0110011111001010" => data_out <= rom_array(26570);
		when "0110011111001011" => data_out <= rom_array(26571);
		when "0110011111001100" => data_out <= rom_array(26572);
		when "0110011111001101" => data_out <= rom_array(26573);
		when "0110011111001110" => data_out <= rom_array(26574);
		when "0110011111001111" => data_out <= rom_array(26575);
		when "0110011111010000" => data_out <= rom_array(26576);
		when "0110011111010001" => data_out <= rom_array(26577);
		when "0110011111010010" => data_out <= rom_array(26578);
		when "0110011111010011" => data_out <= rom_array(26579);
		when "0110011111010100" => data_out <= rom_array(26580);
		when "0110011111010101" => data_out <= rom_array(26581);
		when "0110011111010110" => data_out <= rom_array(26582);
		when "0110011111010111" => data_out <= rom_array(26583);
		when "0110011111011000" => data_out <= rom_array(26584);
		when "0110011111011001" => data_out <= rom_array(26585);
		when "0110011111011010" => data_out <= rom_array(26586);
		when "0110011111011011" => data_out <= rom_array(26587);
		when "0110011111011100" => data_out <= rom_array(26588);
		when "0110011111011101" => data_out <= rom_array(26589);
		when "0110011111011110" => data_out <= rom_array(26590);
		when "0110011111011111" => data_out <= rom_array(26591);
		when "0110011111100000" => data_out <= rom_array(26592);
		when "0110011111100001" => data_out <= rom_array(26593);
		when "0110011111100010" => data_out <= rom_array(26594);
		when "0110011111100011" => data_out <= rom_array(26595);
		when "0110011111100100" => data_out <= rom_array(26596);
		when "0110011111100101" => data_out <= rom_array(26597);
		when "0110011111100110" => data_out <= rom_array(26598);
		when "0110011111100111" => data_out <= rom_array(26599);
		when "0110011111101000" => data_out <= rom_array(26600);
		when "0110011111101001" => data_out <= rom_array(26601);
		when "0110011111101010" => data_out <= rom_array(26602);
		when "0110011111101011" => data_out <= rom_array(26603);
		when "0110011111101100" => data_out <= rom_array(26604);
		when "0110011111101101" => data_out <= rom_array(26605);
		when "0110011111101110" => data_out <= rom_array(26606);
		when "0110011111101111" => data_out <= rom_array(26607);
		when "0110011111110000" => data_out <= rom_array(26608);
		when "0110011111110001" => data_out <= rom_array(26609);
		when "0110011111110010" => data_out <= rom_array(26610);
		when "0110011111110011" => data_out <= rom_array(26611);
		when "0110011111110100" => data_out <= rom_array(26612);
		when "0110011111110101" => data_out <= rom_array(26613);
		when "0110011111110110" => data_out <= rom_array(26614);
		when "0110011111110111" => data_out <= rom_array(26615);
		when "0110011111111000" => data_out <= rom_array(26616);
		when "0110011111111001" => data_out <= rom_array(26617);
		when "0110011111111010" => data_out <= rom_array(26618);
		when "0110011111111011" => data_out <= rom_array(26619);
		when "0110011111111100" => data_out <= rom_array(26620);
		when "0110011111111101" => data_out <= rom_array(26621);
		when "0110011111111110" => data_out <= rom_array(26622);
		when "0110011111111111" => data_out <= rom_array(26623);
		when "0110100000000000" => data_out <= rom_array(26624);
		when "0110100000000001" => data_out <= rom_array(26625);
		when "0110100000000010" => data_out <= rom_array(26626);
		when "0110100000000011" => data_out <= rom_array(26627);
		when "0110100000000100" => data_out <= rom_array(26628);
		when "0110100000000101" => data_out <= rom_array(26629);
		when "0110100000000110" => data_out <= rom_array(26630);
		when "0110100000000111" => data_out <= rom_array(26631);
		when "0110100000001000" => data_out <= rom_array(26632);
		when "0110100000001001" => data_out <= rom_array(26633);
		when "0110100000001010" => data_out <= rom_array(26634);
		when "0110100000001011" => data_out <= rom_array(26635);
		when "0110100000001100" => data_out <= rom_array(26636);
		when "0110100000001101" => data_out <= rom_array(26637);
		when "0110100000001110" => data_out <= rom_array(26638);
		when "0110100000001111" => data_out <= rom_array(26639);
		when "0110100000010000" => data_out <= rom_array(26640);
		when "0110100000010001" => data_out <= rom_array(26641);
		when "0110100000010010" => data_out <= rom_array(26642);
		when "0110100000010011" => data_out <= rom_array(26643);
		when "0110100000010100" => data_out <= rom_array(26644);
		when "0110100000010101" => data_out <= rom_array(26645);
		when "0110100000010110" => data_out <= rom_array(26646);
		when "0110100000010111" => data_out <= rom_array(26647);
		when "0110100000011000" => data_out <= rom_array(26648);
		when "0110100000011001" => data_out <= rom_array(26649);
		when "0110100000011010" => data_out <= rom_array(26650);
		when "0110100000011011" => data_out <= rom_array(26651);
		when "0110100000011100" => data_out <= rom_array(26652);
		when "0110100000011101" => data_out <= rom_array(26653);
		when "0110100000011110" => data_out <= rom_array(26654);
		when "0110100000011111" => data_out <= rom_array(26655);
		when "0110100000100000" => data_out <= rom_array(26656);
		when "0110100000100001" => data_out <= rom_array(26657);
		when "0110100000100010" => data_out <= rom_array(26658);
		when "0110100000100011" => data_out <= rom_array(26659);
		when "0110100000100100" => data_out <= rom_array(26660);
		when "0110100000100101" => data_out <= rom_array(26661);
		when "0110100000100110" => data_out <= rom_array(26662);
		when "0110100000100111" => data_out <= rom_array(26663);
		when "0110100000101000" => data_out <= rom_array(26664);
		when "0110100000101001" => data_out <= rom_array(26665);
		when "0110100000101010" => data_out <= rom_array(26666);
		when "0110100000101011" => data_out <= rom_array(26667);
		when "0110100000101100" => data_out <= rom_array(26668);
		when "0110100000101101" => data_out <= rom_array(26669);
		when "0110100000101110" => data_out <= rom_array(26670);
		when "0110100000101111" => data_out <= rom_array(26671);
		when "0110100000110000" => data_out <= rom_array(26672);
		when "0110100000110001" => data_out <= rom_array(26673);
		when "0110100000110010" => data_out <= rom_array(26674);
		when "0110100000110011" => data_out <= rom_array(26675);
		when "0110100000110100" => data_out <= rom_array(26676);
		when "0110100000110101" => data_out <= rom_array(26677);
		when "0110100000110110" => data_out <= rom_array(26678);
		when "0110100000110111" => data_out <= rom_array(26679);
		when "0110100000111000" => data_out <= rom_array(26680);
		when "0110100000111001" => data_out <= rom_array(26681);
		when "0110100000111010" => data_out <= rom_array(26682);
		when "0110100000111011" => data_out <= rom_array(26683);
		when "0110100000111100" => data_out <= rom_array(26684);
		when "0110100000111101" => data_out <= rom_array(26685);
		when "0110100000111110" => data_out <= rom_array(26686);
		when "0110100000111111" => data_out <= rom_array(26687);
		when "0110100001000000" => data_out <= rom_array(26688);
		when "0110100001000001" => data_out <= rom_array(26689);
		when "0110100001000010" => data_out <= rom_array(26690);
		when "0110100001000011" => data_out <= rom_array(26691);
		when "0110100001000100" => data_out <= rom_array(26692);
		when "0110100001000101" => data_out <= rom_array(26693);
		when "0110100001000110" => data_out <= rom_array(26694);
		when "0110100001000111" => data_out <= rom_array(26695);
		when "0110100001001000" => data_out <= rom_array(26696);
		when "0110100001001001" => data_out <= rom_array(26697);
		when "0110100001001010" => data_out <= rom_array(26698);
		when "0110100001001011" => data_out <= rom_array(26699);
		when "0110100001001100" => data_out <= rom_array(26700);
		when "0110100001001101" => data_out <= rom_array(26701);
		when "0110100001001110" => data_out <= rom_array(26702);
		when "0110100001001111" => data_out <= rom_array(26703);
		when "0110100001010000" => data_out <= rom_array(26704);
		when "0110100001010001" => data_out <= rom_array(26705);
		when "0110100001010010" => data_out <= rom_array(26706);
		when "0110100001010011" => data_out <= rom_array(26707);
		when "0110100001010100" => data_out <= rom_array(26708);
		when "0110100001010101" => data_out <= rom_array(26709);
		when "0110100001010110" => data_out <= rom_array(26710);
		when "0110100001010111" => data_out <= rom_array(26711);
		when "0110100001011000" => data_out <= rom_array(26712);
		when "0110100001011001" => data_out <= rom_array(26713);
		when "0110100001011010" => data_out <= rom_array(26714);
		when "0110100001011011" => data_out <= rom_array(26715);
		when "0110100001011100" => data_out <= rom_array(26716);
		when "0110100001011101" => data_out <= rom_array(26717);
		when "0110100001011110" => data_out <= rom_array(26718);
		when "0110100001011111" => data_out <= rom_array(26719);
		when "0110100001100000" => data_out <= rom_array(26720);
		when "0110100001100001" => data_out <= rom_array(26721);
		when "0110100001100010" => data_out <= rom_array(26722);
		when "0110100001100011" => data_out <= rom_array(26723);
		when "0110100001100100" => data_out <= rom_array(26724);
		when "0110100001100101" => data_out <= rom_array(26725);
		when "0110100001100110" => data_out <= rom_array(26726);
		when "0110100001100111" => data_out <= rom_array(26727);
		when "0110100001101000" => data_out <= rom_array(26728);
		when "0110100001101001" => data_out <= rom_array(26729);
		when "0110100001101010" => data_out <= rom_array(26730);
		when "0110100001101011" => data_out <= rom_array(26731);
		when "0110100001101100" => data_out <= rom_array(26732);
		when "0110100001101101" => data_out <= rom_array(26733);
		when "0110100001101110" => data_out <= rom_array(26734);
		when "0110100001101111" => data_out <= rom_array(26735);
		when "0110100001110000" => data_out <= rom_array(26736);
		when "0110100001110001" => data_out <= rom_array(26737);
		when "0110100001110010" => data_out <= rom_array(26738);
		when "0110100001110011" => data_out <= rom_array(26739);
		when "0110100001110100" => data_out <= rom_array(26740);
		when "0110100001110101" => data_out <= rom_array(26741);
		when "0110100001110110" => data_out <= rom_array(26742);
		when "0110100001110111" => data_out <= rom_array(26743);
		when "0110100001111000" => data_out <= rom_array(26744);
		when "0110100001111001" => data_out <= rom_array(26745);
		when "0110100001111010" => data_out <= rom_array(26746);
		when "0110100001111011" => data_out <= rom_array(26747);
		when "0110100001111100" => data_out <= rom_array(26748);
		when "0110100001111101" => data_out <= rom_array(26749);
		when "0110100001111110" => data_out <= rom_array(26750);
		when "0110100001111111" => data_out <= rom_array(26751);
		when "0110100010000000" => data_out <= rom_array(26752);
		when "0110100010000001" => data_out <= rom_array(26753);
		when "0110100010000010" => data_out <= rom_array(26754);
		when "0110100010000011" => data_out <= rom_array(26755);
		when "0110100010000100" => data_out <= rom_array(26756);
		when "0110100010000101" => data_out <= rom_array(26757);
		when "0110100010000110" => data_out <= rom_array(26758);
		when "0110100010000111" => data_out <= rom_array(26759);
		when "0110100010001000" => data_out <= rom_array(26760);
		when "0110100010001001" => data_out <= rom_array(26761);
		when "0110100010001010" => data_out <= rom_array(26762);
		when "0110100010001011" => data_out <= rom_array(26763);
		when "0110100010001100" => data_out <= rom_array(26764);
		when "0110100010001101" => data_out <= rom_array(26765);
		when "0110100010001110" => data_out <= rom_array(26766);
		when "0110100010001111" => data_out <= rom_array(26767);
		when "0110100010010000" => data_out <= rom_array(26768);
		when "0110100010010001" => data_out <= rom_array(26769);
		when "0110100010010010" => data_out <= rom_array(26770);
		when "0110100010010011" => data_out <= rom_array(26771);
		when "0110100010010100" => data_out <= rom_array(26772);
		when "0110100010010101" => data_out <= rom_array(26773);
		when "0110100010010110" => data_out <= rom_array(26774);
		when "0110100010010111" => data_out <= rom_array(26775);
		when "0110100010011000" => data_out <= rom_array(26776);
		when "0110100010011001" => data_out <= rom_array(26777);
		when "0110100010011010" => data_out <= rom_array(26778);
		when "0110100010011011" => data_out <= rom_array(26779);
		when "0110100010011100" => data_out <= rom_array(26780);
		when "0110100010011101" => data_out <= rom_array(26781);
		when "0110100010011110" => data_out <= rom_array(26782);
		when "0110100010011111" => data_out <= rom_array(26783);
		when "0110100010100000" => data_out <= rom_array(26784);
		when "0110100010100001" => data_out <= rom_array(26785);
		when "0110100010100010" => data_out <= rom_array(26786);
		when "0110100010100011" => data_out <= rom_array(26787);
		when "0110100010100100" => data_out <= rom_array(26788);
		when "0110100010100101" => data_out <= rom_array(26789);
		when "0110100010100110" => data_out <= rom_array(26790);
		when "0110100010100111" => data_out <= rom_array(26791);
		when "0110100010101000" => data_out <= rom_array(26792);
		when "0110100010101001" => data_out <= rom_array(26793);
		when "0110100010101010" => data_out <= rom_array(26794);
		when "0110100010101011" => data_out <= rom_array(26795);
		when "0110100010101100" => data_out <= rom_array(26796);
		when "0110100010101101" => data_out <= rom_array(26797);
		when "0110100010101110" => data_out <= rom_array(26798);
		when "0110100010101111" => data_out <= rom_array(26799);
		when "0110100010110000" => data_out <= rom_array(26800);
		when "0110100010110001" => data_out <= rom_array(26801);
		when "0110100010110010" => data_out <= rom_array(26802);
		when "0110100010110011" => data_out <= rom_array(26803);
		when "0110100010110100" => data_out <= rom_array(26804);
		when "0110100010110101" => data_out <= rom_array(26805);
		when "0110100010110110" => data_out <= rom_array(26806);
		when "0110100010110111" => data_out <= rom_array(26807);
		when "0110100010111000" => data_out <= rom_array(26808);
		when "0110100010111001" => data_out <= rom_array(26809);
		when "0110100010111010" => data_out <= rom_array(26810);
		when "0110100010111011" => data_out <= rom_array(26811);
		when "0110100010111100" => data_out <= rom_array(26812);
		when "0110100010111101" => data_out <= rom_array(26813);
		when "0110100010111110" => data_out <= rom_array(26814);
		when "0110100010111111" => data_out <= rom_array(26815);
		when "0110100011000000" => data_out <= rom_array(26816);
		when "0110100011000001" => data_out <= rom_array(26817);
		when "0110100011000010" => data_out <= rom_array(26818);
		when "0110100011000011" => data_out <= rom_array(26819);
		when "0110100011000100" => data_out <= rom_array(26820);
		when "0110100011000101" => data_out <= rom_array(26821);
		when "0110100011000110" => data_out <= rom_array(26822);
		when "0110100011000111" => data_out <= rom_array(26823);
		when "0110100011001000" => data_out <= rom_array(26824);
		when "0110100011001001" => data_out <= rom_array(26825);
		when "0110100011001010" => data_out <= rom_array(26826);
		when "0110100011001011" => data_out <= rom_array(26827);
		when "0110100011001100" => data_out <= rom_array(26828);
		when "0110100011001101" => data_out <= rom_array(26829);
		when "0110100011001110" => data_out <= rom_array(26830);
		when "0110100011001111" => data_out <= rom_array(26831);
		when "0110100011010000" => data_out <= rom_array(26832);
		when "0110100011010001" => data_out <= rom_array(26833);
		when "0110100011010010" => data_out <= rom_array(26834);
		when "0110100011010011" => data_out <= rom_array(26835);
		when "0110100011010100" => data_out <= rom_array(26836);
		when "0110100011010101" => data_out <= rom_array(26837);
		when "0110100011010110" => data_out <= rom_array(26838);
		when "0110100011010111" => data_out <= rom_array(26839);
		when "0110100011011000" => data_out <= rom_array(26840);
		when "0110100011011001" => data_out <= rom_array(26841);
		when "0110100011011010" => data_out <= rom_array(26842);
		when "0110100011011011" => data_out <= rom_array(26843);
		when "0110100011011100" => data_out <= rom_array(26844);
		when "0110100011011101" => data_out <= rom_array(26845);
		when "0110100011011110" => data_out <= rom_array(26846);
		when "0110100011011111" => data_out <= rom_array(26847);
		when "0110100011100000" => data_out <= rom_array(26848);
		when "0110100011100001" => data_out <= rom_array(26849);
		when "0110100011100010" => data_out <= rom_array(26850);
		when "0110100011100011" => data_out <= rom_array(26851);
		when "0110100011100100" => data_out <= rom_array(26852);
		when "0110100011100101" => data_out <= rom_array(26853);
		when "0110100011100110" => data_out <= rom_array(26854);
		when "0110100011100111" => data_out <= rom_array(26855);
		when "0110100011101000" => data_out <= rom_array(26856);
		when "0110100011101001" => data_out <= rom_array(26857);
		when "0110100011101010" => data_out <= rom_array(26858);
		when "0110100011101011" => data_out <= rom_array(26859);
		when "0110100011101100" => data_out <= rom_array(26860);
		when "0110100011101101" => data_out <= rom_array(26861);
		when "0110100011101110" => data_out <= rom_array(26862);
		when "0110100011101111" => data_out <= rom_array(26863);
		when "0110100011110000" => data_out <= rom_array(26864);
		when "0110100011110001" => data_out <= rom_array(26865);
		when "0110100011110010" => data_out <= rom_array(26866);
		when "0110100011110011" => data_out <= rom_array(26867);
		when "0110100011110100" => data_out <= rom_array(26868);
		when "0110100011110101" => data_out <= rom_array(26869);
		when "0110100011110110" => data_out <= rom_array(26870);
		when "0110100011110111" => data_out <= rom_array(26871);
		when "0110100011111000" => data_out <= rom_array(26872);
		when "0110100011111001" => data_out <= rom_array(26873);
		when "0110100011111010" => data_out <= rom_array(26874);
		when "0110100011111011" => data_out <= rom_array(26875);
		when "0110100011111100" => data_out <= rom_array(26876);
		when "0110100011111101" => data_out <= rom_array(26877);
		when "0110100011111110" => data_out <= rom_array(26878);
		when "0110100011111111" => data_out <= rom_array(26879);
		when "0110100100000000" => data_out <= rom_array(26880);
		when "0110100100000001" => data_out <= rom_array(26881);
		when "0110100100000010" => data_out <= rom_array(26882);
		when "0110100100000011" => data_out <= rom_array(26883);
		when "0110100100000100" => data_out <= rom_array(26884);
		when "0110100100000101" => data_out <= rom_array(26885);
		when "0110100100000110" => data_out <= rom_array(26886);
		when "0110100100000111" => data_out <= rom_array(26887);
		when "0110100100001000" => data_out <= rom_array(26888);
		when "0110100100001001" => data_out <= rom_array(26889);
		when "0110100100001010" => data_out <= rom_array(26890);
		when "0110100100001011" => data_out <= rom_array(26891);
		when "0110100100001100" => data_out <= rom_array(26892);
		when "0110100100001101" => data_out <= rom_array(26893);
		when "0110100100001110" => data_out <= rom_array(26894);
		when "0110100100001111" => data_out <= rom_array(26895);
		when "0110100100010000" => data_out <= rom_array(26896);
		when "0110100100010001" => data_out <= rom_array(26897);
		when "0110100100010010" => data_out <= rom_array(26898);
		when "0110100100010011" => data_out <= rom_array(26899);
		when "0110100100010100" => data_out <= rom_array(26900);
		when "0110100100010101" => data_out <= rom_array(26901);
		when "0110100100010110" => data_out <= rom_array(26902);
		when "0110100100010111" => data_out <= rom_array(26903);
		when "0110100100011000" => data_out <= rom_array(26904);
		when "0110100100011001" => data_out <= rom_array(26905);
		when "0110100100011010" => data_out <= rom_array(26906);
		when "0110100100011011" => data_out <= rom_array(26907);
		when "0110100100011100" => data_out <= rom_array(26908);
		when "0110100100011101" => data_out <= rom_array(26909);
		when "0110100100011110" => data_out <= rom_array(26910);
		when "0110100100011111" => data_out <= rom_array(26911);
		when "0110100100100000" => data_out <= rom_array(26912);
		when "0110100100100001" => data_out <= rom_array(26913);
		when "0110100100100010" => data_out <= rom_array(26914);
		when "0110100100100011" => data_out <= rom_array(26915);
		when "0110100100100100" => data_out <= rom_array(26916);
		when "0110100100100101" => data_out <= rom_array(26917);
		when "0110100100100110" => data_out <= rom_array(26918);
		when "0110100100100111" => data_out <= rom_array(26919);
		when "0110100100101000" => data_out <= rom_array(26920);
		when "0110100100101001" => data_out <= rom_array(26921);
		when "0110100100101010" => data_out <= rom_array(26922);
		when "0110100100101011" => data_out <= rom_array(26923);
		when "0110100100101100" => data_out <= rom_array(26924);
		when "0110100100101101" => data_out <= rom_array(26925);
		when "0110100100101110" => data_out <= rom_array(26926);
		when "0110100100101111" => data_out <= rom_array(26927);
		when "0110100100110000" => data_out <= rom_array(26928);
		when "0110100100110001" => data_out <= rom_array(26929);
		when "0110100100110010" => data_out <= rom_array(26930);
		when "0110100100110011" => data_out <= rom_array(26931);
		when "0110100100110100" => data_out <= rom_array(26932);
		when "0110100100110101" => data_out <= rom_array(26933);
		when "0110100100110110" => data_out <= rom_array(26934);
		when "0110100100110111" => data_out <= rom_array(26935);
		when "0110100100111000" => data_out <= rom_array(26936);
		when "0110100100111001" => data_out <= rom_array(26937);
		when "0110100100111010" => data_out <= rom_array(26938);
		when "0110100100111011" => data_out <= rom_array(26939);
		when "0110100100111100" => data_out <= rom_array(26940);
		when "0110100100111101" => data_out <= rom_array(26941);
		when "0110100100111110" => data_out <= rom_array(26942);
		when "0110100100111111" => data_out <= rom_array(26943);
		when "0110100101000000" => data_out <= rom_array(26944);
		when "0110100101000001" => data_out <= rom_array(26945);
		when "0110100101000010" => data_out <= rom_array(26946);
		when "0110100101000011" => data_out <= rom_array(26947);
		when "0110100101000100" => data_out <= rom_array(26948);
		when "0110100101000101" => data_out <= rom_array(26949);
		when "0110100101000110" => data_out <= rom_array(26950);
		when "0110100101000111" => data_out <= rom_array(26951);
		when "0110100101001000" => data_out <= rom_array(26952);
		when "0110100101001001" => data_out <= rom_array(26953);
		when "0110100101001010" => data_out <= rom_array(26954);
		when "0110100101001011" => data_out <= rom_array(26955);
		when "0110100101001100" => data_out <= rom_array(26956);
		when "0110100101001101" => data_out <= rom_array(26957);
		when "0110100101001110" => data_out <= rom_array(26958);
		when "0110100101001111" => data_out <= rom_array(26959);
		when "0110100101010000" => data_out <= rom_array(26960);
		when "0110100101010001" => data_out <= rom_array(26961);
		when "0110100101010010" => data_out <= rom_array(26962);
		when "0110100101010011" => data_out <= rom_array(26963);
		when "0110100101010100" => data_out <= rom_array(26964);
		when "0110100101010101" => data_out <= rom_array(26965);
		when "0110100101010110" => data_out <= rom_array(26966);
		when "0110100101010111" => data_out <= rom_array(26967);
		when "0110100101011000" => data_out <= rom_array(26968);
		when "0110100101011001" => data_out <= rom_array(26969);
		when "0110100101011010" => data_out <= rom_array(26970);
		when "0110100101011011" => data_out <= rom_array(26971);
		when "0110100101011100" => data_out <= rom_array(26972);
		when "0110100101011101" => data_out <= rom_array(26973);
		when "0110100101011110" => data_out <= rom_array(26974);
		when "0110100101011111" => data_out <= rom_array(26975);
		when "0110100101100000" => data_out <= rom_array(26976);
		when "0110100101100001" => data_out <= rom_array(26977);
		when "0110100101100010" => data_out <= rom_array(26978);
		when "0110100101100011" => data_out <= rom_array(26979);
		when "0110100101100100" => data_out <= rom_array(26980);
		when "0110100101100101" => data_out <= rom_array(26981);
		when "0110100101100110" => data_out <= rom_array(26982);
		when "0110100101100111" => data_out <= rom_array(26983);
		when "0110100101101000" => data_out <= rom_array(26984);
		when "0110100101101001" => data_out <= rom_array(26985);
		when "0110100101101010" => data_out <= rom_array(26986);
		when "0110100101101011" => data_out <= rom_array(26987);
		when "0110100101101100" => data_out <= rom_array(26988);
		when "0110100101101101" => data_out <= rom_array(26989);
		when "0110100101101110" => data_out <= rom_array(26990);
		when "0110100101101111" => data_out <= rom_array(26991);
		when "0110100101110000" => data_out <= rom_array(26992);
		when "0110100101110001" => data_out <= rom_array(26993);
		when "0110100101110010" => data_out <= rom_array(26994);
		when "0110100101110011" => data_out <= rom_array(26995);
		when "0110100101110100" => data_out <= rom_array(26996);
		when "0110100101110101" => data_out <= rom_array(26997);
		when "0110100101110110" => data_out <= rom_array(26998);
		when "0110100101110111" => data_out <= rom_array(26999);
		when "0110100101111000" => data_out <= rom_array(27000);
		when "0110100101111001" => data_out <= rom_array(27001);
		when "0110100101111010" => data_out <= rom_array(27002);
		when "0110100101111011" => data_out <= rom_array(27003);
		when "0110100101111100" => data_out <= rom_array(27004);
		when "0110100101111101" => data_out <= rom_array(27005);
		when "0110100101111110" => data_out <= rom_array(27006);
		when "0110100101111111" => data_out <= rom_array(27007);
		when "0110100110000000" => data_out <= rom_array(27008);
		when "0110100110000001" => data_out <= rom_array(27009);
		when "0110100110000010" => data_out <= rom_array(27010);
		when "0110100110000011" => data_out <= rom_array(27011);
		when "0110100110000100" => data_out <= rom_array(27012);
		when "0110100110000101" => data_out <= rom_array(27013);
		when "0110100110000110" => data_out <= rom_array(27014);
		when "0110100110000111" => data_out <= rom_array(27015);
		when "0110100110001000" => data_out <= rom_array(27016);
		when "0110100110001001" => data_out <= rom_array(27017);
		when "0110100110001010" => data_out <= rom_array(27018);
		when "0110100110001011" => data_out <= rom_array(27019);
		when "0110100110001100" => data_out <= rom_array(27020);
		when "0110100110001101" => data_out <= rom_array(27021);
		when "0110100110001110" => data_out <= rom_array(27022);
		when "0110100110001111" => data_out <= rom_array(27023);
		when "0110100110010000" => data_out <= rom_array(27024);
		when "0110100110010001" => data_out <= rom_array(27025);
		when "0110100110010010" => data_out <= rom_array(27026);
		when "0110100110010011" => data_out <= rom_array(27027);
		when "0110100110010100" => data_out <= rom_array(27028);
		when "0110100110010101" => data_out <= rom_array(27029);
		when "0110100110010110" => data_out <= rom_array(27030);
		when "0110100110010111" => data_out <= rom_array(27031);
		when "0110100110011000" => data_out <= rom_array(27032);
		when "0110100110011001" => data_out <= rom_array(27033);
		when "0110100110011010" => data_out <= rom_array(27034);
		when "0110100110011011" => data_out <= rom_array(27035);
		when "0110100110011100" => data_out <= rom_array(27036);
		when "0110100110011101" => data_out <= rom_array(27037);
		when "0110100110011110" => data_out <= rom_array(27038);
		when "0110100110011111" => data_out <= rom_array(27039);
		when "0110100110100000" => data_out <= rom_array(27040);
		when "0110100110100001" => data_out <= rom_array(27041);
		when "0110100110100010" => data_out <= rom_array(27042);
		when "0110100110100011" => data_out <= rom_array(27043);
		when "0110100110100100" => data_out <= rom_array(27044);
		when "0110100110100101" => data_out <= rom_array(27045);
		when "0110100110100110" => data_out <= rom_array(27046);
		when "0110100110100111" => data_out <= rom_array(27047);
		when "0110100110101000" => data_out <= rom_array(27048);
		when "0110100110101001" => data_out <= rom_array(27049);
		when "0110100110101010" => data_out <= rom_array(27050);
		when "0110100110101011" => data_out <= rom_array(27051);
		when "0110100110101100" => data_out <= rom_array(27052);
		when "0110100110101101" => data_out <= rom_array(27053);
		when "0110100110101110" => data_out <= rom_array(27054);
		when "0110100110101111" => data_out <= rom_array(27055);
		when "0110100110110000" => data_out <= rom_array(27056);
		when "0110100110110001" => data_out <= rom_array(27057);
		when "0110100110110010" => data_out <= rom_array(27058);
		when "0110100110110011" => data_out <= rom_array(27059);
		when "0110100110110100" => data_out <= rom_array(27060);
		when "0110100110110101" => data_out <= rom_array(27061);
		when "0110100110110110" => data_out <= rom_array(27062);
		when "0110100110110111" => data_out <= rom_array(27063);
		when "0110100110111000" => data_out <= rom_array(27064);
		when "0110100110111001" => data_out <= rom_array(27065);
		when "0110100110111010" => data_out <= rom_array(27066);
		when "0110100110111011" => data_out <= rom_array(27067);
		when "0110100110111100" => data_out <= rom_array(27068);
		when "0110100110111101" => data_out <= rom_array(27069);
		when "0110100110111110" => data_out <= rom_array(27070);
		when "0110100110111111" => data_out <= rom_array(27071);
		when "0110100111000000" => data_out <= rom_array(27072);
		when "0110100111000001" => data_out <= rom_array(27073);
		when "0110100111000010" => data_out <= rom_array(27074);
		when "0110100111000011" => data_out <= rom_array(27075);
		when "0110100111000100" => data_out <= rom_array(27076);
		when "0110100111000101" => data_out <= rom_array(27077);
		when "0110100111000110" => data_out <= rom_array(27078);
		when "0110100111000111" => data_out <= rom_array(27079);
		when "0110100111001000" => data_out <= rom_array(27080);
		when "0110100111001001" => data_out <= rom_array(27081);
		when "0110100111001010" => data_out <= rom_array(27082);
		when "0110100111001011" => data_out <= rom_array(27083);
		when "0110100111001100" => data_out <= rom_array(27084);
		when "0110100111001101" => data_out <= rom_array(27085);
		when "0110100111001110" => data_out <= rom_array(27086);
		when "0110100111001111" => data_out <= rom_array(27087);
		when "0110100111010000" => data_out <= rom_array(27088);
		when "0110100111010001" => data_out <= rom_array(27089);
		when "0110100111010010" => data_out <= rom_array(27090);
		when "0110100111010011" => data_out <= rom_array(27091);
		when "0110100111010100" => data_out <= rom_array(27092);
		when "0110100111010101" => data_out <= rom_array(27093);
		when "0110100111010110" => data_out <= rom_array(27094);
		when "0110100111010111" => data_out <= rom_array(27095);
		when "0110100111011000" => data_out <= rom_array(27096);
		when "0110100111011001" => data_out <= rom_array(27097);
		when "0110100111011010" => data_out <= rom_array(27098);
		when "0110100111011011" => data_out <= rom_array(27099);
		when "0110100111011100" => data_out <= rom_array(27100);
		when "0110100111011101" => data_out <= rom_array(27101);
		when "0110100111011110" => data_out <= rom_array(27102);
		when "0110100111011111" => data_out <= rom_array(27103);
		when "0110100111100000" => data_out <= rom_array(27104);
		when "0110100111100001" => data_out <= rom_array(27105);
		when "0110100111100010" => data_out <= rom_array(27106);
		when "0110100111100011" => data_out <= rom_array(27107);
		when "0110100111100100" => data_out <= rom_array(27108);
		when "0110100111100101" => data_out <= rom_array(27109);
		when "0110100111100110" => data_out <= rom_array(27110);
		when "0110100111100111" => data_out <= rom_array(27111);
		when "0110100111101000" => data_out <= rom_array(27112);
		when "0110100111101001" => data_out <= rom_array(27113);
		when "0110100111101010" => data_out <= rom_array(27114);
		when "0110100111101011" => data_out <= rom_array(27115);
		when "0110100111101100" => data_out <= rom_array(27116);
		when "0110100111101101" => data_out <= rom_array(27117);
		when "0110100111101110" => data_out <= rom_array(27118);
		when "0110100111101111" => data_out <= rom_array(27119);
		when "0110100111110000" => data_out <= rom_array(27120);
		when "0110100111110001" => data_out <= rom_array(27121);
		when "0110100111110010" => data_out <= rom_array(27122);
		when "0110100111110011" => data_out <= rom_array(27123);
		when "0110100111110100" => data_out <= rom_array(27124);
		when "0110100111110101" => data_out <= rom_array(27125);
		when "0110100111110110" => data_out <= rom_array(27126);
		when "0110100111110111" => data_out <= rom_array(27127);
		when "0110100111111000" => data_out <= rom_array(27128);
		when "0110100111111001" => data_out <= rom_array(27129);
		when "0110100111111010" => data_out <= rom_array(27130);
		when "0110100111111011" => data_out <= rom_array(27131);
		when "0110100111111100" => data_out <= rom_array(27132);
		when "0110100111111101" => data_out <= rom_array(27133);
		when "0110100111111110" => data_out <= rom_array(27134);
		when "0110100111111111" => data_out <= rom_array(27135);
		when "0110101000000000" => data_out <= rom_array(27136);
		when "0110101000000001" => data_out <= rom_array(27137);
		when "0110101000000010" => data_out <= rom_array(27138);
		when "0110101000000011" => data_out <= rom_array(27139);
		when "0110101000000100" => data_out <= rom_array(27140);
		when "0110101000000101" => data_out <= rom_array(27141);
		when "0110101000000110" => data_out <= rom_array(27142);
		when "0110101000000111" => data_out <= rom_array(27143);
		when "0110101000001000" => data_out <= rom_array(27144);
		when "0110101000001001" => data_out <= rom_array(27145);
		when "0110101000001010" => data_out <= rom_array(27146);
		when "0110101000001011" => data_out <= rom_array(27147);
		when "0110101000001100" => data_out <= rom_array(27148);
		when "0110101000001101" => data_out <= rom_array(27149);
		when "0110101000001110" => data_out <= rom_array(27150);
		when "0110101000001111" => data_out <= rom_array(27151);
		when "0110101000010000" => data_out <= rom_array(27152);
		when "0110101000010001" => data_out <= rom_array(27153);
		when "0110101000010010" => data_out <= rom_array(27154);
		when "0110101000010011" => data_out <= rom_array(27155);
		when "0110101000010100" => data_out <= rom_array(27156);
		when "0110101000010101" => data_out <= rom_array(27157);
		when "0110101000010110" => data_out <= rom_array(27158);
		when "0110101000010111" => data_out <= rom_array(27159);
		when "0110101000011000" => data_out <= rom_array(27160);
		when "0110101000011001" => data_out <= rom_array(27161);
		when "0110101000011010" => data_out <= rom_array(27162);
		when "0110101000011011" => data_out <= rom_array(27163);
		when "0110101000011100" => data_out <= rom_array(27164);
		when "0110101000011101" => data_out <= rom_array(27165);
		when "0110101000011110" => data_out <= rom_array(27166);
		when "0110101000011111" => data_out <= rom_array(27167);
		when "0110101000100000" => data_out <= rom_array(27168);
		when "0110101000100001" => data_out <= rom_array(27169);
		when "0110101000100010" => data_out <= rom_array(27170);
		when "0110101000100011" => data_out <= rom_array(27171);
		when "0110101000100100" => data_out <= rom_array(27172);
		when "0110101000100101" => data_out <= rom_array(27173);
		when "0110101000100110" => data_out <= rom_array(27174);
		when "0110101000100111" => data_out <= rom_array(27175);
		when "0110101000101000" => data_out <= rom_array(27176);
		when "0110101000101001" => data_out <= rom_array(27177);
		when "0110101000101010" => data_out <= rom_array(27178);
		when "0110101000101011" => data_out <= rom_array(27179);
		when "0110101000101100" => data_out <= rom_array(27180);
		when "0110101000101101" => data_out <= rom_array(27181);
		when "0110101000101110" => data_out <= rom_array(27182);
		when "0110101000101111" => data_out <= rom_array(27183);
		when "0110101000110000" => data_out <= rom_array(27184);
		when "0110101000110001" => data_out <= rom_array(27185);
		when "0110101000110010" => data_out <= rom_array(27186);
		when "0110101000110011" => data_out <= rom_array(27187);
		when "0110101000110100" => data_out <= rom_array(27188);
		when "0110101000110101" => data_out <= rom_array(27189);
		when "0110101000110110" => data_out <= rom_array(27190);
		when "0110101000110111" => data_out <= rom_array(27191);
		when "0110101000111000" => data_out <= rom_array(27192);
		when "0110101000111001" => data_out <= rom_array(27193);
		when "0110101000111010" => data_out <= rom_array(27194);
		when "0110101000111011" => data_out <= rom_array(27195);
		when "0110101000111100" => data_out <= rom_array(27196);
		when "0110101000111101" => data_out <= rom_array(27197);
		when "0110101000111110" => data_out <= rom_array(27198);
		when "0110101000111111" => data_out <= rom_array(27199);
		when "0110101001000000" => data_out <= rom_array(27200);
		when "0110101001000001" => data_out <= rom_array(27201);
		when "0110101001000010" => data_out <= rom_array(27202);
		when "0110101001000011" => data_out <= rom_array(27203);
		when "0110101001000100" => data_out <= rom_array(27204);
		when "0110101001000101" => data_out <= rom_array(27205);
		when "0110101001000110" => data_out <= rom_array(27206);
		when "0110101001000111" => data_out <= rom_array(27207);
		when "0110101001001000" => data_out <= rom_array(27208);
		when "0110101001001001" => data_out <= rom_array(27209);
		when "0110101001001010" => data_out <= rom_array(27210);
		when "0110101001001011" => data_out <= rom_array(27211);
		when "0110101001001100" => data_out <= rom_array(27212);
		when "0110101001001101" => data_out <= rom_array(27213);
		when "0110101001001110" => data_out <= rom_array(27214);
		when "0110101001001111" => data_out <= rom_array(27215);
		when "0110101001010000" => data_out <= rom_array(27216);
		when "0110101001010001" => data_out <= rom_array(27217);
		when "0110101001010010" => data_out <= rom_array(27218);
		when "0110101001010011" => data_out <= rom_array(27219);
		when "0110101001010100" => data_out <= rom_array(27220);
		when "0110101001010101" => data_out <= rom_array(27221);
		when "0110101001010110" => data_out <= rom_array(27222);
		when "0110101001010111" => data_out <= rom_array(27223);
		when "0110101001011000" => data_out <= rom_array(27224);
		when "0110101001011001" => data_out <= rom_array(27225);
		when "0110101001011010" => data_out <= rom_array(27226);
		when "0110101001011011" => data_out <= rom_array(27227);
		when "0110101001011100" => data_out <= rom_array(27228);
		when "0110101001011101" => data_out <= rom_array(27229);
		when "0110101001011110" => data_out <= rom_array(27230);
		when "0110101001011111" => data_out <= rom_array(27231);
		when "0110101001100000" => data_out <= rom_array(27232);
		when "0110101001100001" => data_out <= rom_array(27233);
		when "0110101001100010" => data_out <= rom_array(27234);
		when "0110101001100011" => data_out <= rom_array(27235);
		when "0110101001100100" => data_out <= rom_array(27236);
		when "0110101001100101" => data_out <= rom_array(27237);
		when "0110101001100110" => data_out <= rom_array(27238);
		when "0110101001100111" => data_out <= rom_array(27239);
		when "0110101001101000" => data_out <= rom_array(27240);
		when "0110101001101001" => data_out <= rom_array(27241);
		when "0110101001101010" => data_out <= rom_array(27242);
		when "0110101001101011" => data_out <= rom_array(27243);
		when "0110101001101100" => data_out <= rom_array(27244);
		when "0110101001101101" => data_out <= rom_array(27245);
		when "0110101001101110" => data_out <= rom_array(27246);
		when "0110101001101111" => data_out <= rom_array(27247);
		when "0110101001110000" => data_out <= rom_array(27248);
		when "0110101001110001" => data_out <= rom_array(27249);
		when "0110101001110010" => data_out <= rom_array(27250);
		when "0110101001110011" => data_out <= rom_array(27251);
		when "0110101001110100" => data_out <= rom_array(27252);
		when "0110101001110101" => data_out <= rom_array(27253);
		when "0110101001110110" => data_out <= rom_array(27254);
		when "0110101001110111" => data_out <= rom_array(27255);
		when "0110101001111000" => data_out <= rom_array(27256);
		when "0110101001111001" => data_out <= rom_array(27257);
		when "0110101001111010" => data_out <= rom_array(27258);
		when "0110101001111011" => data_out <= rom_array(27259);
		when "0110101001111100" => data_out <= rom_array(27260);
		when "0110101001111101" => data_out <= rom_array(27261);
		when "0110101001111110" => data_out <= rom_array(27262);
		when "0110101001111111" => data_out <= rom_array(27263);
		when "0110101010000000" => data_out <= rom_array(27264);
		when "0110101010000001" => data_out <= rom_array(27265);
		when "0110101010000010" => data_out <= rom_array(27266);
		when "0110101010000011" => data_out <= rom_array(27267);
		when "0110101010000100" => data_out <= rom_array(27268);
		when "0110101010000101" => data_out <= rom_array(27269);
		when "0110101010000110" => data_out <= rom_array(27270);
		when "0110101010000111" => data_out <= rom_array(27271);
		when "0110101010001000" => data_out <= rom_array(27272);
		when "0110101010001001" => data_out <= rom_array(27273);
		when "0110101010001010" => data_out <= rom_array(27274);
		when "0110101010001011" => data_out <= rom_array(27275);
		when "0110101010001100" => data_out <= rom_array(27276);
		when "0110101010001101" => data_out <= rom_array(27277);
		when "0110101010001110" => data_out <= rom_array(27278);
		when "0110101010001111" => data_out <= rom_array(27279);
		when "0110101010010000" => data_out <= rom_array(27280);
		when "0110101010010001" => data_out <= rom_array(27281);
		when "0110101010010010" => data_out <= rom_array(27282);
		when "0110101010010011" => data_out <= rom_array(27283);
		when "0110101010010100" => data_out <= rom_array(27284);
		when "0110101010010101" => data_out <= rom_array(27285);
		when "0110101010010110" => data_out <= rom_array(27286);
		when "0110101010010111" => data_out <= rom_array(27287);
		when "0110101010011000" => data_out <= rom_array(27288);
		when "0110101010011001" => data_out <= rom_array(27289);
		when "0110101010011010" => data_out <= rom_array(27290);
		when "0110101010011011" => data_out <= rom_array(27291);
		when "0110101010011100" => data_out <= rom_array(27292);
		when "0110101010011101" => data_out <= rom_array(27293);
		when "0110101010011110" => data_out <= rom_array(27294);
		when "0110101010011111" => data_out <= rom_array(27295);
		when "0110101010100000" => data_out <= rom_array(27296);
		when "0110101010100001" => data_out <= rom_array(27297);
		when "0110101010100010" => data_out <= rom_array(27298);
		when "0110101010100011" => data_out <= rom_array(27299);
		when "0110101010100100" => data_out <= rom_array(27300);
		when "0110101010100101" => data_out <= rom_array(27301);
		when "0110101010100110" => data_out <= rom_array(27302);
		when "0110101010100111" => data_out <= rom_array(27303);
		when "0110101010101000" => data_out <= rom_array(27304);
		when "0110101010101001" => data_out <= rom_array(27305);
		when "0110101010101010" => data_out <= rom_array(27306);
		when "0110101010101011" => data_out <= rom_array(27307);
		when "0110101010101100" => data_out <= rom_array(27308);
		when "0110101010101101" => data_out <= rom_array(27309);
		when "0110101010101110" => data_out <= rom_array(27310);
		when "0110101010101111" => data_out <= rom_array(27311);
		when "0110101010110000" => data_out <= rom_array(27312);
		when "0110101010110001" => data_out <= rom_array(27313);
		when "0110101010110010" => data_out <= rom_array(27314);
		when "0110101010110011" => data_out <= rom_array(27315);
		when "0110101010110100" => data_out <= rom_array(27316);
		when "0110101010110101" => data_out <= rom_array(27317);
		when "0110101010110110" => data_out <= rom_array(27318);
		when "0110101010110111" => data_out <= rom_array(27319);
		when "0110101010111000" => data_out <= rom_array(27320);
		when "0110101010111001" => data_out <= rom_array(27321);
		when "0110101010111010" => data_out <= rom_array(27322);
		when "0110101010111011" => data_out <= rom_array(27323);
		when "0110101010111100" => data_out <= rom_array(27324);
		when "0110101010111101" => data_out <= rom_array(27325);
		when "0110101010111110" => data_out <= rom_array(27326);
		when "0110101010111111" => data_out <= rom_array(27327);
		when "0110101011000000" => data_out <= rom_array(27328);
		when "0110101011000001" => data_out <= rom_array(27329);
		when "0110101011000010" => data_out <= rom_array(27330);
		when "0110101011000011" => data_out <= rom_array(27331);
		when "0110101011000100" => data_out <= rom_array(27332);
		when "0110101011000101" => data_out <= rom_array(27333);
		when "0110101011000110" => data_out <= rom_array(27334);
		when "0110101011000111" => data_out <= rom_array(27335);
		when "0110101011001000" => data_out <= rom_array(27336);
		when "0110101011001001" => data_out <= rom_array(27337);
		when "0110101011001010" => data_out <= rom_array(27338);
		when "0110101011001011" => data_out <= rom_array(27339);
		when "0110101011001100" => data_out <= rom_array(27340);
		when "0110101011001101" => data_out <= rom_array(27341);
		when "0110101011001110" => data_out <= rom_array(27342);
		when "0110101011001111" => data_out <= rom_array(27343);
		when "0110101011010000" => data_out <= rom_array(27344);
		when "0110101011010001" => data_out <= rom_array(27345);
		when "0110101011010010" => data_out <= rom_array(27346);
		when "0110101011010011" => data_out <= rom_array(27347);
		when "0110101011010100" => data_out <= rom_array(27348);
		when "0110101011010101" => data_out <= rom_array(27349);
		when "0110101011010110" => data_out <= rom_array(27350);
		when "0110101011010111" => data_out <= rom_array(27351);
		when "0110101011011000" => data_out <= rom_array(27352);
		when "0110101011011001" => data_out <= rom_array(27353);
		when "0110101011011010" => data_out <= rom_array(27354);
		when "0110101011011011" => data_out <= rom_array(27355);
		when "0110101011011100" => data_out <= rom_array(27356);
		when "0110101011011101" => data_out <= rom_array(27357);
		when "0110101011011110" => data_out <= rom_array(27358);
		when "0110101011011111" => data_out <= rom_array(27359);
		when "0110101011100000" => data_out <= rom_array(27360);
		when "0110101011100001" => data_out <= rom_array(27361);
		when "0110101011100010" => data_out <= rom_array(27362);
		when "0110101011100011" => data_out <= rom_array(27363);
		when "0110101011100100" => data_out <= rom_array(27364);
		when "0110101011100101" => data_out <= rom_array(27365);
		when "0110101011100110" => data_out <= rom_array(27366);
		when "0110101011100111" => data_out <= rom_array(27367);
		when "0110101011101000" => data_out <= rom_array(27368);
		when "0110101011101001" => data_out <= rom_array(27369);
		when "0110101011101010" => data_out <= rom_array(27370);
		when "0110101011101011" => data_out <= rom_array(27371);
		when "0110101011101100" => data_out <= rom_array(27372);
		when "0110101011101101" => data_out <= rom_array(27373);
		when "0110101011101110" => data_out <= rom_array(27374);
		when "0110101011101111" => data_out <= rom_array(27375);
		when "0110101011110000" => data_out <= rom_array(27376);
		when "0110101011110001" => data_out <= rom_array(27377);
		when "0110101011110010" => data_out <= rom_array(27378);
		when "0110101011110011" => data_out <= rom_array(27379);
		when "0110101011110100" => data_out <= rom_array(27380);
		when "0110101011110101" => data_out <= rom_array(27381);
		when "0110101011110110" => data_out <= rom_array(27382);
		when "0110101011110111" => data_out <= rom_array(27383);
		when "0110101011111000" => data_out <= rom_array(27384);
		when "0110101011111001" => data_out <= rom_array(27385);
		when "0110101011111010" => data_out <= rom_array(27386);
		when "0110101011111011" => data_out <= rom_array(27387);
		when "0110101011111100" => data_out <= rom_array(27388);
		when "0110101011111101" => data_out <= rom_array(27389);
		when "0110101011111110" => data_out <= rom_array(27390);
		when "0110101011111111" => data_out <= rom_array(27391);
		when "0110101100000000" => data_out <= rom_array(27392);
		when "0110101100000001" => data_out <= rom_array(27393);
		when "0110101100000010" => data_out <= rom_array(27394);
		when "0110101100000011" => data_out <= rom_array(27395);
		when "0110101100000100" => data_out <= rom_array(27396);
		when "0110101100000101" => data_out <= rom_array(27397);
		when "0110101100000110" => data_out <= rom_array(27398);
		when "0110101100000111" => data_out <= rom_array(27399);
		when "0110101100001000" => data_out <= rom_array(27400);
		when "0110101100001001" => data_out <= rom_array(27401);
		when "0110101100001010" => data_out <= rom_array(27402);
		when "0110101100001011" => data_out <= rom_array(27403);
		when "0110101100001100" => data_out <= rom_array(27404);
		when "0110101100001101" => data_out <= rom_array(27405);
		when "0110101100001110" => data_out <= rom_array(27406);
		when "0110101100001111" => data_out <= rom_array(27407);
		when "0110101100010000" => data_out <= rom_array(27408);
		when "0110101100010001" => data_out <= rom_array(27409);
		when "0110101100010010" => data_out <= rom_array(27410);
		when "0110101100010011" => data_out <= rom_array(27411);
		when "0110101100010100" => data_out <= rom_array(27412);
		when "0110101100010101" => data_out <= rom_array(27413);
		when "0110101100010110" => data_out <= rom_array(27414);
		when "0110101100010111" => data_out <= rom_array(27415);
		when "0110101100011000" => data_out <= rom_array(27416);
		when "0110101100011001" => data_out <= rom_array(27417);
		when "0110101100011010" => data_out <= rom_array(27418);
		when "0110101100011011" => data_out <= rom_array(27419);
		when "0110101100011100" => data_out <= rom_array(27420);
		when "0110101100011101" => data_out <= rom_array(27421);
		when "0110101100011110" => data_out <= rom_array(27422);
		when "0110101100011111" => data_out <= rom_array(27423);
		when "0110101100100000" => data_out <= rom_array(27424);
		when "0110101100100001" => data_out <= rom_array(27425);
		when "0110101100100010" => data_out <= rom_array(27426);
		when "0110101100100011" => data_out <= rom_array(27427);
		when "0110101100100100" => data_out <= rom_array(27428);
		when "0110101100100101" => data_out <= rom_array(27429);
		when "0110101100100110" => data_out <= rom_array(27430);
		when "0110101100100111" => data_out <= rom_array(27431);
		when "0110101100101000" => data_out <= rom_array(27432);
		when "0110101100101001" => data_out <= rom_array(27433);
		when "0110101100101010" => data_out <= rom_array(27434);
		when "0110101100101011" => data_out <= rom_array(27435);
		when "0110101100101100" => data_out <= rom_array(27436);
		when "0110101100101101" => data_out <= rom_array(27437);
		when "0110101100101110" => data_out <= rom_array(27438);
		when "0110101100101111" => data_out <= rom_array(27439);
		when "0110101100110000" => data_out <= rom_array(27440);
		when "0110101100110001" => data_out <= rom_array(27441);
		when "0110101100110010" => data_out <= rom_array(27442);
		when "0110101100110011" => data_out <= rom_array(27443);
		when "0110101100110100" => data_out <= rom_array(27444);
		when "0110101100110101" => data_out <= rom_array(27445);
		when "0110101100110110" => data_out <= rom_array(27446);
		when "0110101100110111" => data_out <= rom_array(27447);
		when "0110101100111000" => data_out <= rom_array(27448);
		when "0110101100111001" => data_out <= rom_array(27449);
		when "0110101100111010" => data_out <= rom_array(27450);
		when "0110101100111011" => data_out <= rom_array(27451);
		when "0110101100111100" => data_out <= rom_array(27452);
		when "0110101100111101" => data_out <= rom_array(27453);
		when "0110101100111110" => data_out <= rom_array(27454);
		when "0110101100111111" => data_out <= rom_array(27455);
		when "0110101101000000" => data_out <= rom_array(27456);
		when "0110101101000001" => data_out <= rom_array(27457);
		when "0110101101000010" => data_out <= rom_array(27458);
		when "0110101101000011" => data_out <= rom_array(27459);
		when "0110101101000100" => data_out <= rom_array(27460);
		when "0110101101000101" => data_out <= rom_array(27461);
		when "0110101101000110" => data_out <= rom_array(27462);
		when "0110101101000111" => data_out <= rom_array(27463);
		when "0110101101001000" => data_out <= rom_array(27464);
		when "0110101101001001" => data_out <= rom_array(27465);
		when "0110101101001010" => data_out <= rom_array(27466);
		when "0110101101001011" => data_out <= rom_array(27467);
		when "0110101101001100" => data_out <= rom_array(27468);
		when "0110101101001101" => data_out <= rom_array(27469);
		when "0110101101001110" => data_out <= rom_array(27470);
		when "0110101101001111" => data_out <= rom_array(27471);
		when "0110101101010000" => data_out <= rom_array(27472);
		when "0110101101010001" => data_out <= rom_array(27473);
		when "0110101101010010" => data_out <= rom_array(27474);
		when "0110101101010011" => data_out <= rom_array(27475);
		when "0110101101010100" => data_out <= rom_array(27476);
		when "0110101101010101" => data_out <= rom_array(27477);
		when "0110101101010110" => data_out <= rom_array(27478);
		when "0110101101010111" => data_out <= rom_array(27479);
		when "0110101101011000" => data_out <= rom_array(27480);
		when "0110101101011001" => data_out <= rom_array(27481);
		when "0110101101011010" => data_out <= rom_array(27482);
		when "0110101101011011" => data_out <= rom_array(27483);
		when "0110101101011100" => data_out <= rom_array(27484);
		when "0110101101011101" => data_out <= rom_array(27485);
		when "0110101101011110" => data_out <= rom_array(27486);
		when "0110101101011111" => data_out <= rom_array(27487);
		when "0110101101100000" => data_out <= rom_array(27488);
		when "0110101101100001" => data_out <= rom_array(27489);
		when "0110101101100010" => data_out <= rom_array(27490);
		when "0110101101100011" => data_out <= rom_array(27491);
		when "0110101101100100" => data_out <= rom_array(27492);
		when "0110101101100101" => data_out <= rom_array(27493);
		when "0110101101100110" => data_out <= rom_array(27494);
		when "0110101101100111" => data_out <= rom_array(27495);
		when "0110101101101000" => data_out <= rom_array(27496);
		when "0110101101101001" => data_out <= rom_array(27497);
		when "0110101101101010" => data_out <= rom_array(27498);
		when "0110101101101011" => data_out <= rom_array(27499);
		when "0110101101101100" => data_out <= rom_array(27500);
		when "0110101101101101" => data_out <= rom_array(27501);
		when "0110101101101110" => data_out <= rom_array(27502);
		when "0110101101101111" => data_out <= rom_array(27503);
		when "0110101101110000" => data_out <= rom_array(27504);
		when "0110101101110001" => data_out <= rom_array(27505);
		when "0110101101110010" => data_out <= rom_array(27506);
		when "0110101101110011" => data_out <= rom_array(27507);
		when "0110101101110100" => data_out <= rom_array(27508);
		when "0110101101110101" => data_out <= rom_array(27509);
		when "0110101101110110" => data_out <= rom_array(27510);
		when "0110101101110111" => data_out <= rom_array(27511);
		when "0110101101111000" => data_out <= rom_array(27512);
		when "0110101101111001" => data_out <= rom_array(27513);
		when "0110101101111010" => data_out <= rom_array(27514);
		when "0110101101111011" => data_out <= rom_array(27515);
		when "0110101101111100" => data_out <= rom_array(27516);
		when "0110101101111101" => data_out <= rom_array(27517);
		when "0110101101111110" => data_out <= rom_array(27518);
		when "0110101101111111" => data_out <= rom_array(27519);
		when "0110101110000000" => data_out <= rom_array(27520);
		when "0110101110000001" => data_out <= rom_array(27521);
		when "0110101110000010" => data_out <= rom_array(27522);
		when "0110101110000011" => data_out <= rom_array(27523);
		when "0110101110000100" => data_out <= rom_array(27524);
		when "0110101110000101" => data_out <= rom_array(27525);
		when "0110101110000110" => data_out <= rom_array(27526);
		when "0110101110000111" => data_out <= rom_array(27527);
		when "0110101110001000" => data_out <= rom_array(27528);
		when "0110101110001001" => data_out <= rom_array(27529);
		when "0110101110001010" => data_out <= rom_array(27530);
		when "0110101110001011" => data_out <= rom_array(27531);
		when "0110101110001100" => data_out <= rom_array(27532);
		when "0110101110001101" => data_out <= rom_array(27533);
		when "0110101110001110" => data_out <= rom_array(27534);
		when "0110101110001111" => data_out <= rom_array(27535);
		when "0110101110010000" => data_out <= rom_array(27536);
		when "0110101110010001" => data_out <= rom_array(27537);
		when "0110101110010010" => data_out <= rom_array(27538);
		when "0110101110010011" => data_out <= rom_array(27539);
		when "0110101110010100" => data_out <= rom_array(27540);
		when "0110101110010101" => data_out <= rom_array(27541);
		when "0110101110010110" => data_out <= rom_array(27542);
		when "0110101110010111" => data_out <= rom_array(27543);
		when "0110101110011000" => data_out <= rom_array(27544);
		when "0110101110011001" => data_out <= rom_array(27545);
		when "0110101110011010" => data_out <= rom_array(27546);
		when "0110101110011011" => data_out <= rom_array(27547);
		when "0110101110011100" => data_out <= rom_array(27548);
		when "0110101110011101" => data_out <= rom_array(27549);
		when "0110101110011110" => data_out <= rom_array(27550);
		when "0110101110011111" => data_out <= rom_array(27551);
		when "0110101110100000" => data_out <= rom_array(27552);
		when "0110101110100001" => data_out <= rom_array(27553);
		when "0110101110100010" => data_out <= rom_array(27554);
		when "0110101110100011" => data_out <= rom_array(27555);
		when "0110101110100100" => data_out <= rom_array(27556);
		when "0110101110100101" => data_out <= rom_array(27557);
		when "0110101110100110" => data_out <= rom_array(27558);
		when "0110101110100111" => data_out <= rom_array(27559);
		when "0110101110101000" => data_out <= rom_array(27560);
		when "0110101110101001" => data_out <= rom_array(27561);
		when "0110101110101010" => data_out <= rom_array(27562);
		when "0110101110101011" => data_out <= rom_array(27563);
		when "0110101110101100" => data_out <= rom_array(27564);
		when "0110101110101101" => data_out <= rom_array(27565);
		when "0110101110101110" => data_out <= rom_array(27566);
		when "0110101110101111" => data_out <= rom_array(27567);
		when "0110101110110000" => data_out <= rom_array(27568);
		when "0110101110110001" => data_out <= rom_array(27569);
		when "0110101110110010" => data_out <= rom_array(27570);
		when "0110101110110011" => data_out <= rom_array(27571);
		when "0110101110110100" => data_out <= rom_array(27572);
		when "0110101110110101" => data_out <= rom_array(27573);
		when "0110101110110110" => data_out <= rom_array(27574);
		when "0110101110110111" => data_out <= rom_array(27575);
		when "0110101110111000" => data_out <= rom_array(27576);
		when "0110101110111001" => data_out <= rom_array(27577);
		when "0110101110111010" => data_out <= rom_array(27578);
		when "0110101110111011" => data_out <= rom_array(27579);
		when "0110101110111100" => data_out <= rom_array(27580);
		when "0110101110111101" => data_out <= rom_array(27581);
		when "0110101110111110" => data_out <= rom_array(27582);
		when "0110101110111111" => data_out <= rom_array(27583);
		when "0110101111000000" => data_out <= rom_array(27584);
		when "0110101111000001" => data_out <= rom_array(27585);
		when "0110101111000010" => data_out <= rom_array(27586);
		when "0110101111000011" => data_out <= rom_array(27587);
		when "0110101111000100" => data_out <= rom_array(27588);
		when "0110101111000101" => data_out <= rom_array(27589);
		when "0110101111000110" => data_out <= rom_array(27590);
		when "0110101111000111" => data_out <= rom_array(27591);
		when "0110101111001000" => data_out <= rom_array(27592);
		when "0110101111001001" => data_out <= rom_array(27593);
		when "0110101111001010" => data_out <= rom_array(27594);
		when "0110101111001011" => data_out <= rom_array(27595);
		when "0110101111001100" => data_out <= rom_array(27596);
		when "0110101111001101" => data_out <= rom_array(27597);
		when "0110101111001110" => data_out <= rom_array(27598);
		when "0110101111001111" => data_out <= rom_array(27599);
		when "0110101111010000" => data_out <= rom_array(27600);
		when "0110101111010001" => data_out <= rom_array(27601);
		when "0110101111010010" => data_out <= rom_array(27602);
		when "0110101111010011" => data_out <= rom_array(27603);
		when "0110101111010100" => data_out <= rom_array(27604);
		when "0110101111010101" => data_out <= rom_array(27605);
		when "0110101111010110" => data_out <= rom_array(27606);
		when "0110101111010111" => data_out <= rom_array(27607);
		when "0110101111011000" => data_out <= rom_array(27608);
		when "0110101111011001" => data_out <= rom_array(27609);
		when "0110101111011010" => data_out <= rom_array(27610);
		when "0110101111011011" => data_out <= rom_array(27611);
		when "0110101111011100" => data_out <= rom_array(27612);
		when "0110101111011101" => data_out <= rom_array(27613);
		when "0110101111011110" => data_out <= rom_array(27614);
		when "0110101111011111" => data_out <= rom_array(27615);
		when "0110101111100000" => data_out <= rom_array(27616);
		when "0110101111100001" => data_out <= rom_array(27617);
		when "0110101111100010" => data_out <= rom_array(27618);
		when "0110101111100011" => data_out <= rom_array(27619);
		when "0110101111100100" => data_out <= rom_array(27620);
		when "0110101111100101" => data_out <= rom_array(27621);
		when "0110101111100110" => data_out <= rom_array(27622);
		when "0110101111100111" => data_out <= rom_array(27623);
		when "0110101111101000" => data_out <= rom_array(27624);
		when "0110101111101001" => data_out <= rom_array(27625);
		when "0110101111101010" => data_out <= rom_array(27626);
		when "0110101111101011" => data_out <= rom_array(27627);
		when "0110101111101100" => data_out <= rom_array(27628);
		when "0110101111101101" => data_out <= rom_array(27629);
		when "0110101111101110" => data_out <= rom_array(27630);
		when "0110101111101111" => data_out <= rom_array(27631);
		when "0110101111110000" => data_out <= rom_array(27632);
		when "0110101111110001" => data_out <= rom_array(27633);
		when "0110101111110010" => data_out <= rom_array(27634);
		when "0110101111110011" => data_out <= rom_array(27635);
		when "0110101111110100" => data_out <= rom_array(27636);
		when "0110101111110101" => data_out <= rom_array(27637);
		when "0110101111110110" => data_out <= rom_array(27638);
		when "0110101111110111" => data_out <= rom_array(27639);
		when "0110101111111000" => data_out <= rom_array(27640);
		when "0110101111111001" => data_out <= rom_array(27641);
		when "0110101111111010" => data_out <= rom_array(27642);
		when "0110101111111011" => data_out <= rom_array(27643);
		when "0110101111111100" => data_out <= rom_array(27644);
		when "0110101111111101" => data_out <= rom_array(27645);
		when "0110101111111110" => data_out <= rom_array(27646);
		when "0110101111111111" => data_out <= rom_array(27647);
		when "0110110000000000" => data_out <= rom_array(27648);
		when "0110110000000001" => data_out <= rom_array(27649);
		when "0110110000000010" => data_out <= rom_array(27650);
		when "0110110000000011" => data_out <= rom_array(27651);
		when "0110110000000100" => data_out <= rom_array(27652);
		when "0110110000000101" => data_out <= rom_array(27653);
		when "0110110000000110" => data_out <= rom_array(27654);
		when "0110110000000111" => data_out <= rom_array(27655);
		when "0110110000001000" => data_out <= rom_array(27656);
		when "0110110000001001" => data_out <= rom_array(27657);
		when "0110110000001010" => data_out <= rom_array(27658);
		when "0110110000001011" => data_out <= rom_array(27659);
		when "0110110000001100" => data_out <= rom_array(27660);
		when "0110110000001101" => data_out <= rom_array(27661);
		when "0110110000001110" => data_out <= rom_array(27662);
		when "0110110000001111" => data_out <= rom_array(27663);
		when "0110110000010000" => data_out <= rom_array(27664);
		when "0110110000010001" => data_out <= rom_array(27665);
		when "0110110000010010" => data_out <= rom_array(27666);
		when "0110110000010011" => data_out <= rom_array(27667);
		when "0110110000010100" => data_out <= rom_array(27668);
		when "0110110000010101" => data_out <= rom_array(27669);
		when "0110110000010110" => data_out <= rom_array(27670);
		when "0110110000010111" => data_out <= rom_array(27671);
		when "0110110000011000" => data_out <= rom_array(27672);
		when "0110110000011001" => data_out <= rom_array(27673);
		when "0110110000011010" => data_out <= rom_array(27674);
		when "0110110000011011" => data_out <= rom_array(27675);
		when "0110110000011100" => data_out <= rom_array(27676);
		when "0110110000011101" => data_out <= rom_array(27677);
		when "0110110000011110" => data_out <= rom_array(27678);
		when "0110110000011111" => data_out <= rom_array(27679);
		when "0110110000100000" => data_out <= rom_array(27680);
		when "0110110000100001" => data_out <= rom_array(27681);
		when "0110110000100010" => data_out <= rom_array(27682);
		when "0110110000100011" => data_out <= rom_array(27683);
		when "0110110000100100" => data_out <= rom_array(27684);
		when "0110110000100101" => data_out <= rom_array(27685);
		when "0110110000100110" => data_out <= rom_array(27686);
		when "0110110000100111" => data_out <= rom_array(27687);
		when "0110110000101000" => data_out <= rom_array(27688);
		when "0110110000101001" => data_out <= rom_array(27689);
		when "0110110000101010" => data_out <= rom_array(27690);
		when "0110110000101011" => data_out <= rom_array(27691);
		when "0110110000101100" => data_out <= rom_array(27692);
		when "0110110000101101" => data_out <= rom_array(27693);
		when "0110110000101110" => data_out <= rom_array(27694);
		when "0110110000101111" => data_out <= rom_array(27695);
		when "0110110000110000" => data_out <= rom_array(27696);
		when "0110110000110001" => data_out <= rom_array(27697);
		when "0110110000110010" => data_out <= rom_array(27698);
		when "0110110000110011" => data_out <= rom_array(27699);
		when "0110110000110100" => data_out <= rom_array(27700);
		when "0110110000110101" => data_out <= rom_array(27701);
		when "0110110000110110" => data_out <= rom_array(27702);
		when "0110110000110111" => data_out <= rom_array(27703);
		when "0110110000111000" => data_out <= rom_array(27704);
		when "0110110000111001" => data_out <= rom_array(27705);
		when "0110110000111010" => data_out <= rom_array(27706);
		when "0110110000111011" => data_out <= rom_array(27707);
		when "0110110000111100" => data_out <= rom_array(27708);
		when "0110110000111101" => data_out <= rom_array(27709);
		when "0110110000111110" => data_out <= rom_array(27710);
		when "0110110000111111" => data_out <= rom_array(27711);
		when "0110110001000000" => data_out <= rom_array(27712);
		when "0110110001000001" => data_out <= rom_array(27713);
		when "0110110001000010" => data_out <= rom_array(27714);
		when "0110110001000011" => data_out <= rom_array(27715);
		when "0110110001000100" => data_out <= rom_array(27716);
		when "0110110001000101" => data_out <= rom_array(27717);
		when "0110110001000110" => data_out <= rom_array(27718);
		when "0110110001000111" => data_out <= rom_array(27719);
		when "0110110001001000" => data_out <= rom_array(27720);
		when "0110110001001001" => data_out <= rom_array(27721);
		when "0110110001001010" => data_out <= rom_array(27722);
		when "0110110001001011" => data_out <= rom_array(27723);
		when "0110110001001100" => data_out <= rom_array(27724);
		when "0110110001001101" => data_out <= rom_array(27725);
		when "0110110001001110" => data_out <= rom_array(27726);
		when "0110110001001111" => data_out <= rom_array(27727);
		when "0110110001010000" => data_out <= rom_array(27728);
		when "0110110001010001" => data_out <= rom_array(27729);
		when "0110110001010010" => data_out <= rom_array(27730);
		when "0110110001010011" => data_out <= rom_array(27731);
		when "0110110001010100" => data_out <= rom_array(27732);
		when "0110110001010101" => data_out <= rom_array(27733);
		when "0110110001010110" => data_out <= rom_array(27734);
		when "0110110001010111" => data_out <= rom_array(27735);
		when "0110110001011000" => data_out <= rom_array(27736);
		when "0110110001011001" => data_out <= rom_array(27737);
		when "0110110001011010" => data_out <= rom_array(27738);
		when "0110110001011011" => data_out <= rom_array(27739);
		when "0110110001011100" => data_out <= rom_array(27740);
		when "0110110001011101" => data_out <= rom_array(27741);
		when "0110110001011110" => data_out <= rom_array(27742);
		when "0110110001011111" => data_out <= rom_array(27743);
		when "0110110001100000" => data_out <= rom_array(27744);
		when "0110110001100001" => data_out <= rom_array(27745);
		when "0110110001100010" => data_out <= rom_array(27746);
		when "0110110001100011" => data_out <= rom_array(27747);
		when "0110110001100100" => data_out <= rom_array(27748);
		when "0110110001100101" => data_out <= rom_array(27749);
		when "0110110001100110" => data_out <= rom_array(27750);
		when "0110110001100111" => data_out <= rom_array(27751);
		when "0110110001101000" => data_out <= rom_array(27752);
		when "0110110001101001" => data_out <= rom_array(27753);
		when "0110110001101010" => data_out <= rom_array(27754);
		when "0110110001101011" => data_out <= rom_array(27755);
		when "0110110001101100" => data_out <= rom_array(27756);
		when "0110110001101101" => data_out <= rom_array(27757);
		when "0110110001101110" => data_out <= rom_array(27758);
		when "0110110001101111" => data_out <= rom_array(27759);
		when "0110110001110000" => data_out <= rom_array(27760);
		when "0110110001110001" => data_out <= rom_array(27761);
		when "0110110001110010" => data_out <= rom_array(27762);
		when "0110110001110011" => data_out <= rom_array(27763);
		when "0110110001110100" => data_out <= rom_array(27764);
		when "0110110001110101" => data_out <= rom_array(27765);
		when "0110110001110110" => data_out <= rom_array(27766);
		when "0110110001110111" => data_out <= rom_array(27767);
		when "0110110001111000" => data_out <= rom_array(27768);
		when "0110110001111001" => data_out <= rom_array(27769);
		when "0110110001111010" => data_out <= rom_array(27770);
		when "0110110001111011" => data_out <= rom_array(27771);
		when "0110110001111100" => data_out <= rom_array(27772);
		when "0110110001111101" => data_out <= rom_array(27773);
		when "0110110001111110" => data_out <= rom_array(27774);
		when "0110110001111111" => data_out <= rom_array(27775);
		when "0110110010000000" => data_out <= rom_array(27776);
		when "0110110010000001" => data_out <= rom_array(27777);
		when "0110110010000010" => data_out <= rom_array(27778);
		when "0110110010000011" => data_out <= rom_array(27779);
		when "0110110010000100" => data_out <= rom_array(27780);
		when "0110110010000101" => data_out <= rom_array(27781);
		when "0110110010000110" => data_out <= rom_array(27782);
		when "0110110010000111" => data_out <= rom_array(27783);
		when "0110110010001000" => data_out <= rom_array(27784);
		when "0110110010001001" => data_out <= rom_array(27785);
		when "0110110010001010" => data_out <= rom_array(27786);
		when "0110110010001011" => data_out <= rom_array(27787);
		when "0110110010001100" => data_out <= rom_array(27788);
		when "0110110010001101" => data_out <= rom_array(27789);
		when "0110110010001110" => data_out <= rom_array(27790);
		when "0110110010001111" => data_out <= rom_array(27791);
		when "0110110010010000" => data_out <= rom_array(27792);
		when "0110110010010001" => data_out <= rom_array(27793);
		when "0110110010010010" => data_out <= rom_array(27794);
		when "0110110010010011" => data_out <= rom_array(27795);
		when "0110110010010100" => data_out <= rom_array(27796);
		when "0110110010010101" => data_out <= rom_array(27797);
		when "0110110010010110" => data_out <= rom_array(27798);
		when "0110110010010111" => data_out <= rom_array(27799);
		when "0110110010011000" => data_out <= rom_array(27800);
		when "0110110010011001" => data_out <= rom_array(27801);
		when "0110110010011010" => data_out <= rom_array(27802);
		when "0110110010011011" => data_out <= rom_array(27803);
		when "0110110010011100" => data_out <= rom_array(27804);
		when "0110110010011101" => data_out <= rom_array(27805);
		when "0110110010011110" => data_out <= rom_array(27806);
		when "0110110010011111" => data_out <= rom_array(27807);
		when "0110110010100000" => data_out <= rom_array(27808);
		when "0110110010100001" => data_out <= rom_array(27809);
		when "0110110010100010" => data_out <= rom_array(27810);
		when "0110110010100011" => data_out <= rom_array(27811);
		when "0110110010100100" => data_out <= rom_array(27812);
		when "0110110010100101" => data_out <= rom_array(27813);
		when "0110110010100110" => data_out <= rom_array(27814);
		when "0110110010100111" => data_out <= rom_array(27815);
		when "0110110010101000" => data_out <= rom_array(27816);
		when "0110110010101001" => data_out <= rom_array(27817);
		when "0110110010101010" => data_out <= rom_array(27818);
		when "0110110010101011" => data_out <= rom_array(27819);
		when "0110110010101100" => data_out <= rom_array(27820);
		when "0110110010101101" => data_out <= rom_array(27821);
		when "0110110010101110" => data_out <= rom_array(27822);
		when "0110110010101111" => data_out <= rom_array(27823);
		when "0110110010110000" => data_out <= rom_array(27824);
		when "0110110010110001" => data_out <= rom_array(27825);
		when "0110110010110010" => data_out <= rom_array(27826);
		when "0110110010110011" => data_out <= rom_array(27827);
		when "0110110010110100" => data_out <= rom_array(27828);
		when "0110110010110101" => data_out <= rom_array(27829);
		when "0110110010110110" => data_out <= rom_array(27830);
		when "0110110010110111" => data_out <= rom_array(27831);
		when "0110110010111000" => data_out <= rom_array(27832);
		when "0110110010111001" => data_out <= rom_array(27833);
		when "0110110010111010" => data_out <= rom_array(27834);
		when "0110110010111011" => data_out <= rom_array(27835);
		when "0110110010111100" => data_out <= rom_array(27836);
		when "0110110010111101" => data_out <= rom_array(27837);
		when "0110110010111110" => data_out <= rom_array(27838);
		when "0110110010111111" => data_out <= rom_array(27839);
		when "0110110011000000" => data_out <= rom_array(27840);
		when "0110110011000001" => data_out <= rom_array(27841);
		when "0110110011000010" => data_out <= rom_array(27842);
		when "0110110011000011" => data_out <= rom_array(27843);
		when "0110110011000100" => data_out <= rom_array(27844);
		when "0110110011000101" => data_out <= rom_array(27845);
		when "0110110011000110" => data_out <= rom_array(27846);
		when "0110110011000111" => data_out <= rom_array(27847);
		when "0110110011001000" => data_out <= rom_array(27848);
		when "0110110011001001" => data_out <= rom_array(27849);
		when "0110110011001010" => data_out <= rom_array(27850);
		when "0110110011001011" => data_out <= rom_array(27851);
		when "0110110011001100" => data_out <= rom_array(27852);
		when "0110110011001101" => data_out <= rom_array(27853);
		when "0110110011001110" => data_out <= rom_array(27854);
		when "0110110011001111" => data_out <= rom_array(27855);
		when "0110110011010000" => data_out <= rom_array(27856);
		when "0110110011010001" => data_out <= rom_array(27857);
		when "0110110011010010" => data_out <= rom_array(27858);
		when "0110110011010011" => data_out <= rom_array(27859);
		when "0110110011010100" => data_out <= rom_array(27860);
		when "0110110011010101" => data_out <= rom_array(27861);
		when "0110110011010110" => data_out <= rom_array(27862);
		when "0110110011010111" => data_out <= rom_array(27863);
		when "0110110011011000" => data_out <= rom_array(27864);
		when "0110110011011001" => data_out <= rom_array(27865);
		when "0110110011011010" => data_out <= rom_array(27866);
		when "0110110011011011" => data_out <= rom_array(27867);
		when "0110110011011100" => data_out <= rom_array(27868);
		when "0110110011011101" => data_out <= rom_array(27869);
		when "0110110011011110" => data_out <= rom_array(27870);
		when "0110110011011111" => data_out <= rom_array(27871);
		when "0110110011100000" => data_out <= rom_array(27872);
		when "0110110011100001" => data_out <= rom_array(27873);
		when "0110110011100010" => data_out <= rom_array(27874);
		when "0110110011100011" => data_out <= rom_array(27875);
		when "0110110011100100" => data_out <= rom_array(27876);
		when "0110110011100101" => data_out <= rom_array(27877);
		when "0110110011100110" => data_out <= rom_array(27878);
		when "0110110011100111" => data_out <= rom_array(27879);
		when "0110110011101000" => data_out <= rom_array(27880);
		when "0110110011101001" => data_out <= rom_array(27881);
		when "0110110011101010" => data_out <= rom_array(27882);
		when "0110110011101011" => data_out <= rom_array(27883);
		when "0110110011101100" => data_out <= rom_array(27884);
		when "0110110011101101" => data_out <= rom_array(27885);
		when "0110110011101110" => data_out <= rom_array(27886);
		when "0110110011101111" => data_out <= rom_array(27887);
		when "0110110011110000" => data_out <= rom_array(27888);
		when "0110110011110001" => data_out <= rom_array(27889);
		when "0110110011110010" => data_out <= rom_array(27890);
		when "0110110011110011" => data_out <= rom_array(27891);
		when "0110110011110100" => data_out <= rom_array(27892);
		when "0110110011110101" => data_out <= rom_array(27893);
		when "0110110011110110" => data_out <= rom_array(27894);
		when "0110110011110111" => data_out <= rom_array(27895);
		when "0110110011111000" => data_out <= rom_array(27896);
		when "0110110011111001" => data_out <= rom_array(27897);
		when "0110110011111010" => data_out <= rom_array(27898);
		when "0110110011111011" => data_out <= rom_array(27899);
		when "0110110011111100" => data_out <= rom_array(27900);
		when "0110110011111101" => data_out <= rom_array(27901);
		when "0110110011111110" => data_out <= rom_array(27902);
		when "0110110011111111" => data_out <= rom_array(27903);
		when "0110110100000000" => data_out <= rom_array(27904);
		when "0110110100000001" => data_out <= rom_array(27905);
		when "0110110100000010" => data_out <= rom_array(27906);
		when "0110110100000011" => data_out <= rom_array(27907);
		when "0110110100000100" => data_out <= rom_array(27908);
		when "0110110100000101" => data_out <= rom_array(27909);
		when "0110110100000110" => data_out <= rom_array(27910);
		when "0110110100000111" => data_out <= rom_array(27911);
		when "0110110100001000" => data_out <= rom_array(27912);
		when "0110110100001001" => data_out <= rom_array(27913);
		when "0110110100001010" => data_out <= rom_array(27914);
		when "0110110100001011" => data_out <= rom_array(27915);
		when "0110110100001100" => data_out <= rom_array(27916);
		when "0110110100001101" => data_out <= rom_array(27917);
		when "0110110100001110" => data_out <= rom_array(27918);
		when "0110110100001111" => data_out <= rom_array(27919);
		when "0110110100010000" => data_out <= rom_array(27920);
		when "0110110100010001" => data_out <= rom_array(27921);
		when "0110110100010010" => data_out <= rom_array(27922);
		when "0110110100010011" => data_out <= rom_array(27923);
		when "0110110100010100" => data_out <= rom_array(27924);
		when "0110110100010101" => data_out <= rom_array(27925);
		when "0110110100010110" => data_out <= rom_array(27926);
		when "0110110100010111" => data_out <= rom_array(27927);
		when "0110110100011000" => data_out <= rom_array(27928);
		when "0110110100011001" => data_out <= rom_array(27929);
		when "0110110100011010" => data_out <= rom_array(27930);
		when "0110110100011011" => data_out <= rom_array(27931);
		when "0110110100011100" => data_out <= rom_array(27932);
		when "0110110100011101" => data_out <= rom_array(27933);
		when "0110110100011110" => data_out <= rom_array(27934);
		when "0110110100011111" => data_out <= rom_array(27935);
		when "0110110100100000" => data_out <= rom_array(27936);
		when "0110110100100001" => data_out <= rom_array(27937);
		when "0110110100100010" => data_out <= rom_array(27938);
		when "0110110100100011" => data_out <= rom_array(27939);
		when "0110110100100100" => data_out <= rom_array(27940);
		when "0110110100100101" => data_out <= rom_array(27941);
		when "0110110100100110" => data_out <= rom_array(27942);
		when "0110110100100111" => data_out <= rom_array(27943);
		when "0110110100101000" => data_out <= rom_array(27944);
		when "0110110100101001" => data_out <= rom_array(27945);
		when "0110110100101010" => data_out <= rom_array(27946);
		when "0110110100101011" => data_out <= rom_array(27947);
		when "0110110100101100" => data_out <= rom_array(27948);
		when "0110110100101101" => data_out <= rom_array(27949);
		when "0110110100101110" => data_out <= rom_array(27950);
		when "0110110100101111" => data_out <= rom_array(27951);
		when "0110110100110000" => data_out <= rom_array(27952);
		when "0110110100110001" => data_out <= rom_array(27953);
		when "0110110100110010" => data_out <= rom_array(27954);
		when "0110110100110011" => data_out <= rom_array(27955);
		when "0110110100110100" => data_out <= rom_array(27956);
		when "0110110100110101" => data_out <= rom_array(27957);
		when "0110110100110110" => data_out <= rom_array(27958);
		when "0110110100110111" => data_out <= rom_array(27959);
		when "0110110100111000" => data_out <= rom_array(27960);
		when "0110110100111001" => data_out <= rom_array(27961);
		when "0110110100111010" => data_out <= rom_array(27962);
		when "0110110100111011" => data_out <= rom_array(27963);
		when "0110110100111100" => data_out <= rom_array(27964);
		when "0110110100111101" => data_out <= rom_array(27965);
		when "0110110100111110" => data_out <= rom_array(27966);
		when "0110110100111111" => data_out <= rom_array(27967);
		when "0110110101000000" => data_out <= rom_array(27968);
		when "0110110101000001" => data_out <= rom_array(27969);
		when "0110110101000010" => data_out <= rom_array(27970);
		when "0110110101000011" => data_out <= rom_array(27971);
		when "0110110101000100" => data_out <= rom_array(27972);
		when "0110110101000101" => data_out <= rom_array(27973);
		when "0110110101000110" => data_out <= rom_array(27974);
		when "0110110101000111" => data_out <= rom_array(27975);
		when "0110110101001000" => data_out <= rom_array(27976);
		when "0110110101001001" => data_out <= rom_array(27977);
		when "0110110101001010" => data_out <= rom_array(27978);
		when "0110110101001011" => data_out <= rom_array(27979);
		when "0110110101001100" => data_out <= rom_array(27980);
		when "0110110101001101" => data_out <= rom_array(27981);
		when "0110110101001110" => data_out <= rom_array(27982);
		when "0110110101001111" => data_out <= rom_array(27983);
		when "0110110101010000" => data_out <= rom_array(27984);
		when "0110110101010001" => data_out <= rom_array(27985);
		when "0110110101010010" => data_out <= rom_array(27986);
		when "0110110101010011" => data_out <= rom_array(27987);
		when "0110110101010100" => data_out <= rom_array(27988);
		when "0110110101010101" => data_out <= rom_array(27989);
		when "0110110101010110" => data_out <= rom_array(27990);
		when "0110110101010111" => data_out <= rom_array(27991);
		when "0110110101011000" => data_out <= rom_array(27992);
		when "0110110101011001" => data_out <= rom_array(27993);
		when "0110110101011010" => data_out <= rom_array(27994);
		when "0110110101011011" => data_out <= rom_array(27995);
		when "0110110101011100" => data_out <= rom_array(27996);
		when "0110110101011101" => data_out <= rom_array(27997);
		when "0110110101011110" => data_out <= rom_array(27998);
		when "0110110101011111" => data_out <= rom_array(27999);
		when "0110110101100000" => data_out <= rom_array(28000);
		when "0110110101100001" => data_out <= rom_array(28001);
		when "0110110101100010" => data_out <= rom_array(28002);
		when "0110110101100011" => data_out <= rom_array(28003);
		when "0110110101100100" => data_out <= rom_array(28004);
		when "0110110101100101" => data_out <= rom_array(28005);
		when "0110110101100110" => data_out <= rom_array(28006);
		when "0110110101100111" => data_out <= rom_array(28007);
		when "0110110101101000" => data_out <= rom_array(28008);
		when "0110110101101001" => data_out <= rom_array(28009);
		when "0110110101101010" => data_out <= rom_array(28010);
		when "0110110101101011" => data_out <= rom_array(28011);
		when "0110110101101100" => data_out <= rom_array(28012);
		when "0110110101101101" => data_out <= rom_array(28013);
		when "0110110101101110" => data_out <= rom_array(28014);
		when "0110110101101111" => data_out <= rom_array(28015);
		when "0110110101110000" => data_out <= rom_array(28016);
		when "0110110101110001" => data_out <= rom_array(28017);
		when "0110110101110010" => data_out <= rom_array(28018);
		when "0110110101110011" => data_out <= rom_array(28019);
		when "0110110101110100" => data_out <= rom_array(28020);
		when "0110110101110101" => data_out <= rom_array(28021);
		when "0110110101110110" => data_out <= rom_array(28022);
		when "0110110101110111" => data_out <= rom_array(28023);
		when "0110110101111000" => data_out <= rom_array(28024);
		when "0110110101111001" => data_out <= rom_array(28025);
		when "0110110101111010" => data_out <= rom_array(28026);
		when "0110110101111011" => data_out <= rom_array(28027);
		when "0110110101111100" => data_out <= rom_array(28028);
		when "0110110101111101" => data_out <= rom_array(28029);
		when "0110110101111110" => data_out <= rom_array(28030);
		when "0110110101111111" => data_out <= rom_array(28031);
		when "0110110110000000" => data_out <= rom_array(28032);
		when "0110110110000001" => data_out <= rom_array(28033);
		when "0110110110000010" => data_out <= rom_array(28034);
		when "0110110110000011" => data_out <= rom_array(28035);
		when "0110110110000100" => data_out <= rom_array(28036);
		when "0110110110000101" => data_out <= rom_array(28037);
		when "0110110110000110" => data_out <= rom_array(28038);
		when "0110110110000111" => data_out <= rom_array(28039);
		when "0110110110001000" => data_out <= rom_array(28040);
		when "0110110110001001" => data_out <= rom_array(28041);
		when "0110110110001010" => data_out <= rom_array(28042);
		when "0110110110001011" => data_out <= rom_array(28043);
		when "0110110110001100" => data_out <= rom_array(28044);
		when "0110110110001101" => data_out <= rom_array(28045);
		when "0110110110001110" => data_out <= rom_array(28046);
		when "0110110110001111" => data_out <= rom_array(28047);
		when "0110110110010000" => data_out <= rom_array(28048);
		when "0110110110010001" => data_out <= rom_array(28049);
		when "0110110110010010" => data_out <= rom_array(28050);
		when "0110110110010011" => data_out <= rom_array(28051);
		when "0110110110010100" => data_out <= rom_array(28052);
		when "0110110110010101" => data_out <= rom_array(28053);
		when "0110110110010110" => data_out <= rom_array(28054);
		when "0110110110010111" => data_out <= rom_array(28055);
		when "0110110110011000" => data_out <= rom_array(28056);
		when "0110110110011001" => data_out <= rom_array(28057);
		when "0110110110011010" => data_out <= rom_array(28058);
		when "0110110110011011" => data_out <= rom_array(28059);
		when "0110110110011100" => data_out <= rom_array(28060);
		when "0110110110011101" => data_out <= rom_array(28061);
		when "0110110110011110" => data_out <= rom_array(28062);
		when "0110110110011111" => data_out <= rom_array(28063);
		when "0110110110100000" => data_out <= rom_array(28064);
		when "0110110110100001" => data_out <= rom_array(28065);
		when "0110110110100010" => data_out <= rom_array(28066);
		when "0110110110100011" => data_out <= rom_array(28067);
		when "0110110110100100" => data_out <= rom_array(28068);
		when "0110110110100101" => data_out <= rom_array(28069);
		when "0110110110100110" => data_out <= rom_array(28070);
		when "0110110110100111" => data_out <= rom_array(28071);
		when "0110110110101000" => data_out <= rom_array(28072);
		when "0110110110101001" => data_out <= rom_array(28073);
		when "0110110110101010" => data_out <= rom_array(28074);
		when "0110110110101011" => data_out <= rom_array(28075);
		when "0110110110101100" => data_out <= rom_array(28076);
		when "0110110110101101" => data_out <= rom_array(28077);
		when "0110110110101110" => data_out <= rom_array(28078);
		when "0110110110101111" => data_out <= rom_array(28079);
		when "0110110110110000" => data_out <= rom_array(28080);
		when "0110110110110001" => data_out <= rom_array(28081);
		when "0110110110110010" => data_out <= rom_array(28082);
		when "0110110110110011" => data_out <= rom_array(28083);
		when "0110110110110100" => data_out <= rom_array(28084);
		when "0110110110110101" => data_out <= rom_array(28085);
		when "0110110110110110" => data_out <= rom_array(28086);
		when "0110110110110111" => data_out <= rom_array(28087);
		when "0110110110111000" => data_out <= rom_array(28088);
		when "0110110110111001" => data_out <= rom_array(28089);
		when "0110110110111010" => data_out <= rom_array(28090);
		when "0110110110111011" => data_out <= rom_array(28091);
		when "0110110110111100" => data_out <= rom_array(28092);
		when "0110110110111101" => data_out <= rom_array(28093);
		when "0110110110111110" => data_out <= rom_array(28094);
		when "0110110110111111" => data_out <= rom_array(28095);
		when "0110110111000000" => data_out <= rom_array(28096);
		when "0110110111000001" => data_out <= rom_array(28097);
		when "0110110111000010" => data_out <= rom_array(28098);
		when "0110110111000011" => data_out <= rom_array(28099);
		when "0110110111000100" => data_out <= rom_array(28100);
		when "0110110111000101" => data_out <= rom_array(28101);
		when "0110110111000110" => data_out <= rom_array(28102);
		when "0110110111000111" => data_out <= rom_array(28103);
		when "0110110111001000" => data_out <= rom_array(28104);
		when "0110110111001001" => data_out <= rom_array(28105);
		when "0110110111001010" => data_out <= rom_array(28106);
		when "0110110111001011" => data_out <= rom_array(28107);
		when "0110110111001100" => data_out <= rom_array(28108);
		when "0110110111001101" => data_out <= rom_array(28109);
		when "0110110111001110" => data_out <= rom_array(28110);
		when "0110110111001111" => data_out <= rom_array(28111);
		when "0110110111010000" => data_out <= rom_array(28112);
		when "0110110111010001" => data_out <= rom_array(28113);
		when "0110110111010010" => data_out <= rom_array(28114);
		when "0110110111010011" => data_out <= rom_array(28115);
		when "0110110111010100" => data_out <= rom_array(28116);
		when "0110110111010101" => data_out <= rom_array(28117);
		when "0110110111010110" => data_out <= rom_array(28118);
		when "0110110111010111" => data_out <= rom_array(28119);
		when "0110110111011000" => data_out <= rom_array(28120);
		when "0110110111011001" => data_out <= rom_array(28121);
		when "0110110111011010" => data_out <= rom_array(28122);
		when "0110110111011011" => data_out <= rom_array(28123);
		when "0110110111011100" => data_out <= rom_array(28124);
		when "0110110111011101" => data_out <= rom_array(28125);
		when "0110110111011110" => data_out <= rom_array(28126);
		when "0110110111011111" => data_out <= rom_array(28127);
		when "0110110111100000" => data_out <= rom_array(28128);
		when "0110110111100001" => data_out <= rom_array(28129);
		when "0110110111100010" => data_out <= rom_array(28130);
		when "0110110111100011" => data_out <= rom_array(28131);
		when "0110110111100100" => data_out <= rom_array(28132);
		when "0110110111100101" => data_out <= rom_array(28133);
		when "0110110111100110" => data_out <= rom_array(28134);
		when "0110110111100111" => data_out <= rom_array(28135);
		when "0110110111101000" => data_out <= rom_array(28136);
		when "0110110111101001" => data_out <= rom_array(28137);
		when "0110110111101010" => data_out <= rom_array(28138);
		when "0110110111101011" => data_out <= rom_array(28139);
		when "0110110111101100" => data_out <= rom_array(28140);
		when "0110110111101101" => data_out <= rom_array(28141);
		when "0110110111101110" => data_out <= rom_array(28142);
		when "0110110111101111" => data_out <= rom_array(28143);
		when "0110110111110000" => data_out <= rom_array(28144);
		when "0110110111110001" => data_out <= rom_array(28145);
		when "0110110111110010" => data_out <= rom_array(28146);
		when "0110110111110011" => data_out <= rom_array(28147);
		when "0110110111110100" => data_out <= rom_array(28148);
		when "0110110111110101" => data_out <= rom_array(28149);
		when "0110110111110110" => data_out <= rom_array(28150);
		when "0110110111110111" => data_out <= rom_array(28151);
		when "0110110111111000" => data_out <= rom_array(28152);
		when "0110110111111001" => data_out <= rom_array(28153);
		when "0110110111111010" => data_out <= rom_array(28154);
		when "0110110111111011" => data_out <= rom_array(28155);
		when "0110110111111100" => data_out <= rom_array(28156);
		when "0110110111111101" => data_out <= rom_array(28157);
		when "0110110111111110" => data_out <= rom_array(28158);
		when "0110110111111111" => data_out <= rom_array(28159);
		when "0110111000000000" => data_out <= rom_array(28160);
		when "0110111000000001" => data_out <= rom_array(28161);
		when "0110111000000010" => data_out <= rom_array(28162);
		when "0110111000000011" => data_out <= rom_array(28163);
		when "0110111000000100" => data_out <= rom_array(28164);
		when "0110111000000101" => data_out <= rom_array(28165);
		when "0110111000000110" => data_out <= rom_array(28166);
		when "0110111000000111" => data_out <= rom_array(28167);
		when "0110111000001000" => data_out <= rom_array(28168);
		when "0110111000001001" => data_out <= rom_array(28169);
		when "0110111000001010" => data_out <= rom_array(28170);
		when "0110111000001011" => data_out <= rom_array(28171);
		when "0110111000001100" => data_out <= rom_array(28172);
		when "0110111000001101" => data_out <= rom_array(28173);
		when "0110111000001110" => data_out <= rom_array(28174);
		when "0110111000001111" => data_out <= rom_array(28175);
		when "0110111000010000" => data_out <= rom_array(28176);
		when "0110111000010001" => data_out <= rom_array(28177);
		when "0110111000010010" => data_out <= rom_array(28178);
		when "0110111000010011" => data_out <= rom_array(28179);
		when "0110111000010100" => data_out <= rom_array(28180);
		when "0110111000010101" => data_out <= rom_array(28181);
		when "0110111000010110" => data_out <= rom_array(28182);
		when "0110111000010111" => data_out <= rom_array(28183);
		when "0110111000011000" => data_out <= rom_array(28184);
		when "0110111000011001" => data_out <= rom_array(28185);
		when "0110111000011010" => data_out <= rom_array(28186);
		when "0110111000011011" => data_out <= rom_array(28187);
		when "0110111000011100" => data_out <= rom_array(28188);
		when "0110111000011101" => data_out <= rom_array(28189);
		when "0110111000011110" => data_out <= rom_array(28190);
		when "0110111000011111" => data_out <= rom_array(28191);
		when "0110111000100000" => data_out <= rom_array(28192);
		when "0110111000100001" => data_out <= rom_array(28193);
		when "0110111000100010" => data_out <= rom_array(28194);
		when "0110111000100011" => data_out <= rom_array(28195);
		when "0110111000100100" => data_out <= rom_array(28196);
		when "0110111000100101" => data_out <= rom_array(28197);
		when "0110111000100110" => data_out <= rom_array(28198);
		when "0110111000100111" => data_out <= rom_array(28199);
		when "0110111000101000" => data_out <= rom_array(28200);
		when "0110111000101001" => data_out <= rom_array(28201);
		when "0110111000101010" => data_out <= rom_array(28202);
		when "0110111000101011" => data_out <= rom_array(28203);
		when "0110111000101100" => data_out <= rom_array(28204);
		when "0110111000101101" => data_out <= rom_array(28205);
		when "0110111000101110" => data_out <= rom_array(28206);
		when "0110111000101111" => data_out <= rom_array(28207);
		when "0110111000110000" => data_out <= rom_array(28208);
		when "0110111000110001" => data_out <= rom_array(28209);
		when "0110111000110010" => data_out <= rom_array(28210);
		when "0110111000110011" => data_out <= rom_array(28211);
		when "0110111000110100" => data_out <= rom_array(28212);
		when "0110111000110101" => data_out <= rom_array(28213);
		when "0110111000110110" => data_out <= rom_array(28214);
		when "0110111000110111" => data_out <= rom_array(28215);
		when "0110111000111000" => data_out <= rom_array(28216);
		when "0110111000111001" => data_out <= rom_array(28217);
		when "0110111000111010" => data_out <= rom_array(28218);
		when "0110111000111011" => data_out <= rom_array(28219);
		when "0110111000111100" => data_out <= rom_array(28220);
		when "0110111000111101" => data_out <= rom_array(28221);
		when "0110111000111110" => data_out <= rom_array(28222);
		when "0110111000111111" => data_out <= rom_array(28223);
		when "0110111001000000" => data_out <= rom_array(28224);
		when "0110111001000001" => data_out <= rom_array(28225);
		when "0110111001000010" => data_out <= rom_array(28226);
		when "0110111001000011" => data_out <= rom_array(28227);
		when "0110111001000100" => data_out <= rom_array(28228);
		when "0110111001000101" => data_out <= rom_array(28229);
		when "0110111001000110" => data_out <= rom_array(28230);
		when "0110111001000111" => data_out <= rom_array(28231);
		when "0110111001001000" => data_out <= rom_array(28232);
		when "0110111001001001" => data_out <= rom_array(28233);
		when "0110111001001010" => data_out <= rom_array(28234);
		when "0110111001001011" => data_out <= rom_array(28235);
		when "0110111001001100" => data_out <= rom_array(28236);
		when "0110111001001101" => data_out <= rom_array(28237);
		when "0110111001001110" => data_out <= rom_array(28238);
		when "0110111001001111" => data_out <= rom_array(28239);
		when "0110111001010000" => data_out <= rom_array(28240);
		when "0110111001010001" => data_out <= rom_array(28241);
		when "0110111001010010" => data_out <= rom_array(28242);
		when "0110111001010011" => data_out <= rom_array(28243);
		when "0110111001010100" => data_out <= rom_array(28244);
		when "0110111001010101" => data_out <= rom_array(28245);
		when "0110111001010110" => data_out <= rom_array(28246);
		when "0110111001010111" => data_out <= rom_array(28247);
		when "0110111001011000" => data_out <= rom_array(28248);
		when "0110111001011001" => data_out <= rom_array(28249);
		when "0110111001011010" => data_out <= rom_array(28250);
		when "0110111001011011" => data_out <= rom_array(28251);
		when "0110111001011100" => data_out <= rom_array(28252);
		when "0110111001011101" => data_out <= rom_array(28253);
		when "0110111001011110" => data_out <= rom_array(28254);
		when "0110111001011111" => data_out <= rom_array(28255);
		when "0110111001100000" => data_out <= rom_array(28256);
		when "0110111001100001" => data_out <= rom_array(28257);
		when "0110111001100010" => data_out <= rom_array(28258);
		when "0110111001100011" => data_out <= rom_array(28259);
		when "0110111001100100" => data_out <= rom_array(28260);
		when "0110111001100101" => data_out <= rom_array(28261);
		when "0110111001100110" => data_out <= rom_array(28262);
		when "0110111001100111" => data_out <= rom_array(28263);
		when "0110111001101000" => data_out <= rom_array(28264);
		when "0110111001101001" => data_out <= rom_array(28265);
		when "0110111001101010" => data_out <= rom_array(28266);
		when "0110111001101011" => data_out <= rom_array(28267);
		when "0110111001101100" => data_out <= rom_array(28268);
		when "0110111001101101" => data_out <= rom_array(28269);
		when "0110111001101110" => data_out <= rom_array(28270);
		when "0110111001101111" => data_out <= rom_array(28271);
		when "0110111001110000" => data_out <= rom_array(28272);
		when "0110111001110001" => data_out <= rom_array(28273);
		when "0110111001110010" => data_out <= rom_array(28274);
		when "0110111001110011" => data_out <= rom_array(28275);
		when "0110111001110100" => data_out <= rom_array(28276);
		when "0110111001110101" => data_out <= rom_array(28277);
		when "0110111001110110" => data_out <= rom_array(28278);
		when "0110111001110111" => data_out <= rom_array(28279);
		when "0110111001111000" => data_out <= rom_array(28280);
		when "0110111001111001" => data_out <= rom_array(28281);
		when "0110111001111010" => data_out <= rom_array(28282);
		when "0110111001111011" => data_out <= rom_array(28283);
		when "0110111001111100" => data_out <= rom_array(28284);
		when "0110111001111101" => data_out <= rom_array(28285);
		when "0110111001111110" => data_out <= rom_array(28286);
		when "0110111001111111" => data_out <= rom_array(28287);
		when "0110111010000000" => data_out <= rom_array(28288);
		when "0110111010000001" => data_out <= rom_array(28289);
		when "0110111010000010" => data_out <= rom_array(28290);
		when "0110111010000011" => data_out <= rom_array(28291);
		when "0110111010000100" => data_out <= rom_array(28292);
		when "0110111010000101" => data_out <= rom_array(28293);
		when "0110111010000110" => data_out <= rom_array(28294);
		when "0110111010000111" => data_out <= rom_array(28295);
		when "0110111010001000" => data_out <= rom_array(28296);
		when "0110111010001001" => data_out <= rom_array(28297);
		when "0110111010001010" => data_out <= rom_array(28298);
		when "0110111010001011" => data_out <= rom_array(28299);
		when "0110111010001100" => data_out <= rom_array(28300);
		when "0110111010001101" => data_out <= rom_array(28301);
		when "0110111010001110" => data_out <= rom_array(28302);
		when "0110111010001111" => data_out <= rom_array(28303);
		when "0110111010010000" => data_out <= rom_array(28304);
		when "0110111010010001" => data_out <= rom_array(28305);
		when "0110111010010010" => data_out <= rom_array(28306);
		when "0110111010010011" => data_out <= rom_array(28307);
		when "0110111010010100" => data_out <= rom_array(28308);
		when "0110111010010101" => data_out <= rom_array(28309);
		when "0110111010010110" => data_out <= rom_array(28310);
		when "0110111010010111" => data_out <= rom_array(28311);
		when "0110111010011000" => data_out <= rom_array(28312);
		when "0110111010011001" => data_out <= rom_array(28313);
		when "0110111010011010" => data_out <= rom_array(28314);
		when "0110111010011011" => data_out <= rom_array(28315);
		when "0110111010011100" => data_out <= rom_array(28316);
		when "0110111010011101" => data_out <= rom_array(28317);
		when "0110111010011110" => data_out <= rom_array(28318);
		when "0110111010011111" => data_out <= rom_array(28319);
		when "0110111010100000" => data_out <= rom_array(28320);
		when "0110111010100001" => data_out <= rom_array(28321);
		when "0110111010100010" => data_out <= rom_array(28322);
		when "0110111010100011" => data_out <= rom_array(28323);
		when "0110111010100100" => data_out <= rom_array(28324);
		when "0110111010100101" => data_out <= rom_array(28325);
		when "0110111010100110" => data_out <= rom_array(28326);
		when "0110111010100111" => data_out <= rom_array(28327);
		when "0110111010101000" => data_out <= rom_array(28328);
		when "0110111010101001" => data_out <= rom_array(28329);
		when "0110111010101010" => data_out <= rom_array(28330);
		when "0110111010101011" => data_out <= rom_array(28331);
		when "0110111010101100" => data_out <= rom_array(28332);
		when "0110111010101101" => data_out <= rom_array(28333);
		when "0110111010101110" => data_out <= rom_array(28334);
		when "0110111010101111" => data_out <= rom_array(28335);
		when "0110111010110000" => data_out <= rom_array(28336);
		when "0110111010110001" => data_out <= rom_array(28337);
		when "0110111010110010" => data_out <= rom_array(28338);
		when "0110111010110011" => data_out <= rom_array(28339);
		when "0110111010110100" => data_out <= rom_array(28340);
		when "0110111010110101" => data_out <= rom_array(28341);
		when "0110111010110110" => data_out <= rom_array(28342);
		when "0110111010110111" => data_out <= rom_array(28343);
		when "0110111010111000" => data_out <= rom_array(28344);
		when "0110111010111001" => data_out <= rom_array(28345);
		when "0110111010111010" => data_out <= rom_array(28346);
		when "0110111010111011" => data_out <= rom_array(28347);
		when "0110111010111100" => data_out <= rom_array(28348);
		when "0110111010111101" => data_out <= rom_array(28349);
		when "0110111010111110" => data_out <= rom_array(28350);
		when "0110111010111111" => data_out <= rom_array(28351);
		when "0110111011000000" => data_out <= rom_array(28352);
		when "0110111011000001" => data_out <= rom_array(28353);
		when "0110111011000010" => data_out <= rom_array(28354);
		when "0110111011000011" => data_out <= rom_array(28355);
		when "0110111011000100" => data_out <= rom_array(28356);
		when "0110111011000101" => data_out <= rom_array(28357);
		when "0110111011000110" => data_out <= rom_array(28358);
		when "0110111011000111" => data_out <= rom_array(28359);
		when "0110111011001000" => data_out <= rom_array(28360);
		when "0110111011001001" => data_out <= rom_array(28361);
		when "0110111011001010" => data_out <= rom_array(28362);
		when "0110111011001011" => data_out <= rom_array(28363);
		when "0110111011001100" => data_out <= rom_array(28364);
		when "0110111011001101" => data_out <= rom_array(28365);
		when "0110111011001110" => data_out <= rom_array(28366);
		when "0110111011001111" => data_out <= rom_array(28367);
		when "0110111011010000" => data_out <= rom_array(28368);
		when "0110111011010001" => data_out <= rom_array(28369);
		when "0110111011010010" => data_out <= rom_array(28370);
		when "0110111011010011" => data_out <= rom_array(28371);
		when "0110111011010100" => data_out <= rom_array(28372);
		when "0110111011010101" => data_out <= rom_array(28373);
		when "0110111011010110" => data_out <= rom_array(28374);
		when "0110111011010111" => data_out <= rom_array(28375);
		when "0110111011011000" => data_out <= rom_array(28376);
		when "0110111011011001" => data_out <= rom_array(28377);
		when "0110111011011010" => data_out <= rom_array(28378);
		when "0110111011011011" => data_out <= rom_array(28379);
		when "0110111011011100" => data_out <= rom_array(28380);
		when "0110111011011101" => data_out <= rom_array(28381);
		when "0110111011011110" => data_out <= rom_array(28382);
		when "0110111011011111" => data_out <= rom_array(28383);
		when "0110111011100000" => data_out <= rom_array(28384);
		when "0110111011100001" => data_out <= rom_array(28385);
		when "0110111011100010" => data_out <= rom_array(28386);
		when "0110111011100011" => data_out <= rom_array(28387);
		when "0110111011100100" => data_out <= rom_array(28388);
		when "0110111011100101" => data_out <= rom_array(28389);
		when "0110111011100110" => data_out <= rom_array(28390);
		when "0110111011100111" => data_out <= rom_array(28391);
		when "0110111011101000" => data_out <= rom_array(28392);
		when "0110111011101001" => data_out <= rom_array(28393);
		when "0110111011101010" => data_out <= rom_array(28394);
		when "0110111011101011" => data_out <= rom_array(28395);
		when "0110111011101100" => data_out <= rom_array(28396);
		when "0110111011101101" => data_out <= rom_array(28397);
		when "0110111011101110" => data_out <= rom_array(28398);
		when "0110111011101111" => data_out <= rom_array(28399);
		when "0110111011110000" => data_out <= rom_array(28400);
		when "0110111011110001" => data_out <= rom_array(28401);
		when "0110111011110010" => data_out <= rom_array(28402);
		when "0110111011110011" => data_out <= rom_array(28403);
		when "0110111011110100" => data_out <= rom_array(28404);
		when "0110111011110101" => data_out <= rom_array(28405);
		when "0110111011110110" => data_out <= rom_array(28406);
		when "0110111011110111" => data_out <= rom_array(28407);
		when "0110111011111000" => data_out <= rom_array(28408);
		when "0110111011111001" => data_out <= rom_array(28409);
		when "0110111011111010" => data_out <= rom_array(28410);
		when "0110111011111011" => data_out <= rom_array(28411);
		when "0110111011111100" => data_out <= rom_array(28412);
		when "0110111011111101" => data_out <= rom_array(28413);
		when "0110111011111110" => data_out <= rom_array(28414);
		when "0110111011111111" => data_out <= rom_array(28415);
		when "0110111100000000" => data_out <= rom_array(28416);
		when "0110111100000001" => data_out <= rom_array(28417);
		when "0110111100000010" => data_out <= rom_array(28418);
		when "0110111100000011" => data_out <= rom_array(28419);
		when "0110111100000100" => data_out <= rom_array(28420);
		when "0110111100000101" => data_out <= rom_array(28421);
		when "0110111100000110" => data_out <= rom_array(28422);
		when "0110111100000111" => data_out <= rom_array(28423);
		when "0110111100001000" => data_out <= rom_array(28424);
		when "0110111100001001" => data_out <= rom_array(28425);
		when "0110111100001010" => data_out <= rom_array(28426);
		when "0110111100001011" => data_out <= rom_array(28427);
		when "0110111100001100" => data_out <= rom_array(28428);
		when "0110111100001101" => data_out <= rom_array(28429);
		when "0110111100001110" => data_out <= rom_array(28430);
		when "0110111100001111" => data_out <= rom_array(28431);
		when "0110111100010000" => data_out <= rom_array(28432);
		when "0110111100010001" => data_out <= rom_array(28433);
		when "0110111100010010" => data_out <= rom_array(28434);
		when "0110111100010011" => data_out <= rom_array(28435);
		when "0110111100010100" => data_out <= rom_array(28436);
		when "0110111100010101" => data_out <= rom_array(28437);
		when "0110111100010110" => data_out <= rom_array(28438);
		when "0110111100010111" => data_out <= rom_array(28439);
		when "0110111100011000" => data_out <= rom_array(28440);
		when "0110111100011001" => data_out <= rom_array(28441);
		when "0110111100011010" => data_out <= rom_array(28442);
		when "0110111100011011" => data_out <= rom_array(28443);
		when "0110111100011100" => data_out <= rom_array(28444);
		when "0110111100011101" => data_out <= rom_array(28445);
		when "0110111100011110" => data_out <= rom_array(28446);
		when "0110111100011111" => data_out <= rom_array(28447);
		when "0110111100100000" => data_out <= rom_array(28448);
		when "0110111100100001" => data_out <= rom_array(28449);
		when "0110111100100010" => data_out <= rom_array(28450);
		when "0110111100100011" => data_out <= rom_array(28451);
		when "0110111100100100" => data_out <= rom_array(28452);
		when "0110111100100101" => data_out <= rom_array(28453);
		when "0110111100100110" => data_out <= rom_array(28454);
		when "0110111100100111" => data_out <= rom_array(28455);
		when "0110111100101000" => data_out <= rom_array(28456);
		when "0110111100101001" => data_out <= rom_array(28457);
		when "0110111100101010" => data_out <= rom_array(28458);
		when "0110111100101011" => data_out <= rom_array(28459);
		when "0110111100101100" => data_out <= rom_array(28460);
		when "0110111100101101" => data_out <= rom_array(28461);
		when "0110111100101110" => data_out <= rom_array(28462);
		when "0110111100101111" => data_out <= rom_array(28463);
		when "0110111100110000" => data_out <= rom_array(28464);
		when "0110111100110001" => data_out <= rom_array(28465);
		when "0110111100110010" => data_out <= rom_array(28466);
		when "0110111100110011" => data_out <= rom_array(28467);
		when "0110111100110100" => data_out <= rom_array(28468);
		when "0110111100110101" => data_out <= rom_array(28469);
		when "0110111100110110" => data_out <= rom_array(28470);
		when "0110111100110111" => data_out <= rom_array(28471);
		when "0110111100111000" => data_out <= rom_array(28472);
		when "0110111100111001" => data_out <= rom_array(28473);
		when "0110111100111010" => data_out <= rom_array(28474);
		when "0110111100111011" => data_out <= rom_array(28475);
		when "0110111100111100" => data_out <= rom_array(28476);
		when "0110111100111101" => data_out <= rom_array(28477);
		when "0110111100111110" => data_out <= rom_array(28478);
		when "0110111100111111" => data_out <= rom_array(28479);
		when "0110111101000000" => data_out <= rom_array(28480);
		when "0110111101000001" => data_out <= rom_array(28481);
		when "0110111101000010" => data_out <= rom_array(28482);
		when "0110111101000011" => data_out <= rom_array(28483);
		when "0110111101000100" => data_out <= rom_array(28484);
		when "0110111101000101" => data_out <= rom_array(28485);
		when "0110111101000110" => data_out <= rom_array(28486);
		when "0110111101000111" => data_out <= rom_array(28487);
		when "0110111101001000" => data_out <= rom_array(28488);
		when "0110111101001001" => data_out <= rom_array(28489);
		when "0110111101001010" => data_out <= rom_array(28490);
		when "0110111101001011" => data_out <= rom_array(28491);
		when "0110111101001100" => data_out <= rom_array(28492);
		when "0110111101001101" => data_out <= rom_array(28493);
		when "0110111101001110" => data_out <= rom_array(28494);
		when "0110111101001111" => data_out <= rom_array(28495);
		when "0110111101010000" => data_out <= rom_array(28496);
		when "0110111101010001" => data_out <= rom_array(28497);
		when "0110111101010010" => data_out <= rom_array(28498);
		when "0110111101010011" => data_out <= rom_array(28499);
		when "0110111101010100" => data_out <= rom_array(28500);
		when "0110111101010101" => data_out <= rom_array(28501);
		when "0110111101010110" => data_out <= rom_array(28502);
		when "0110111101010111" => data_out <= rom_array(28503);
		when "0110111101011000" => data_out <= rom_array(28504);
		when "0110111101011001" => data_out <= rom_array(28505);
		when "0110111101011010" => data_out <= rom_array(28506);
		when "0110111101011011" => data_out <= rom_array(28507);
		when "0110111101011100" => data_out <= rom_array(28508);
		when "0110111101011101" => data_out <= rom_array(28509);
		when "0110111101011110" => data_out <= rom_array(28510);
		when "0110111101011111" => data_out <= rom_array(28511);
		when "0110111101100000" => data_out <= rom_array(28512);
		when "0110111101100001" => data_out <= rom_array(28513);
		when "0110111101100010" => data_out <= rom_array(28514);
		when "0110111101100011" => data_out <= rom_array(28515);
		when "0110111101100100" => data_out <= rom_array(28516);
		when "0110111101100101" => data_out <= rom_array(28517);
		when "0110111101100110" => data_out <= rom_array(28518);
		when "0110111101100111" => data_out <= rom_array(28519);
		when "0110111101101000" => data_out <= rom_array(28520);
		when "0110111101101001" => data_out <= rom_array(28521);
		when "0110111101101010" => data_out <= rom_array(28522);
		when "0110111101101011" => data_out <= rom_array(28523);
		when "0110111101101100" => data_out <= rom_array(28524);
		when "0110111101101101" => data_out <= rom_array(28525);
		when "0110111101101110" => data_out <= rom_array(28526);
		when "0110111101101111" => data_out <= rom_array(28527);
		when "0110111101110000" => data_out <= rom_array(28528);
		when "0110111101110001" => data_out <= rom_array(28529);
		when "0110111101110010" => data_out <= rom_array(28530);
		when "0110111101110011" => data_out <= rom_array(28531);
		when "0110111101110100" => data_out <= rom_array(28532);
		when "0110111101110101" => data_out <= rom_array(28533);
		when "0110111101110110" => data_out <= rom_array(28534);
		when "0110111101110111" => data_out <= rom_array(28535);
		when "0110111101111000" => data_out <= rom_array(28536);
		when "0110111101111001" => data_out <= rom_array(28537);
		when "0110111101111010" => data_out <= rom_array(28538);
		when "0110111101111011" => data_out <= rom_array(28539);
		when "0110111101111100" => data_out <= rom_array(28540);
		when "0110111101111101" => data_out <= rom_array(28541);
		when "0110111101111110" => data_out <= rom_array(28542);
		when "0110111101111111" => data_out <= rom_array(28543);
		when "0110111110000000" => data_out <= rom_array(28544);
		when "0110111110000001" => data_out <= rom_array(28545);
		when "0110111110000010" => data_out <= rom_array(28546);
		when "0110111110000011" => data_out <= rom_array(28547);
		when "0110111110000100" => data_out <= rom_array(28548);
		when "0110111110000101" => data_out <= rom_array(28549);
		when "0110111110000110" => data_out <= rom_array(28550);
		when "0110111110000111" => data_out <= rom_array(28551);
		when "0110111110001000" => data_out <= rom_array(28552);
		when "0110111110001001" => data_out <= rom_array(28553);
		when "0110111110001010" => data_out <= rom_array(28554);
		when "0110111110001011" => data_out <= rom_array(28555);
		when "0110111110001100" => data_out <= rom_array(28556);
		when "0110111110001101" => data_out <= rom_array(28557);
		when "0110111110001110" => data_out <= rom_array(28558);
		when "0110111110001111" => data_out <= rom_array(28559);
		when "0110111110010000" => data_out <= rom_array(28560);
		when "0110111110010001" => data_out <= rom_array(28561);
		when "0110111110010010" => data_out <= rom_array(28562);
		when "0110111110010011" => data_out <= rom_array(28563);
		when "0110111110010100" => data_out <= rom_array(28564);
		when "0110111110010101" => data_out <= rom_array(28565);
		when "0110111110010110" => data_out <= rom_array(28566);
		when "0110111110010111" => data_out <= rom_array(28567);
		when "0110111110011000" => data_out <= rom_array(28568);
		when "0110111110011001" => data_out <= rom_array(28569);
		when "0110111110011010" => data_out <= rom_array(28570);
		when "0110111110011011" => data_out <= rom_array(28571);
		when "0110111110011100" => data_out <= rom_array(28572);
		when "0110111110011101" => data_out <= rom_array(28573);
		when "0110111110011110" => data_out <= rom_array(28574);
		when "0110111110011111" => data_out <= rom_array(28575);
		when "0110111110100000" => data_out <= rom_array(28576);
		when "0110111110100001" => data_out <= rom_array(28577);
		when "0110111110100010" => data_out <= rom_array(28578);
		when "0110111110100011" => data_out <= rom_array(28579);
		when "0110111110100100" => data_out <= rom_array(28580);
		when "0110111110100101" => data_out <= rom_array(28581);
		when "0110111110100110" => data_out <= rom_array(28582);
		when "0110111110100111" => data_out <= rom_array(28583);
		when "0110111110101000" => data_out <= rom_array(28584);
		when "0110111110101001" => data_out <= rom_array(28585);
		when "0110111110101010" => data_out <= rom_array(28586);
		when "0110111110101011" => data_out <= rom_array(28587);
		when "0110111110101100" => data_out <= rom_array(28588);
		when "0110111110101101" => data_out <= rom_array(28589);
		when "0110111110101110" => data_out <= rom_array(28590);
		when "0110111110101111" => data_out <= rom_array(28591);
		when "0110111110110000" => data_out <= rom_array(28592);
		when "0110111110110001" => data_out <= rom_array(28593);
		when "0110111110110010" => data_out <= rom_array(28594);
		when "0110111110110011" => data_out <= rom_array(28595);
		when "0110111110110100" => data_out <= rom_array(28596);
		when "0110111110110101" => data_out <= rom_array(28597);
		when "0110111110110110" => data_out <= rom_array(28598);
		when "0110111110110111" => data_out <= rom_array(28599);
		when "0110111110111000" => data_out <= rom_array(28600);
		when "0110111110111001" => data_out <= rom_array(28601);
		when "0110111110111010" => data_out <= rom_array(28602);
		when "0110111110111011" => data_out <= rom_array(28603);
		when "0110111110111100" => data_out <= rom_array(28604);
		when "0110111110111101" => data_out <= rom_array(28605);
		when "0110111110111110" => data_out <= rom_array(28606);
		when "0110111110111111" => data_out <= rom_array(28607);
		when "0110111111000000" => data_out <= rom_array(28608);
		when "0110111111000001" => data_out <= rom_array(28609);
		when "0110111111000010" => data_out <= rom_array(28610);
		when "0110111111000011" => data_out <= rom_array(28611);
		when "0110111111000100" => data_out <= rom_array(28612);
		when "0110111111000101" => data_out <= rom_array(28613);
		when "0110111111000110" => data_out <= rom_array(28614);
		when "0110111111000111" => data_out <= rom_array(28615);
		when "0110111111001000" => data_out <= rom_array(28616);
		when "0110111111001001" => data_out <= rom_array(28617);
		when "0110111111001010" => data_out <= rom_array(28618);
		when "0110111111001011" => data_out <= rom_array(28619);
		when "0110111111001100" => data_out <= rom_array(28620);
		when "0110111111001101" => data_out <= rom_array(28621);
		when "0110111111001110" => data_out <= rom_array(28622);
		when "0110111111001111" => data_out <= rom_array(28623);
		when "0110111111010000" => data_out <= rom_array(28624);
		when "0110111111010001" => data_out <= rom_array(28625);
		when "0110111111010010" => data_out <= rom_array(28626);
		when "0110111111010011" => data_out <= rom_array(28627);
		when "0110111111010100" => data_out <= rom_array(28628);
		when "0110111111010101" => data_out <= rom_array(28629);
		when "0110111111010110" => data_out <= rom_array(28630);
		when "0110111111010111" => data_out <= rom_array(28631);
		when "0110111111011000" => data_out <= rom_array(28632);
		when "0110111111011001" => data_out <= rom_array(28633);
		when "0110111111011010" => data_out <= rom_array(28634);
		when "0110111111011011" => data_out <= rom_array(28635);
		when "0110111111011100" => data_out <= rom_array(28636);
		when "0110111111011101" => data_out <= rom_array(28637);
		when "0110111111011110" => data_out <= rom_array(28638);
		when "0110111111011111" => data_out <= rom_array(28639);
		when "0110111111100000" => data_out <= rom_array(28640);
		when "0110111111100001" => data_out <= rom_array(28641);
		when "0110111111100010" => data_out <= rom_array(28642);
		when "0110111111100011" => data_out <= rom_array(28643);
		when "0110111111100100" => data_out <= rom_array(28644);
		when "0110111111100101" => data_out <= rom_array(28645);
		when "0110111111100110" => data_out <= rom_array(28646);
		when "0110111111100111" => data_out <= rom_array(28647);
		when "0110111111101000" => data_out <= rom_array(28648);
		when "0110111111101001" => data_out <= rom_array(28649);
		when "0110111111101010" => data_out <= rom_array(28650);
		when "0110111111101011" => data_out <= rom_array(28651);
		when "0110111111101100" => data_out <= rom_array(28652);
		when "0110111111101101" => data_out <= rom_array(28653);
		when "0110111111101110" => data_out <= rom_array(28654);
		when "0110111111101111" => data_out <= rom_array(28655);
		when "0110111111110000" => data_out <= rom_array(28656);
		when "0110111111110001" => data_out <= rom_array(28657);
		when "0110111111110010" => data_out <= rom_array(28658);
		when "0110111111110011" => data_out <= rom_array(28659);
		when "0110111111110100" => data_out <= rom_array(28660);
		when "0110111111110101" => data_out <= rom_array(28661);
		when "0110111111110110" => data_out <= rom_array(28662);
		when "0110111111110111" => data_out <= rom_array(28663);
		when "0110111111111000" => data_out <= rom_array(28664);
		when "0110111111111001" => data_out <= rom_array(28665);
		when "0110111111111010" => data_out <= rom_array(28666);
		when "0110111111111011" => data_out <= rom_array(28667);
		when "0110111111111100" => data_out <= rom_array(28668);
		when "0110111111111101" => data_out <= rom_array(28669);
		when "0110111111111110" => data_out <= rom_array(28670);
		when "0110111111111111" => data_out <= rom_array(28671);
		when "0111000000000000" => data_out <= rom_array(28672);
		when "0111000000000001" => data_out <= rom_array(28673);
		when "0111000000000010" => data_out <= rom_array(28674);
		when "0111000000000011" => data_out <= rom_array(28675);
		when "0111000000000100" => data_out <= rom_array(28676);
		when "0111000000000101" => data_out <= rom_array(28677);
		when "0111000000000110" => data_out <= rom_array(28678);
		when "0111000000000111" => data_out <= rom_array(28679);
		when "0111000000001000" => data_out <= rom_array(28680);
		when "0111000000001001" => data_out <= rom_array(28681);
		when "0111000000001010" => data_out <= rom_array(28682);
		when "0111000000001011" => data_out <= rom_array(28683);
		when "0111000000001100" => data_out <= rom_array(28684);
		when "0111000000001101" => data_out <= rom_array(28685);
		when "0111000000001110" => data_out <= rom_array(28686);
		when "0111000000001111" => data_out <= rom_array(28687);
		when "0111000000010000" => data_out <= rom_array(28688);
		when "0111000000010001" => data_out <= rom_array(28689);
		when "0111000000010010" => data_out <= rom_array(28690);
		when "0111000000010011" => data_out <= rom_array(28691);
		when "0111000000010100" => data_out <= rom_array(28692);
		when "0111000000010101" => data_out <= rom_array(28693);
		when "0111000000010110" => data_out <= rom_array(28694);
		when "0111000000010111" => data_out <= rom_array(28695);
		when "0111000000011000" => data_out <= rom_array(28696);
		when "0111000000011001" => data_out <= rom_array(28697);
		when "0111000000011010" => data_out <= rom_array(28698);
		when "0111000000011011" => data_out <= rom_array(28699);
		when "0111000000011100" => data_out <= rom_array(28700);
		when "0111000000011101" => data_out <= rom_array(28701);
		when "0111000000011110" => data_out <= rom_array(28702);
		when "0111000000011111" => data_out <= rom_array(28703);
		when "0111000000100000" => data_out <= rom_array(28704);
		when "0111000000100001" => data_out <= rom_array(28705);
		when "0111000000100010" => data_out <= rom_array(28706);
		when "0111000000100011" => data_out <= rom_array(28707);
		when "0111000000100100" => data_out <= rom_array(28708);
		when "0111000000100101" => data_out <= rom_array(28709);
		when "0111000000100110" => data_out <= rom_array(28710);
		when "0111000000100111" => data_out <= rom_array(28711);
		when "0111000000101000" => data_out <= rom_array(28712);
		when "0111000000101001" => data_out <= rom_array(28713);
		when "0111000000101010" => data_out <= rom_array(28714);
		when "0111000000101011" => data_out <= rom_array(28715);
		when "0111000000101100" => data_out <= rom_array(28716);
		when "0111000000101101" => data_out <= rom_array(28717);
		when "0111000000101110" => data_out <= rom_array(28718);
		when "0111000000101111" => data_out <= rom_array(28719);
		when "0111000000110000" => data_out <= rom_array(28720);
		when "0111000000110001" => data_out <= rom_array(28721);
		when "0111000000110010" => data_out <= rom_array(28722);
		when "0111000000110011" => data_out <= rom_array(28723);
		when "0111000000110100" => data_out <= rom_array(28724);
		when "0111000000110101" => data_out <= rom_array(28725);
		when "0111000000110110" => data_out <= rom_array(28726);
		when "0111000000110111" => data_out <= rom_array(28727);
		when "0111000000111000" => data_out <= rom_array(28728);
		when "0111000000111001" => data_out <= rom_array(28729);
		when "0111000000111010" => data_out <= rom_array(28730);
		when "0111000000111011" => data_out <= rom_array(28731);
		when "0111000000111100" => data_out <= rom_array(28732);
		when "0111000000111101" => data_out <= rom_array(28733);
		when "0111000000111110" => data_out <= rom_array(28734);
		when "0111000000111111" => data_out <= rom_array(28735);
		when "0111000001000000" => data_out <= rom_array(28736);
		when "0111000001000001" => data_out <= rom_array(28737);
		when "0111000001000010" => data_out <= rom_array(28738);
		when "0111000001000011" => data_out <= rom_array(28739);
		when "0111000001000100" => data_out <= rom_array(28740);
		when "0111000001000101" => data_out <= rom_array(28741);
		when "0111000001000110" => data_out <= rom_array(28742);
		when "0111000001000111" => data_out <= rom_array(28743);
		when "0111000001001000" => data_out <= rom_array(28744);
		when "0111000001001001" => data_out <= rom_array(28745);
		when "0111000001001010" => data_out <= rom_array(28746);
		when "0111000001001011" => data_out <= rom_array(28747);
		when "0111000001001100" => data_out <= rom_array(28748);
		when "0111000001001101" => data_out <= rom_array(28749);
		when "0111000001001110" => data_out <= rom_array(28750);
		when "0111000001001111" => data_out <= rom_array(28751);
		when "0111000001010000" => data_out <= rom_array(28752);
		when "0111000001010001" => data_out <= rom_array(28753);
		when "0111000001010010" => data_out <= rom_array(28754);
		when "0111000001010011" => data_out <= rom_array(28755);
		when "0111000001010100" => data_out <= rom_array(28756);
		when "0111000001010101" => data_out <= rom_array(28757);
		when "0111000001010110" => data_out <= rom_array(28758);
		when "0111000001010111" => data_out <= rom_array(28759);
		when "0111000001011000" => data_out <= rom_array(28760);
		when "0111000001011001" => data_out <= rom_array(28761);
		when "0111000001011010" => data_out <= rom_array(28762);
		when "0111000001011011" => data_out <= rom_array(28763);
		when "0111000001011100" => data_out <= rom_array(28764);
		when "0111000001011101" => data_out <= rom_array(28765);
		when "0111000001011110" => data_out <= rom_array(28766);
		when "0111000001011111" => data_out <= rom_array(28767);
		when "0111000001100000" => data_out <= rom_array(28768);
		when "0111000001100001" => data_out <= rom_array(28769);
		when "0111000001100010" => data_out <= rom_array(28770);
		when "0111000001100011" => data_out <= rom_array(28771);
		when "0111000001100100" => data_out <= rom_array(28772);
		when "0111000001100101" => data_out <= rom_array(28773);
		when "0111000001100110" => data_out <= rom_array(28774);
		when "0111000001100111" => data_out <= rom_array(28775);
		when "0111000001101000" => data_out <= rom_array(28776);
		when "0111000001101001" => data_out <= rom_array(28777);
		when "0111000001101010" => data_out <= rom_array(28778);
		when "0111000001101011" => data_out <= rom_array(28779);
		when "0111000001101100" => data_out <= rom_array(28780);
		when "0111000001101101" => data_out <= rom_array(28781);
		when "0111000001101110" => data_out <= rom_array(28782);
		when "0111000001101111" => data_out <= rom_array(28783);
		when "0111000001110000" => data_out <= rom_array(28784);
		when "0111000001110001" => data_out <= rom_array(28785);
		when "0111000001110010" => data_out <= rom_array(28786);
		when "0111000001110011" => data_out <= rom_array(28787);
		when "0111000001110100" => data_out <= rom_array(28788);
		when "0111000001110101" => data_out <= rom_array(28789);
		when "0111000001110110" => data_out <= rom_array(28790);
		when "0111000001110111" => data_out <= rom_array(28791);
		when "0111000001111000" => data_out <= rom_array(28792);
		when "0111000001111001" => data_out <= rom_array(28793);
		when "0111000001111010" => data_out <= rom_array(28794);
		when "0111000001111011" => data_out <= rom_array(28795);
		when "0111000001111100" => data_out <= rom_array(28796);
		when "0111000001111101" => data_out <= rom_array(28797);
		when "0111000001111110" => data_out <= rom_array(28798);
		when "0111000001111111" => data_out <= rom_array(28799);
		when "0111000010000000" => data_out <= rom_array(28800);
		when "0111000010000001" => data_out <= rom_array(28801);
		when "0111000010000010" => data_out <= rom_array(28802);
		when "0111000010000011" => data_out <= rom_array(28803);
		when "0111000010000100" => data_out <= rom_array(28804);
		when "0111000010000101" => data_out <= rom_array(28805);
		when "0111000010000110" => data_out <= rom_array(28806);
		when "0111000010000111" => data_out <= rom_array(28807);
		when "0111000010001000" => data_out <= rom_array(28808);
		when "0111000010001001" => data_out <= rom_array(28809);
		when "0111000010001010" => data_out <= rom_array(28810);
		when "0111000010001011" => data_out <= rom_array(28811);
		when "0111000010001100" => data_out <= rom_array(28812);
		when "0111000010001101" => data_out <= rom_array(28813);
		when "0111000010001110" => data_out <= rom_array(28814);
		when "0111000010001111" => data_out <= rom_array(28815);
		when "0111000010010000" => data_out <= rom_array(28816);
		when "0111000010010001" => data_out <= rom_array(28817);
		when "0111000010010010" => data_out <= rom_array(28818);
		when "0111000010010011" => data_out <= rom_array(28819);
		when "0111000010010100" => data_out <= rom_array(28820);
		when "0111000010010101" => data_out <= rom_array(28821);
		when "0111000010010110" => data_out <= rom_array(28822);
		when "0111000010010111" => data_out <= rom_array(28823);
		when "0111000010011000" => data_out <= rom_array(28824);
		when "0111000010011001" => data_out <= rom_array(28825);
		when "0111000010011010" => data_out <= rom_array(28826);
		when "0111000010011011" => data_out <= rom_array(28827);
		when "0111000010011100" => data_out <= rom_array(28828);
		when "0111000010011101" => data_out <= rom_array(28829);
		when "0111000010011110" => data_out <= rom_array(28830);
		when "0111000010011111" => data_out <= rom_array(28831);
		when "0111000010100000" => data_out <= rom_array(28832);
		when "0111000010100001" => data_out <= rom_array(28833);
		when "0111000010100010" => data_out <= rom_array(28834);
		when "0111000010100011" => data_out <= rom_array(28835);
		when "0111000010100100" => data_out <= rom_array(28836);
		when "0111000010100101" => data_out <= rom_array(28837);
		when "0111000010100110" => data_out <= rom_array(28838);
		when "0111000010100111" => data_out <= rom_array(28839);
		when "0111000010101000" => data_out <= rom_array(28840);
		when "0111000010101001" => data_out <= rom_array(28841);
		when "0111000010101010" => data_out <= rom_array(28842);
		when "0111000010101011" => data_out <= rom_array(28843);
		when "0111000010101100" => data_out <= rom_array(28844);
		when "0111000010101101" => data_out <= rom_array(28845);
		when "0111000010101110" => data_out <= rom_array(28846);
		when "0111000010101111" => data_out <= rom_array(28847);
		when "0111000010110000" => data_out <= rom_array(28848);
		when "0111000010110001" => data_out <= rom_array(28849);
		when "0111000010110010" => data_out <= rom_array(28850);
		when "0111000010110011" => data_out <= rom_array(28851);
		when "0111000010110100" => data_out <= rom_array(28852);
		when "0111000010110101" => data_out <= rom_array(28853);
		when "0111000010110110" => data_out <= rom_array(28854);
		when "0111000010110111" => data_out <= rom_array(28855);
		when "0111000010111000" => data_out <= rom_array(28856);
		when "0111000010111001" => data_out <= rom_array(28857);
		when "0111000010111010" => data_out <= rom_array(28858);
		when "0111000010111011" => data_out <= rom_array(28859);
		when "0111000010111100" => data_out <= rom_array(28860);
		when "0111000010111101" => data_out <= rom_array(28861);
		when "0111000010111110" => data_out <= rom_array(28862);
		when "0111000010111111" => data_out <= rom_array(28863);
		when "0111000011000000" => data_out <= rom_array(28864);
		when "0111000011000001" => data_out <= rom_array(28865);
		when "0111000011000010" => data_out <= rom_array(28866);
		when "0111000011000011" => data_out <= rom_array(28867);
		when "0111000011000100" => data_out <= rom_array(28868);
		when "0111000011000101" => data_out <= rom_array(28869);
		when "0111000011000110" => data_out <= rom_array(28870);
		when "0111000011000111" => data_out <= rom_array(28871);
		when "0111000011001000" => data_out <= rom_array(28872);
		when "0111000011001001" => data_out <= rom_array(28873);
		when "0111000011001010" => data_out <= rom_array(28874);
		when "0111000011001011" => data_out <= rom_array(28875);
		when "0111000011001100" => data_out <= rom_array(28876);
		when "0111000011001101" => data_out <= rom_array(28877);
		when "0111000011001110" => data_out <= rom_array(28878);
		when "0111000011001111" => data_out <= rom_array(28879);
		when "0111000011010000" => data_out <= rom_array(28880);
		when "0111000011010001" => data_out <= rom_array(28881);
		when "0111000011010010" => data_out <= rom_array(28882);
		when "0111000011010011" => data_out <= rom_array(28883);
		when "0111000011010100" => data_out <= rom_array(28884);
		when "0111000011010101" => data_out <= rom_array(28885);
		when "0111000011010110" => data_out <= rom_array(28886);
		when "0111000011010111" => data_out <= rom_array(28887);
		when "0111000011011000" => data_out <= rom_array(28888);
		when "0111000011011001" => data_out <= rom_array(28889);
		when "0111000011011010" => data_out <= rom_array(28890);
		when "0111000011011011" => data_out <= rom_array(28891);
		when "0111000011011100" => data_out <= rom_array(28892);
		when "0111000011011101" => data_out <= rom_array(28893);
		when "0111000011011110" => data_out <= rom_array(28894);
		when "0111000011011111" => data_out <= rom_array(28895);
		when "0111000011100000" => data_out <= rom_array(28896);
		when "0111000011100001" => data_out <= rom_array(28897);
		when "0111000011100010" => data_out <= rom_array(28898);
		when "0111000011100011" => data_out <= rom_array(28899);
		when "0111000011100100" => data_out <= rom_array(28900);
		when "0111000011100101" => data_out <= rom_array(28901);
		when "0111000011100110" => data_out <= rom_array(28902);
		when "0111000011100111" => data_out <= rom_array(28903);
		when "0111000011101000" => data_out <= rom_array(28904);
		when "0111000011101001" => data_out <= rom_array(28905);
		when "0111000011101010" => data_out <= rom_array(28906);
		when "0111000011101011" => data_out <= rom_array(28907);
		when "0111000011101100" => data_out <= rom_array(28908);
		when "0111000011101101" => data_out <= rom_array(28909);
		when "0111000011101110" => data_out <= rom_array(28910);
		when "0111000011101111" => data_out <= rom_array(28911);
		when "0111000011110000" => data_out <= rom_array(28912);
		when "0111000011110001" => data_out <= rom_array(28913);
		when "0111000011110010" => data_out <= rom_array(28914);
		when "0111000011110011" => data_out <= rom_array(28915);
		when "0111000011110100" => data_out <= rom_array(28916);
		when "0111000011110101" => data_out <= rom_array(28917);
		when "0111000011110110" => data_out <= rom_array(28918);
		when "0111000011110111" => data_out <= rom_array(28919);
		when "0111000011111000" => data_out <= rom_array(28920);
		when "0111000011111001" => data_out <= rom_array(28921);
		when "0111000011111010" => data_out <= rom_array(28922);
		when "0111000011111011" => data_out <= rom_array(28923);
		when "0111000011111100" => data_out <= rom_array(28924);
		when "0111000011111101" => data_out <= rom_array(28925);
		when "0111000011111110" => data_out <= rom_array(28926);
		when "0111000011111111" => data_out <= rom_array(28927);
		when "0111000100000000" => data_out <= rom_array(28928);
		when "0111000100000001" => data_out <= rom_array(28929);
		when "0111000100000010" => data_out <= rom_array(28930);
		when "0111000100000011" => data_out <= rom_array(28931);
		when "0111000100000100" => data_out <= rom_array(28932);
		when "0111000100000101" => data_out <= rom_array(28933);
		when "0111000100000110" => data_out <= rom_array(28934);
		when "0111000100000111" => data_out <= rom_array(28935);
		when "0111000100001000" => data_out <= rom_array(28936);
		when "0111000100001001" => data_out <= rom_array(28937);
		when "0111000100001010" => data_out <= rom_array(28938);
		when "0111000100001011" => data_out <= rom_array(28939);
		when "0111000100001100" => data_out <= rom_array(28940);
		when "0111000100001101" => data_out <= rom_array(28941);
		when "0111000100001110" => data_out <= rom_array(28942);
		when "0111000100001111" => data_out <= rom_array(28943);
		when "0111000100010000" => data_out <= rom_array(28944);
		when "0111000100010001" => data_out <= rom_array(28945);
		when "0111000100010010" => data_out <= rom_array(28946);
		when "0111000100010011" => data_out <= rom_array(28947);
		when "0111000100010100" => data_out <= rom_array(28948);
		when "0111000100010101" => data_out <= rom_array(28949);
		when "0111000100010110" => data_out <= rom_array(28950);
		when "0111000100010111" => data_out <= rom_array(28951);
		when "0111000100011000" => data_out <= rom_array(28952);
		when "0111000100011001" => data_out <= rom_array(28953);
		when "0111000100011010" => data_out <= rom_array(28954);
		when "0111000100011011" => data_out <= rom_array(28955);
		when "0111000100011100" => data_out <= rom_array(28956);
		when "0111000100011101" => data_out <= rom_array(28957);
		when "0111000100011110" => data_out <= rom_array(28958);
		when "0111000100011111" => data_out <= rom_array(28959);
		when "0111000100100000" => data_out <= rom_array(28960);
		when "0111000100100001" => data_out <= rom_array(28961);
		when "0111000100100010" => data_out <= rom_array(28962);
		when "0111000100100011" => data_out <= rom_array(28963);
		when "0111000100100100" => data_out <= rom_array(28964);
		when "0111000100100101" => data_out <= rom_array(28965);
		when "0111000100100110" => data_out <= rom_array(28966);
		when "0111000100100111" => data_out <= rom_array(28967);
		when "0111000100101000" => data_out <= rom_array(28968);
		when "0111000100101001" => data_out <= rom_array(28969);
		when "0111000100101010" => data_out <= rom_array(28970);
		when "0111000100101011" => data_out <= rom_array(28971);
		when "0111000100101100" => data_out <= rom_array(28972);
		when "0111000100101101" => data_out <= rom_array(28973);
		when "0111000100101110" => data_out <= rom_array(28974);
		when "0111000100101111" => data_out <= rom_array(28975);
		when "0111000100110000" => data_out <= rom_array(28976);
		when "0111000100110001" => data_out <= rom_array(28977);
		when "0111000100110010" => data_out <= rom_array(28978);
		when "0111000100110011" => data_out <= rom_array(28979);
		when "0111000100110100" => data_out <= rom_array(28980);
		when "0111000100110101" => data_out <= rom_array(28981);
		when "0111000100110110" => data_out <= rom_array(28982);
		when "0111000100110111" => data_out <= rom_array(28983);
		when "0111000100111000" => data_out <= rom_array(28984);
		when "0111000100111001" => data_out <= rom_array(28985);
		when "0111000100111010" => data_out <= rom_array(28986);
		when "0111000100111011" => data_out <= rom_array(28987);
		when "0111000100111100" => data_out <= rom_array(28988);
		when "0111000100111101" => data_out <= rom_array(28989);
		when "0111000100111110" => data_out <= rom_array(28990);
		when "0111000100111111" => data_out <= rom_array(28991);
		when "0111000101000000" => data_out <= rom_array(28992);
		when "0111000101000001" => data_out <= rom_array(28993);
		when "0111000101000010" => data_out <= rom_array(28994);
		when "0111000101000011" => data_out <= rom_array(28995);
		when "0111000101000100" => data_out <= rom_array(28996);
		when "0111000101000101" => data_out <= rom_array(28997);
		when "0111000101000110" => data_out <= rom_array(28998);
		when "0111000101000111" => data_out <= rom_array(28999);
		when "0111000101001000" => data_out <= rom_array(29000);
		when "0111000101001001" => data_out <= rom_array(29001);
		when "0111000101001010" => data_out <= rom_array(29002);
		when "0111000101001011" => data_out <= rom_array(29003);
		when "0111000101001100" => data_out <= rom_array(29004);
		when "0111000101001101" => data_out <= rom_array(29005);
		when "0111000101001110" => data_out <= rom_array(29006);
		when "0111000101001111" => data_out <= rom_array(29007);
		when "0111000101010000" => data_out <= rom_array(29008);
		when "0111000101010001" => data_out <= rom_array(29009);
		when "0111000101010010" => data_out <= rom_array(29010);
		when "0111000101010011" => data_out <= rom_array(29011);
		when "0111000101010100" => data_out <= rom_array(29012);
		when "0111000101010101" => data_out <= rom_array(29013);
		when "0111000101010110" => data_out <= rom_array(29014);
		when "0111000101010111" => data_out <= rom_array(29015);
		when "0111000101011000" => data_out <= rom_array(29016);
		when "0111000101011001" => data_out <= rom_array(29017);
		when "0111000101011010" => data_out <= rom_array(29018);
		when "0111000101011011" => data_out <= rom_array(29019);
		when "0111000101011100" => data_out <= rom_array(29020);
		when "0111000101011101" => data_out <= rom_array(29021);
		when "0111000101011110" => data_out <= rom_array(29022);
		when "0111000101011111" => data_out <= rom_array(29023);
		when "0111000101100000" => data_out <= rom_array(29024);
		when "0111000101100001" => data_out <= rom_array(29025);
		when "0111000101100010" => data_out <= rom_array(29026);
		when "0111000101100011" => data_out <= rom_array(29027);
		when "0111000101100100" => data_out <= rom_array(29028);
		when "0111000101100101" => data_out <= rom_array(29029);
		when "0111000101100110" => data_out <= rom_array(29030);
		when "0111000101100111" => data_out <= rom_array(29031);
		when "0111000101101000" => data_out <= rom_array(29032);
		when "0111000101101001" => data_out <= rom_array(29033);
		when "0111000101101010" => data_out <= rom_array(29034);
		when "0111000101101011" => data_out <= rom_array(29035);
		when "0111000101101100" => data_out <= rom_array(29036);
		when "0111000101101101" => data_out <= rom_array(29037);
		when "0111000101101110" => data_out <= rom_array(29038);
		when "0111000101101111" => data_out <= rom_array(29039);
		when "0111000101110000" => data_out <= rom_array(29040);
		when "0111000101110001" => data_out <= rom_array(29041);
		when "0111000101110010" => data_out <= rom_array(29042);
		when "0111000101110011" => data_out <= rom_array(29043);
		when "0111000101110100" => data_out <= rom_array(29044);
		when "0111000101110101" => data_out <= rom_array(29045);
		when "0111000101110110" => data_out <= rom_array(29046);
		when "0111000101110111" => data_out <= rom_array(29047);
		when "0111000101111000" => data_out <= rom_array(29048);
		when "0111000101111001" => data_out <= rom_array(29049);
		when "0111000101111010" => data_out <= rom_array(29050);
		when "0111000101111011" => data_out <= rom_array(29051);
		when "0111000101111100" => data_out <= rom_array(29052);
		when "0111000101111101" => data_out <= rom_array(29053);
		when "0111000101111110" => data_out <= rom_array(29054);
		when "0111000101111111" => data_out <= rom_array(29055);
		when "0111000110000000" => data_out <= rom_array(29056);
		when "0111000110000001" => data_out <= rom_array(29057);
		when "0111000110000010" => data_out <= rom_array(29058);
		when "0111000110000011" => data_out <= rom_array(29059);
		when "0111000110000100" => data_out <= rom_array(29060);
		when "0111000110000101" => data_out <= rom_array(29061);
		when "0111000110000110" => data_out <= rom_array(29062);
		when "0111000110000111" => data_out <= rom_array(29063);
		when "0111000110001000" => data_out <= rom_array(29064);
		when "0111000110001001" => data_out <= rom_array(29065);
		when "0111000110001010" => data_out <= rom_array(29066);
		when "0111000110001011" => data_out <= rom_array(29067);
		when "0111000110001100" => data_out <= rom_array(29068);
		when "0111000110001101" => data_out <= rom_array(29069);
		when "0111000110001110" => data_out <= rom_array(29070);
		when "0111000110001111" => data_out <= rom_array(29071);
		when "0111000110010000" => data_out <= rom_array(29072);
		when "0111000110010001" => data_out <= rom_array(29073);
		when "0111000110010010" => data_out <= rom_array(29074);
		when "0111000110010011" => data_out <= rom_array(29075);
		when "0111000110010100" => data_out <= rom_array(29076);
		when "0111000110010101" => data_out <= rom_array(29077);
		when "0111000110010110" => data_out <= rom_array(29078);
		when "0111000110010111" => data_out <= rom_array(29079);
		when "0111000110011000" => data_out <= rom_array(29080);
		when "0111000110011001" => data_out <= rom_array(29081);
		when "0111000110011010" => data_out <= rom_array(29082);
		when "0111000110011011" => data_out <= rom_array(29083);
		when "0111000110011100" => data_out <= rom_array(29084);
		when "0111000110011101" => data_out <= rom_array(29085);
		when "0111000110011110" => data_out <= rom_array(29086);
		when "0111000110011111" => data_out <= rom_array(29087);
		when "0111000110100000" => data_out <= rom_array(29088);
		when "0111000110100001" => data_out <= rom_array(29089);
		when "0111000110100010" => data_out <= rom_array(29090);
		when "0111000110100011" => data_out <= rom_array(29091);
		when "0111000110100100" => data_out <= rom_array(29092);
		when "0111000110100101" => data_out <= rom_array(29093);
		when "0111000110100110" => data_out <= rom_array(29094);
		when "0111000110100111" => data_out <= rom_array(29095);
		when "0111000110101000" => data_out <= rom_array(29096);
		when "0111000110101001" => data_out <= rom_array(29097);
		when "0111000110101010" => data_out <= rom_array(29098);
		when "0111000110101011" => data_out <= rom_array(29099);
		when "0111000110101100" => data_out <= rom_array(29100);
		when "0111000110101101" => data_out <= rom_array(29101);
		when "0111000110101110" => data_out <= rom_array(29102);
		when "0111000110101111" => data_out <= rom_array(29103);
		when "0111000110110000" => data_out <= rom_array(29104);
		when "0111000110110001" => data_out <= rom_array(29105);
		when "0111000110110010" => data_out <= rom_array(29106);
		when "0111000110110011" => data_out <= rom_array(29107);
		when "0111000110110100" => data_out <= rom_array(29108);
		when "0111000110110101" => data_out <= rom_array(29109);
		when "0111000110110110" => data_out <= rom_array(29110);
		when "0111000110110111" => data_out <= rom_array(29111);
		when "0111000110111000" => data_out <= rom_array(29112);
		when "0111000110111001" => data_out <= rom_array(29113);
		when "0111000110111010" => data_out <= rom_array(29114);
		when "0111000110111011" => data_out <= rom_array(29115);
		when "0111000110111100" => data_out <= rom_array(29116);
		when "0111000110111101" => data_out <= rom_array(29117);
		when "0111000110111110" => data_out <= rom_array(29118);
		when "0111000110111111" => data_out <= rom_array(29119);
		when "0111000111000000" => data_out <= rom_array(29120);
		when "0111000111000001" => data_out <= rom_array(29121);
		when "0111000111000010" => data_out <= rom_array(29122);
		when "0111000111000011" => data_out <= rom_array(29123);
		when "0111000111000100" => data_out <= rom_array(29124);
		when "0111000111000101" => data_out <= rom_array(29125);
		when "0111000111000110" => data_out <= rom_array(29126);
		when "0111000111000111" => data_out <= rom_array(29127);
		when "0111000111001000" => data_out <= rom_array(29128);
		when "0111000111001001" => data_out <= rom_array(29129);
		when "0111000111001010" => data_out <= rom_array(29130);
		when "0111000111001011" => data_out <= rom_array(29131);
		when "0111000111001100" => data_out <= rom_array(29132);
		when "0111000111001101" => data_out <= rom_array(29133);
		when "0111000111001110" => data_out <= rom_array(29134);
		when "0111000111001111" => data_out <= rom_array(29135);
		when "0111000111010000" => data_out <= rom_array(29136);
		when "0111000111010001" => data_out <= rom_array(29137);
		when "0111000111010010" => data_out <= rom_array(29138);
		when "0111000111010011" => data_out <= rom_array(29139);
		when "0111000111010100" => data_out <= rom_array(29140);
		when "0111000111010101" => data_out <= rom_array(29141);
		when "0111000111010110" => data_out <= rom_array(29142);
		when "0111000111010111" => data_out <= rom_array(29143);
		when "0111000111011000" => data_out <= rom_array(29144);
		when "0111000111011001" => data_out <= rom_array(29145);
		when "0111000111011010" => data_out <= rom_array(29146);
		when "0111000111011011" => data_out <= rom_array(29147);
		when "0111000111011100" => data_out <= rom_array(29148);
		when "0111000111011101" => data_out <= rom_array(29149);
		when "0111000111011110" => data_out <= rom_array(29150);
		when "0111000111011111" => data_out <= rom_array(29151);
		when "0111000111100000" => data_out <= rom_array(29152);
		when "0111000111100001" => data_out <= rom_array(29153);
		when "0111000111100010" => data_out <= rom_array(29154);
		when "0111000111100011" => data_out <= rom_array(29155);
		when "0111000111100100" => data_out <= rom_array(29156);
		when "0111000111100101" => data_out <= rom_array(29157);
		when "0111000111100110" => data_out <= rom_array(29158);
		when "0111000111100111" => data_out <= rom_array(29159);
		when "0111000111101000" => data_out <= rom_array(29160);
		when "0111000111101001" => data_out <= rom_array(29161);
		when "0111000111101010" => data_out <= rom_array(29162);
		when "0111000111101011" => data_out <= rom_array(29163);
		when "0111000111101100" => data_out <= rom_array(29164);
		when "0111000111101101" => data_out <= rom_array(29165);
		when "0111000111101110" => data_out <= rom_array(29166);
		when "0111000111101111" => data_out <= rom_array(29167);
		when "0111000111110000" => data_out <= rom_array(29168);
		when "0111000111110001" => data_out <= rom_array(29169);
		when "0111000111110010" => data_out <= rom_array(29170);
		when "0111000111110011" => data_out <= rom_array(29171);
		when "0111000111110100" => data_out <= rom_array(29172);
		when "0111000111110101" => data_out <= rom_array(29173);
		when "0111000111110110" => data_out <= rom_array(29174);
		when "0111000111110111" => data_out <= rom_array(29175);
		when "0111000111111000" => data_out <= rom_array(29176);
		when "0111000111111001" => data_out <= rom_array(29177);
		when "0111000111111010" => data_out <= rom_array(29178);
		when "0111000111111011" => data_out <= rom_array(29179);
		when "0111000111111100" => data_out <= rom_array(29180);
		when "0111000111111101" => data_out <= rom_array(29181);
		when "0111000111111110" => data_out <= rom_array(29182);
		when "0111000111111111" => data_out <= rom_array(29183);
		when "0111001000000000" => data_out <= rom_array(29184);
		when "0111001000000001" => data_out <= rom_array(29185);
		when "0111001000000010" => data_out <= rom_array(29186);
		when "0111001000000011" => data_out <= rom_array(29187);
		when "0111001000000100" => data_out <= rom_array(29188);
		when "0111001000000101" => data_out <= rom_array(29189);
		when "0111001000000110" => data_out <= rom_array(29190);
		when "0111001000000111" => data_out <= rom_array(29191);
		when "0111001000001000" => data_out <= rom_array(29192);
		when "0111001000001001" => data_out <= rom_array(29193);
		when "0111001000001010" => data_out <= rom_array(29194);
		when "0111001000001011" => data_out <= rom_array(29195);
		when "0111001000001100" => data_out <= rom_array(29196);
		when "0111001000001101" => data_out <= rom_array(29197);
		when "0111001000001110" => data_out <= rom_array(29198);
		when "0111001000001111" => data_out <= rom_array(29199);
		when "0111001000010000" => data_out <= rom_array(29200);
		when "0111001000010001" => data_out <= rom_array(29201);
		when "0111001000010010" => data_out <= rom_array(29202);
		when "0111001000010011" => data_out <= rom_array(29203);
		when "0111001000010100" => data_out <= rom_array(29204);
		when "0111001000010101" => data_out <= rom_array(29205);
		when "0111001000010110" => data_out <= rom_array(29206);
		when "0111001000010111" => data_out <= rom_array(29207);
		when "0111001000011000" => data_out <= rom_array(29208);
		when "0111001000011001" => data_out <= rom_array(29209);
		when "0111001000011010" => data_out <= rom_array(29210);
		when "0111001000011011" => data_out <= rom_array(29211);
		when "0111001000011100" => data_out <= rom_array(29212);
		when "0111001000011101" => data_out <= rom_array(29213);
		when "0111001000011110" => data_out <= rom_array(29214);
		when "0111001000011111" => data_out <= rom_array(29215);
		when "0111001000100000" => data_out <= rom_array(29216);
		when "0111001000100001" => data_out <= rom_array(29217);
		when "0111001000100010" => data_out <= rom_array(29218);
		when "0111001000100011" => data_out <= rom_array(29219);
		when "0111001000100100" => data_out <= rom_array(29220);
		when "0111001000100101" => data_out <= rom_array(29221);
		when "0111001000100110" => data_out <= rom_array(29222);
		when "0111001000100111" => data_out <= rom_array(29223);
		when "0111001000101000" => data_out <= rom_array(29224);
		when "0111001000101001" => data_out <= rom_array(29225);
		when "0111001000101010" => data_out <= rom_array(29226);
		when "0111001000101011" => data_out <= rom_array(29227);
		when "0111001000101100" => data_out <= rom_array(29228);
		when "0111001000101101" => data_out <= rom_array(29229);
		when "0111001000101110" => data_out <= rom_array(29230);
		when "0111001000101111" => data_out <= rom_array(29231);
		when "0111001000110000" => data_out <= rom_array(29232);
		when "0111001000110001" => data_out <= rom_array(29233);
		when "0111001000110010" => data_out <= rom_array(29234);
		when "0111001000110011" => data_out <= rom_array(29235);
		when "0111001000110100" => data_out <= rom_array(29236);
		when "0111001000110101" => data_out <= rom_array(29237);
		when "0111001000110110" => data_out <= rom_array(29238);
		when "0111001000110111" => data_out <= rom_array(29239);
		when "0111001000111000" => data_out <= rom_array(29240);
		when "0111001000111001" => data_out <= rom_array(29241);
		when "0111001000111010" => data_out <= rom_array(29242);
		when "0111001000111011" => data_out <= rom_array(29243);
		when "0111001000111100" => data_out <= rom_array(29244);
		when "0111001000111101" => data_out <= rom_array(29245);
		when "0111001000111110" => data_out <= rom_array(29246);
		when "0111001000111111" => data_out <= rom_array(29247);
		when "0111001001000000" => data_out <= rom_array(29248);
		when "0111001001000001" => data_out <= rom_array(29249);
		when "0111001001000010" => data_out <= rom_array(29250);
		when "0111001001000011" => data_out <= rom_array(29251);
		when "0111001001000100" => data_out <= rom_array(29252);
		when "0111001001000101" => data_out <= rom_array(29253);
		when "0111001001000110" => data_out <= rom_array(29254);
		when "0111001001000111" => data_out <= rom_array(29255);
		when "0111001001001000" => data_out <= rom_array(29256);
		when "0111001001001001" => data_out <= rom_array(29257);
		when "0111001001001010" => data_out <= rom_array(29258);
		when "0111001001001011" => data_out <= rom_array(29259);
		when "0111001001001100" => data_out <= rom_array(29260);
		when "0111001001001101" => data_out <= rom_array(29261);
		when "0111001001001110" => data_out <= rom_array(29262);
		when "0111001001001111" => data_out <= rom_array(29263);
		when "0111001001010000" => data_out <= rom_array(29264);
		when "0111001001010001" => data_out <= rom_array(29265);
		when "0111001001010010" => data_out <= rom_array(29266);
		when "0111001001010011" => data_out <= rom_array(29267);
		when "0111001001010100" => data_out <= rom_array(29268);
		when "0111001001010101" => data_out <= rom_array(29269);
		when "0111001001010110" => data_out <= rom_array(29270);
		when "0111001001010111" => data_out <= rom_array(29271);
		when "0111001001011000" => data_out <= rom_array(29272);
		when "0111001001011001" => data_out <= rom_array(29273);
		when "0111001001011010" => data_out <= rom_array(29274);
		when "0111001001011011" => data_out <= rom_array(29275);
		when "0111001001011100" => data_out <= rom_array(29276);
		when "0111001001011101" => data_out <= rom_array(29277);
		when "0111001001011110" => data_out <= rom_array(29278);
		when "0111001001011111" => data_out <= rom_array(29279);
		when "0111001001100000" => data_out <= rom_array(29280);
		when "0111001001100001" => data_out <= rom_array(29281);
		when "0111001001100010" => data_out <= rom_array(29282);
		when "0111001001100011" => data_out <= rom_array(29283);
		when "0111001001100100" => data_out <= rom_array(29284);
		when "0111001001100101" => data_out <= rom_array(29285);
		when "0111001001100110" => data_out <= rom_array(29286);
		when "0111001001100111" => data_out <= rom_array(29287);
		when "0111001001101000" => data_out <= rom_array(29288);
		when "0111001001101001" => data_out <= rom_array(29289);
		when "0111001001101010" => data_out <= rom_array(29290);
		when "0111001001101011" => data_out <= rom_array(29291);
		when "0111001001101100" => data_out <= rom_array(29292);
		when "0111001001101101" => data_out <= rom_array(29293);
		when "0111001001101110" => data_out <= rom_array(29294);
		when "0111001001101111" => data_out <= rom_array(29295);
		when "0111001001110000" => data_out <= rom_array(29296);
		when "0111001001110001" => data_out <= rom_array(29297);
		when "0111001001110010" => data_out <= rom_array(29298);
		when "0111001001110011" => data_out <= rom_array(29299);
		when "0111001001110100" => data_out <= rom_array(29300);
		when "0111001001110101" => data_out <= rom_array(29301);
		when "0111001001110110" => data_out <= rom_array(29302);
		when "0111001001110111" => data_out <= rom_array(29303);
		when "0111001001111000" => data_out <= rom_array(29304);
		when "0111001001111001" => data_out <= rom_array(29305);
		when "0111001001111010" => data_out <= rom_array(29306);
		when "0111001001111011" => data_out <= rom_array(29307);
		when "0111001001111100" => data_out <= rom_array(29308);
		when "0111001001111101" => data_out <= rom_array(29309);
		when "0111001001111110" => data_out <= rom_array(29310);
		when "0111001001111111" => data_out <= rom_array(29311);
		when "0111001010000000" => data_out <= rom_array(29312);
		when "0111001010000001" => data_out <= rom_array(29313);
		when "0111001010000010" => data_out <= rom_array(29314);
		when "0111001010000011" => data_out <= rom_array(29315);
		when "0111001010000100" => data_out <= rom_array(29316);
		when "0111001010000101" => data_out <= rom_array(29317);
		when "0111001010000110" => data_out <= rom_array(29318);
		when "0111001010000111" => data_out <= rom_array(29319);
		when "0111001010001000" => data_out <= rom_array(29320);
		when "0111001010001001" => data_out <= rom_array(29321);
		when "0111001010001010" => data_out <= rom_array(29322);
		when "0111001010001011" => data_out <= rom_array(29323);
		when "0111001010001100" => data_out <= rom_array(29324);
		when "0111001010001101" => data_out <= rom_array(29325);
		when "0111001010001110" => data_out <= rom_array(29326);
		when "0111001010001111" => data_out <= rom_array(29327);
		when "0111001010010000" => data_out <= rom_array(29328);
		when "0111001010010001" => data_out <= rom_array(29329);
		when "0111001010010010" => data_out <= rom_array(29330);
		when "0111001010010011" => data_out <= rom_array(29331);
		when "0111001010010100" => data_out <= rom_array(29332);
		when "0111001010010101" => data_out <= rom_array(29333);
		when "0111001010010110" => data_out <= rom_array(29334);
		when "0111001010010111" => data_out <= rom_array(29335);
		when "0111001010011000" => data_out <= rom_array(29336);
		when "0111001010011001" => data_out <= rom_array(29337);
		when "0111001010011010" => data_out <= rom_array(29338);
		when "0111001010011011" => data_out <= rom_array(29339);
		when "0111001010011100" => data_out <= rom_array(29340);
		when "0111001010011101" => data_out <= rom_array(29341);
		when "0111001010011110" => data_out <= rom_array(29342);
		when "0111001010011111" => data_out <= rom_array(29343);
		when "0111001010100000" => data_out <= rom_array(29344);
		when "0111001010100001" => data_out <= rom_array(29345);
		when "0111001010100010" => data_out <= rom_array(29346);
		when "0111001010100011" => data_out <= rom_array(29347);
		when "0111001010100100" => data_out <= rom_array(29348);
		when "0111001010100101" => data_out <= rom_array(29349);
		when "0111001010100110" => data_out <= rom_array(29350);
		when "0111001010100111" => data_out <= rom_array(29351);
		when "0111001010101000" => data_out <= rom_array(29352);
		when "0111001010101001" => data_out <= rom_array(29353);
		when "0111001010101010" => data_out <= rom_array(29354);
		when "0111001010101011" => data_out <= rom_array(29355);
		when "0111001010101100" => data_out <= rom_array(29356);
		when "0111001010101101" => data_out <= rom_array(29357);
		when "0111001010101110" => data_out <= rom_array(29358);
		when "0111001010101111" => data_out <= rom_array(29359);
		when "0111001010110000" => data_out <= rom_array(29360);
		when "0111001010110001" => data_out <= rom_array(29361);
		when "0111001010110010" => data_out <= rom_array(29362);
		when "0111001010110011" => data_out <= rom_array(29363);
		when "0111001010110100" => data_out <= rom_array(29364);
		when "0111001010110101" => data_out <= rom_array(29365);
		when "0111001010110110" => data_out <= rom_array(29366);
		when "0111001010110111" => data_out <= rom_array(29367);
		when "0111001010111000" => data_out <= rom_array(29368);
		when "0111001010111001" => data_out <= rom_array(29369);
		when "0111001010111010" => data_out <= rom_array(29370);
		when "0111001010111011" => data_out <= rom_array(29371);
		when "0111001010111100" => data_out <= rom_array(29372);
		when "0111001010111101" => data_out <= rom_array(29373);
		when "0111001010111110" => data_out <= rom_array(29374);
		when "0111001010111111" => data_out <= rom_array(29375);
		when "0111001011000000" => data_out <= rom_array(29376);
		when "0111001011000001" => data_out <= rom_array(29377);
		when "0111001011000010" => data_out <= rom_array(29378);
		when "0111001011000011" => data_out <= rom_array(29379);
		when "0111001011000100" => data_out <= rom_array(29380);
		when "0111001011000101" => data_out <= rom_array(29381);
		when "0111001011000110" => data_out <= rom_array(29382);
		when "0111001011000111" => data_out <= rom_array(29383);
		when "0111001011001000" => data_out <= rom_array(29384);
		when "0111001011001001" => data_out <= rom_array(29385);
		when "0111001011001010" => data_out <= rom_array(29386);
		when "0111001011001011" => data_out <= rom_array(29387);
		when "0111001011001100" => data_out <= rom_array(29388);
		when "0111001011001101" => data_out <= rom_array(29389);
		when "0111001011001110" => data_out <= rom_array(29390);
		when "0111001011001111" => data_out <= rom_array(29391);
		when "0111001011010000" => data_out <= rom_array(29392);
		when "0111001011010001" => data_out <= rom_array(29393);
		when "0111001011010010" => data_out <= rom_array(29394);
		when "0111001011010011" => data_out <= rom_array(29395);
		when "0111001011010100" => data_out <= rom_array(29396);
		when "0111001011010101" => data_out <= rom_array(29397);
		when "0111001011010110" => data_out <= rom_array(29398);
		when "0111001011010111" => data_out <= rom_array(29399);
		when "0111001011011000" => data_out <= rom_array(29400);
		when "0111001011011001" => data_out <= rom_array(29401);
		when "0111001011011010" => data_out <= rom_array(29402);
		when "0111001011011011" => data_out <= rom_array(29403);
		when "0111001011011100" => data_out <= rom_array(29404);
		when "0111001011011101" => data_out <= rom_array(29405);
		when "0111001011011110" => data_out <= rom_array(29406);
		when "0111001011011111" => data_out <= rom_array(29407);
		when "0111001011100000" => data_out <= rom_array(29408);
		when "0111001011100001" => data_out <= rom_array(29409);
		when "0111001011100010" => data_out <= rom_array(29410);
		when "0111001011100011" => data_out <= rom_array(29411);
		when "0111001011100100" => data_out <= rom_array(29412);
		when "0111001011100101" => data_out <= rom_array(29413);
		when "0111001011100110" => data_out <= rom_array(29414);
		when "0111001011100111" => data_out <= rom_array(29415);
		when "0111001011101000" => data_out <= rom_array(29416);
		when "0111001011101001" => data_out <= rom_array(29417);
		when "0111001011101010" => data_out <= rom_array(29418);
		when "0111001011101011" => data_out <= rom_array(29419);
		when "0111001011101100" => data_out <= rom_array(29420);
		when "0111001011101101" => data_out <= rom_array(29421);
		when "0111001011101110" => data_out <= rom_array(29422);
		when "0111001011101111" => data_out <= rom_array(29423);
		when "0111001011110000" => data_out <= rom_array(29424);
		when "0111001011110001" => data_out <= rom_array(29425);
		when "0111001011110010" => data_out <= rom_array(29426);
		when "0111001011110011" => data_out <= rom_array(29427);
		when "0111001011110100" => data_out <= rom_array(29428);
		when "0111001011110101" => data_out <= rom_array(29429);
		when "0111001011110110" => data_out <= rom_array(29430);
		when "0111001011110111" => data_out <= rom_array(29431);
		when "0111001011111000" => data_out <= rom_array(29432);
		when "0111001011111001" => data_out <= rom_array(29433);
		when "0111001011111010" => data_out <= rom_array(29434);
		when "0111001011111011" => data_out <= rom_array(29435);
		when "0111001011111100" => data_out <= rom_array(29436);
		when "0111001011111101" => data_out <= rom_array(29437);
		when "0111001011111110" => data_out <= rom_array(29438);
		when "0111001011111111" => data_out <= rom_array(29439);
		when "0111001100000000" => data_out <= rom_array(29440);
		when "0111001100000001" => data_out <= rom_array(29441);
		when "0111001100000010" => data_out <= rom_array(29442);
		when "0111001100000011" => data_out <= rom_array(29443);
		when "0111001100000100" => data_out <= rom_array(29444);
		when "0111001100000101" => data_out <= rom_array(29445);
		when "0111001100000110" => data_out <= rom_array(29446);
		when "0111001100000111" => data_out <= rom_array(29447);
		when "0111001100001000" => data_out <= rom_array(29448);
		when "0111001100001001" => data_out <= rom_array(29449);
		when "0111001100001010" => data_out <= rom_array(29450);
		when "0111001100001011" => data_out <= rom_array(29451);
		when "0111001100001100" => data_out <= rom_array(29452);
		when "0111001100001101" => data_out <= rom_array(29453);
		when "0111001100001110" => data_out <= rom_array(29454);
		when "0111001100001111" => data_out <= rom_array(29455);
		when "0111001100010000" => data_out <= rom_array(29456);
		when "0111001100010001" => data_out <= rom_array(29457);
		when "0111001100010010" => data_out <= rom_array(29458);
		when "0111001100010011" => data_out <= rom_array(29459);
		when "0111001100010100" => data_out <= rom_array(29460);
		when "0111001100010101" => data_out <= rom_array(29461);
		when "0111001100010110" => data_out <= rom_array(29462);
		when "0111001100010111" => data_out <= rom_array(29463);
		when "0111001100011000" => data_out <= rom_array(29464);
		when "0111001100011001" => data_out <= rom_array(29465);
		when "0111001100011010" => data_out <= rom_array(29466);
		when "0111001100011011" => data_out <= rom_array(29467);
		when "0111001100011100" => data_out <= rom_array(29468);
		when "0111001100011101" => data_out <= rom_array(29469);
		when "0111001100011110" => data_out <= rom_array(29470);
		when "0111001100011111" => data_out <= rom_array(29471);
		when "0111001100100000" => data_out <= rom_array(29472);
		when "0111001100100001" => data_out <= rom_array(29473);
		when "0111001100100010" => data_out <= rom_array(29474);
		when "0111001100100011" => data_out <= rom_array(29475);
		when "0111001100100100" => data_out <= rom_array(29476);
		when "0111001100100101" => data_out <= rom_array(29477);
		when "0111001100100110" => data_out <= rom_array(29478);
		when "0111001100100111" => data_out <= rom_array(29479);
		when "0111001100101000" => data_out <= rom_array(29480);
		when "0111001100101001" => data_out <= rom_array(29481);
		when "0111001100101010" => data_out <= rom_array(29482);
		when "0111001100101011" => data_out <= rom_array(29483);
		when "0111001100101100" => data_out <= rom_array(29484);
		when "0111001100101101" => data_out <= rom_array(29485);
		when "0111001100101110" => data_out <= rom_array(29486);
		when "0111001100101111" => data_out <= rom_array(29487);
		when "0111001100110000" => data_out <= rom_array(29488);
		when "0111001100110001" => data_out <= rom_array(29489);
		when "0111001100110010" => data_out <= rom_array(29490);
		when "0111001100110011" => data_out <= rom_array(29491);
		when "0111001100110100" => data_out <= rom_array(29492);
		when "0111001100110101" => data_out <= rom_array(29493);
		when "0111001100110110" => data_out <= rom_array(29494);
		when "0111001100110111" => data_out <= rom_array(29495);
		when "0111001100111000" => data_out <= rom_array(29496);
		when "0111001100111001" => data_out <= rom_array(29497);
		when "0111001100111010" => data_out <= rom_array(29498);
		when "0111001100111011" => data_out <= rom_array(29499);
		when "0111001100111100" => data_out <= rom_array(29500);
		when "0111001100111101" => data_out <= rom_array(29501);
		when "0111001100111110" => data_out <= rom_array(29502);
		when "0111001100111111" => data_out <= rom_array(29503);
		when "0111001101000000" => data_out <= rom_array(29504);
		when "0111001101000001" => data_out <= rom_array(29505);
		when "0111001101000010" => data_out <= rom_array(29506);
		when "0111001101000011" => data_out <= rom_array(29507);
		when "0111001101000100" => data_out <= rom_array(29508);
		when "0111001101000101" => data_out <= rom_array(29509);
		when "0111001101000110" => data_out <= rom_array(29510);
		when "0111001101000111" => data_out <= rom_array(29511);
		when "0111001101001000" => data_out <= rom_array(29512);
		when "0111001101001001" => data_out <= rom_array(29513);
		when "0111001101001010" => data_out <= rom_array(29514);
		when "0111001101001011" => data_out <= rom_array(29515);
		when "0111001101001100" => data_out <= rom_array(29516);
		when "0111001101001101" => data_out <= rom_array(29517);
		when "0111001101001110" => data_out <= rom_array(29518);
		when "0111001101001111" => data_out <= rom_array(29519);
		when "0111001101010000" => data_out <= rom_array(29520);
		when "0111001101010001" => data_out <= rom_array(29521);
		when "0111001101010010" => data_out <= rom_array(29522);
		when "0111001101010011" => data_out <= rom_array(29523);
		when "0111001101010100" => data_out <= rom_array(29524);
		when "0111001101010101" => data_out <= rom_array(29525);
		when "0111001101010110" => data_out <= rom_array(29526);
		when "0111001101010111" => data_out <= rom_array(29527);
		when "0111001101011000" => data_out <= rom_array(29528);
		when "0111001101011001" => data_out <= rom_array(29529);
		when "0111001101011010" => data_out <= rom_array(29530);
		when "0111001101011011" => data_out <= rom_array(29531);
		when "0111001101011100" => data_out <= rom_array(29532);
		when "0111001101011101" => data_out <= rom_array(29533);
		when "0111001101011110" => data_out <= rom_array(29534);
		when "0111001101011111" => data_out <= rom_array(29535);
		when "0111001101100000" => data_out <= rom_array(29536);
		when "0111001101100001" => data_out <= rom_array(29537);
		when "0111001101100010" => data_out <= rom_array(29538);
		when "0111001101100011" => data_out <= rom_array(29539);
		when "0111001101100100" => data_out <= rom_array(29540);
		when "0111001101100101" => data_out <= rom_array(29541);
		when "0111001101100110" => data_out <= rom_array(29542);
		when "0111001101100111" => data_out <= rom_array(29543);
		when "0111001101101000" => data_out <= rom_array(29544);
		when "0111001101101001" => data_out <= rom_array(29545);
		when "0111001101101010" => data_out <= rom_array(29546);
		when "0111001101101011" => data_out <= rom_array(29547);
		when "0111001101101100" => data_out <= rom_array(29548);
		when "0111001101101101" => data_out <= rom_array(29549);
		when "0111001101101110" => data_out <= rom_array(29550);
		when "0111001101101111" => data_out <= rom_array(29551);
		when "0111001101110000" => data_out <= rom_array(29552);
		when "0111001101110001" => data_out <= rom_array(29553);
		when "0111001101110010" => data_out <= rom_array(29554);
		when "0111001101110011" => data_out <= rom_array(29555);
		when "0111001101110100" => data_out <= rom_array(29556);
		when "0111001101110101" => data_out <= rom_array(29557);
		when "0111001101110110" => data_out <= rom_array(29558);
		when "0111001101110111" => data_out <= rom_array(29559);
		when "0111001101111000" => data_out <= rom_array(29560);
		when "0111001101111001" => data_out <= rom_array(29561);
		when "0111001101111010" => data_out <= rom_array(29562);
		when "0111001101111011" => data_out <= rom_array(29563);
		when "0111001101111100" => data_out <= rom_array(29564);
		when "0111001101111101" => data_out <= rom_array(29565);
		when "0111001101111110" => data_out <= rom_array(29566);
		when "0111001101111111" => data_out <= rom_array(29567);
		when "0111001110000000" => data_out <= rom_array(29568);
		when "0111001110000001" => data_out <= rom_array(29569);
		when "0111001110000010" => data_out <= rom_array(29570);
		when "0111001110000011" => data_out <= rom_array(29571);
		when "0111001110000100" => data_out <= rom_array(29572);
		when "0111001110000101" => data_out <= rom_array(29573);
		when "0111001110000110" => data_out <= rom_array(29574);
		when "0111001110000111" => data_out <= rom_array(29575);
		when "0111001110001000" => data_out <= rom_array(29576);
		when "0111001110001001" => data_out <= rom_array(29577);
		when "0111001110001010" => data_out <= rom_array(29578);
		when "0111001110001011" => data_out <= rom_array(29579);
		when "0111001110001100" => data_out <= rom_array(29580);
		when "0111001110001101" => data_out <= rom_array(29581);
		when "0111001110001110" => data_out <= rom_array(29582);
		when "0111001110001111" => data_out <= rom_array(29583);
		when "0111001110010000" => data_out <= rom_array(29584);
		when "0111001110010001" => data_out <= rom_array(29585);
		when "0111001110010010" => data_out <= rom_array(29586);
		when "0111001110010011" => data_out <= rom_array(29587);
		when "0111001110010100" => data_out <= rom_array(29588);
		when "0111001110010101" => data_out <= rom_array(29589);
		when "0111001110010110" => data_out <= rom_array(29590);
		when "0111001110010111" => data_out <= rom_array(29591);
		when "0111001110011000" => data_out <= rom_array(29592);
		when "0111001110011001" => data_out <= rom_array(29593);
		when "0111001110011010" => data_out <= rom_array(29594);
		when "0111001110011011" => data_out <= rom_array(29595);
		when "0111001110011100" => data_out <= rom_array(29596);
		when "0111001110011101" => data_out <= rom_array(29597);
		when "0111001110011110" => data_out <= rom_array(29598);
		when "0111001110011111" => data_out <= rom_array(29599);
		when "0111001110100000" => data_out <= rom_array(29600);
		when "0111001110100001" => data_out <= rom_array(29601);
		when "0111001110100010" => data_out <= rom_array(29602);
		when "0111001110100011" => data_out <= rom_array(29603);
		when "0111001110100100" => data_out <= rom_array(29604);
		when "0111001110100101" => data_out <= rom_array(29605);
		when "0111001110100110" => data_out <= rom_array(29606);
		when "0111001110100111" => data_out <= rom_array(29607);
		when "0111001110101000" => data_out <= rom_array(29608);
		when "0111001110101001" => data_out <= rom_array(29609);
		when "0111001110101010" => data_out <= rom_array(29610);
		when "0111001110101011" => data_out <= rom_array(29611);
		when "0111001110101100" => data_out <= rom_array(29612);
		when "0111001110101101" => data_out <= rom_array(29613);
		when "0111001110101110" => data_out <= rom_array(29614);
		when "0111001110101111" => data_out <= rom_array(29615);
		when "0111001110110000" => data_out <= rom_array(29616);
		when "0111001110110001" => data_out <= rom_array(29617);
		when "0111001110110010" => data_out <= rom_array(29618);
		when "0111001110110011" => data_out <= rom_array(29619);
		when "0111001110110100" => data_out <= rom_array(29620);
		when "0111001110110101" => data_out <= rom_array(29621);
		when "0111001110110110" => data_out <= rom_array(29622);
		when "0111001110110111" => data_out <= rom_array(29623);
		when "0111001110111000" => data_out <= rom_array(29624);
		when "0111001110111001" => data_out <= rom_array(29625);
		when "0111001110111010" => data_out <= rom_array(29626);
		when "0111001110111011" => data_out <= rom_array(29627);
		when "0111001110111100" => data_out <= rom_array(29628);
		when "0111001110111101" => data_out <= rom_array(29629);
		when "0111001110111110" => data_out <= rom_array(29630);
		when "0111001110111111" => data_out <= rom_array(29631);
		when "0111001111000000" => data_out <= rom_array(29632);
		when "0111001111000001" => data_out <= rom_array(29633);
		when "0111001111000010" => data_out <= rom_array(29634);
		when "0111001111000011" => data_out <= rom_array(29635);
		when "0111001111000100" => data_out <= rom_array(29636);
		when "0111001111000101" => data_out <= rom_array(29637);
		when "0111001111000110" => data_out <= rom_array(29638);
		when "0111001111000111" => data_out <= rom_array(29639);
		when "0111001111001000" => data_out <= rom_array(29640);
		when "0111001111001001" => data_out <= rom_array(29641);
		when "0111001111001010" => data_out <= rom_array(29642);
		when "0111001111001011" => data_out <= rom_array(29643);
		when "0111001111001100" => data_out <= rom_array(29644);
		when "0111001111001101" => data_out <= rom_array(29645);
		when "0111001111001110" => data_out <= rom_array(29646);
		when "0111001111001111" => data_out <= rom_array(29647);
		when "0111001111010000" => data_out <= rom_array(29648);
		when "0111001111010001" => data_out <= rom_array(29649);
		when "0111001111010010" => data_out <= rom_array(29650);
		when "0111001111010011" => data_out <= rom_array(29651);
		when "0111001111010100" => data_out <= rom_array(29652);
		when "0111001111010101" => data_out <= rom_array(29653);
		when "0111001111010110" => data_out <= rom_array(29654);
		when "0111001111010111" => data_out <= rom_array(29655);
		when "0111001111011000" => data_out <= rom_array(29656);
		when "0111001111011001" => data_out <= rom_array(29657);
		when "0111001111011010" => data_out <= rom_array(29658);
		when "0111001111011011" => data_out <= rom_array(29659);
		when "0111001111011100" => data_out <= rom_array(29660);
		when "0111001111011101" => data_out <= rom_array(29661);
		when "0111001111011110" => data_out <= rom_array(29662);
		when "0111001111011111" => data_out <= rom_array(29663);
		when "0111001111100000" => data_out <= rom_array(29664);
		when "0111001111100001" => data_out <= rom_array(29665);
		when "0111001111100010" => data_out <= rom_array(29666);
		when "0111001111100011" => data_out <= rom_array(29667);
		when "0111001111100100" => data_out <= rom_array(29668);
		when "0111001111100101" => data_out <= rom_array(29669);
		when "0111001111100110" => data_out <= rom_array(29670);
		when "0111001111100111" => data_out <= rom_array(29671);
		when "0111001111101000" => data_out <= rom_array(29672);
		when "0111001111101001" => data_out <= rom_array(29673);
		when "0111001111101010" => data_out <= rom_array(29674);
		when "0111001111101011" => data_out <= rom_array(29675);
		when "0111001111101100" => data_out <= rom_array(29676);
		when "0111001111101101" => data_out <= rom_array(29677);
		when "0111001111101110" => data_out <= rom_array(29678);
		when "0111001111101111" => data_out <= rom_array(29679);
		when "0111001111110000" => data_out <= rom_array(29680);
		when "0111001111110001" => data_out <= rom_array(29681);
		when "0111001111110010" => data_out <= rom_array(29682);
		when "0111001111110011" => data_out <= rom_array(29683);
		when "0111001111110100" => data_out <= rom_array(29684);
		when "0111001111110101" => data_out <= rom_array(29685);
		when "0111001111110110" => data_out <= rom_array(29686);
		when "0111001111110111" => data_out <= rom_array(29687);
		when "0111001111111000" => data_out <= rom_array(29688);
		when "0111001111111001" => data_out <= rom_array(29689);
		when "0111001111111010" => data_out <= rom_array(29690);
		when "0111001111111011" => data_out <= rom_array(29691);
		when "0111001111111100" => data_out <= rom_array(29692);
		when "0111001111111101" => data_out <= rom_array(29693);
		when "0111001111111110" => data_out <= rom_array(29694);
		when "0111001111111111" => data_out <= rom_array(29695);
		when "0111010000000000" => data_out <= rom_array(29696);
		when "0111010000000001" => data_out <= rom_array(29697);
		when "0111010000000010" => data_out <= rom_array(29698);
		when "0111010000000011" => data_out <= rom_array(29699);
		when "0111010000000100" => data_out <= rom_array(29700);
		when "0111010000000101" => data_out <= rom_array(29701);
		when "0111010000000110" => data_out <= rom_array(29702);
		when "0111010000000111" => data_out <= rom_array(29703);
		when "0111010000001000" => data_out <= rom_array(29704);
		when "0111010000001001" => data_out <= rom_array(29705);
		when "0111010000001010" => data_out <= rom_array(29706);
		when "0111010000001011" => data_out <= rom_array(29707);
		when "0111010000001100" => data_out <= rom_array(29708);
		when "0111010000001101" => data_out <= rom_array(29709);
		when "0111010000001110" => data_out <= rom_array(29710);
		when "0111010000001111" => data_out <= rom_array(29711);
		when "0111010000010000" => data_out <= rom_array(29712);
		when "0111010000010001" => data_out <= rom_array(29713);
		when "0111010000010010" => data_out <= rom_array(29714);
		when "0111010000010011" => data_out <= rom_array(29715);
		when "0111010000010100" => data_out <= rom_array(29716);
		when "0111010000010101" => data_out <= rom_array(29717);
		when "0111010000010110" => data_out <= rom_array(29718);
		when "0111010000010111" => data_out <= rom_array(29719);
		when "0111010000011000" => data_out <= rom_array(29720);
		when "0111010000011001" => data_out <= rom_array(29721);
		when "0111010000011010" => data_out <= rom_array(29722);
		when "0111010000011011" => data_out <= rom_array(29723);
		when "0111010000011100" => data_out <= rom_array(29724);
		when "0111010000011101" => data_out <= rom_array(29725);
		when "0111010000011110" => data_out <= rom_array(29726);
		when "0111010000011111" => data_out <= rom_array(29727);
		when "0111010000100000" => data_out <= rom_array(29728);
		when "0111010000100001" => data_out <= rom_array(29729);
		when "0111010000100010" => data_out <= rom_array(29730);
		when "0111010000100011" => data_out <= rom_array(29731);
		when "0111010000100100" => data_out <= rom_array(29732);
		when "0111010000100101" => data_out <= rom_array(29733);
		when "0111010000100110" => data_out <= rom_array(29734);
		when "0111010000100111" => data_out <= rom_array(29735);
		when "0111010000101000" => data_out <= rom_array(29736);
		when "0111010000101001" => data_out <= rom_array(29737);
		when "0111010000101010" => data_out <= rom_array(29738);
		when "0111010000101011" => data_out <= rom_array(29739);
		when "0111010000101100" => data_out <= rom_array(29740);
		when "0111010000101101" => data_out <= rom_array(29741);
		when "0111010000101110" => data_out <= rom_array(29742);
		when "0111010000101111" => data_out <= rom_array(29743);
		when "0111010000110000" => data_out <= rom_array(29744);
		when "0111010000110001" => data_out <= rom_array(29745);
		when "0111010000110010" => data_out <= rom_array(29746);
		when "0111010000110011" => data_out <= rom_array(29747);
		when "0111010000110100" => data_out <= rom_array(29748);
		when "0111010000110101" => data_out <= rom_array(29749);
		when "0111010000110110" => data_out <= rom_array(29750);
		when "0111010000110111" => data_out <= rom_array(29751);
		when "0111010000111000" => data_out <= rom_array(29752);
		when "0111010000111001" => data_out <= rom_array(29753);
		when "0111010000111010" => data_out <= rom_array(29754);
		when "0111010000111011" => data_out <= rom_array(29755);
		when "0111010000111100" => data_out <= rom_array(29756);
		when "0111010000111101" => data_out <= rom_array(29757);
		when "0111010000111110" => data_out <= rom_array(29758);
		when "0111010000111111" => data_out <= rom_array(29759);
		when "0111010001000000" => data_out <= rom_array(29760);
		when "0111010001000001" => data_out <= rom_array(29761);
		when "0111010001000010" => data_out <= rom_array(29762);
		when "0111010001000011" => data_out <= rom_array(29763);
		when "0111010001000100" => data_out <= rom_array(29764);
		when "0111010001000101" => data_out <= rom_array(29765);
		when "0111010001000110" => data_out <= rom_array(29766);
		when "0111010001000111" => data_out <= rom_array(29767);
		when "0111010001001000" => data_out <= rom_array(29768);
		when "0111010001001001" => data_out <= rom_array(29769);
		when "0111010001001010" => data_out <= rom_array(29770);
		when "0111010001001011" => data_out <= rom_array(29771);
		when "0111010001001100" => data_out <= rom_array(29772);
		when "0111010001001101" => data_out <= rom_array(29773);
		when "0111010001001110" => data_out <= rom_array(29774);
		when "0111010001001111" => data_out <= rom_array(29775);
		when "0111010001010000" => data_out <= rom_array(29776);
		when "0111010001010001" => data_out <= rom_array(29777);
		when "0111010001010010" => data_out <= rom_array(29778);
		when "0111010001010011" => data_out <= rom_array(29779);
		when "0111010001010100" => data_out <= rom_array(29780);
		when "0111010001010101" => data_out <= rom_array(29781);
		when "0111010001010110" => data_out <= rom_array(29782);
		when "0111010001010111" => data_out <= rom_array(29783);
		when "0111010001011000" => data_out <= rom_array(29784);
		when "0111010001011001" => data_out <= rom_array(29785);
		when "0111010001011010" => data_out <= rom_array(29786);
		when "0111010001011011" => data_out <= rom_array(29787);
		when "0111010001011100" => data_out <= rom_array(29788);
		when "0111010001011101" => data_out <= rom_array(29789);
		when "0111010001011110" => data_out <= rom_array(29790);
		when "0111010001011111" => data_out <= rom_array(29791);
		when "0111010001100000" => data_out <= rom_array(29792);
		when "0111010001100001" => data_out <= rom_array(29793);
		when "0111010001100010" => data_out <= rom_array(29794);
		when "0111010001100011" => data_out <= rom_array(29795);
		when "0111010001100100" => data_out <= rom_array(29796);
		when "0111010001100101" => data_out <= rom_array(29797);
		when "0111010001100110" => data_out <= rom_array(29798);
		when "0111010001100111" => data_out <= rom_array(29799);
		when "0111010001101000" => data_out <= rom_array(29800);
		when "0111010001101001" => data_out <= rom_array(29801);
		when "0111010001101010" => data_out <= rom_array(29802);
		when "0111010001101011" => data_out <= rom_array(29803);
		when "0111010001101100" => data_out <= rom_array(29804);
		when "0111010001101101" => data_out <= rom_array(29805);
		when "0111010001101110" => data_out <= rom_array(29806);
		when "0111010001101111" => data_out <= rom_array(29807);
		when "0111010001110000" => data_out <= rom_array(29808);
		when "0111010001110001" => data_out <= rom_array(29809);
		when "0111010001110010" => data_out <= rom_array(29810);
		when "0111010001110011" => data_out <= rom_array(29811);
		when "0111010001110100" => data_out <= rom_array(29812);
		when "0111010001110101" => data_out <= rom_array(29813);
		when "0111010001110110" => data_out <= rom_array(29814);
		when "0111010001110111" => data_out <= rom_array(29815);
		when "0111010001111000" => data_out <= rom_array(29816);
		when "0111010001111001" => data_out <= rom_array(29817);
		when "0111010001111010" => data_out <= rom_array(29818);
		when "0111010001111011" => data_out <= rom_array(29819);
		when "0111010001111100" => data_out <= rom_array(29820);
		when "0111010001111101" => data_out <= rom_array(29821);
		when "0111010001111110" => data_out <= rom_array(29822);
		when "0111010001111111" => data_out <= rom_array(29823);
		when "0111010010000000" => data_out <= rom_array(29824);
		when "0111010010000001" => data_out <= rom_array(29825);
		when "0111010010000010" => data_out <= rom_array(29826);
		when "0111010010000011" => data_out <= rom_array(29827);
		when "0111010010000100" => data_out <= rom_array(29828);
		when "0111010010000101" => data_out <= rom_array(29829);
		when "0111010010000110" => data_out <= rom_array(29830);
		when "0111010010000111" => data_out <= rom_array(29831);
		when "0111010010001000" => data_out <= rom_array(29832);
		when "0111010010001001" => data_out <= rom_array(29833);
		when "0111010010001010" => data_out <= rom_array(29834);
		when "0111010010001011" => data_out <= rom_array(29835);
		when "0111010010001100" => data_out <= rom_array(29836);
		when "0111010010001101" => data_out <= rom_array(29837);
		when "0111010010001110" => data_out <= rom_array(29838);
		when "0111010010001111" => data_out <= rom_array(29839);
		when "0111010010010000" => data_out <= rom_array(29840);
		when "0111010010010001" => data_out <= rom_array(29841);
		when "0111010010010010" => data_out <= rom_array(29842);
		when "0111010010010011" => data_out <= rom_array(29843);
		when "0111010010010100" => data_out <= rom_array(29844);
		when "0111010010010101" => data_out <= rom_array(29845);
		when "0111010010010110" => data_out <= rom_array(29846);
		when "0111010010010111" => data_out <= rom_array(29847);
		when "0111010010011000" => data_out <= rom_array(29848);
		when "0111010010011001" => data_out <= rom_array(29849);
		when "0111010010011010" => data_out <= rom_array(29850);
		when "0111010010011011" => data_out <= rom_array(29851);
		when "0111010010011100" => data_out <= rom_array(29852);
		when "0111010010011101" => data_out <= rom_array(29853);
		when "0111010010011110" => data_out <= rom_array(29854);
		when "0111010010011111" => data_out <= rom_array(29855);
		when "0111010010100000" => data_out <= rom_array(29856);
		when "0111010010100001" => data_out <= rom_array(29857);
		when "0111010010100010" => data_out <= rom_array(29858);
		when "0111010010100011" => data_out <= rom_array(29859);
		when "0111010010100100" => data_out <= rom_array(29860);
		when "0111010010100101" => data_out <= rom_array(29861);
		when "0111010010100110" => data_out <= rom_array(29862);
		when "0111010010100111" => data_out <= rom_array(29863);
		when "0111010010101000" => data_out <= rom_array(29864);
		when "0111010010101001" => data_out <= rom_array(29865);
		when "0111010010101010" => data_out <= rom_array(29866);
		when "0111010010101011" => data_out <= rom_array(29867);
		when "0111010010101100" => data_out <= rom_array(29868);
		when "0111010010101101" => data_out <= rom_array(29869);
		when "0111010010101110" => data_out <= rom_array(29870);
		when "0111010010101111" => data_out <= rom_array(29871);
		when "0111010010110000" => data_out <= rom_array(29872);
		when "0111010010110001" => data_out <= rom_array(29873);
		when "0111010010110010" => data_out <= rom_array(29874);
		when "0111010010110011" => data_out <= rom_array(29875);
		when "0111010010110100" => data_out <= rom_array(29876);
		when "0111010010110101" => data_out <= rom_array(29877);
		when "0111010010110110" => data_out <= rom_array(29878);
		when "0111010010110111" => data_out <= rom_array(29879);
		when "0111010010111000" => data_out <= rom_array(29880);
		when "0111010010111001" => data_out <= rom_array(29881);
		when "0111010010111010" => data_out <= rom_array(29882);
		when "0111010010111011" => data_out <= rom_array(29883);
		when "0111010010111100" => data_out <= rom_array(29884);
		when "0111010010111101" => data_out <= rom_array(29885);
		when "0111010010111110" => data_out <= rom_array(29886);
		when "0111010010111111" => data_out <= rom_array(29887);
		when "0111010011000000" => data_out <= rom_array(29888);
		when "0111010011000001" => data_out <= rom_array(29889);
		when "0111010011000010" => data_out <= rom_array(29890);
		when "0111010011000011" => data_out <= rom_array(29891);
		when "0111010011000100" => data_out <= rom_array(29892);
		when "0111010011000101" => data_out <= rom_array(29893);
		when "0111010011000110" => data_out <= rom_array(29894);
		when "0111010011000111" => data_out <= rom_array(29895);
		when "0111010011001000" => data_out <= rom_array(29896);
		when "0111010011001001" => data_out <= rom_array(29897);
		when "0111010011001010" => data_out <= rom_array(29898);
		when "0111010011001011" => data_out <= rom_array(29899);
		when "0111010011001100" => data_out <= rom_array(29900);
		when "0111010011001101" => data_out <= rom_array(29901);
		when "0111010011001110" => data_out <= rom_array(29902);
		when "0111010011001111" => data_out <= rom_array(29903);
		when "0111010011010000" => data_out <= rom_array(29904);
		when "0111010011010001" => data_out <= rom_array(29905);
		when "0111010011010010" => data_out <= rom_array(29906);
		when "0111010011010011" => data_out <= rom_array(29907);
		when "0111010011010100" => data_out <= rom_array(29908);
		when "0111010011010101" => data_out <= rom_array(29909);
		when "0111010011010110" => data_out <= rom_array(29910);
		when "0111010011010111" => data_out <= rom_array(29911);
		when "0111010011011000" => data_out <= rom_array(29912);
		when "0111010011011001" => data_out <= rom_array(29913);
		when "0111010011011010" => data_out <= rom_array(29914);
		when "0111010011011011" => data_out <= rom_array(29915);
		when "0111010011011100" => data_out <= rom_array(29916);
		when "0111010011011101" => data_out <= rom_array(29917);
		when "0111010011011110" => data_out <= rom_array(29918);
		when "0111010011011111" => data_out <= rom_array(29919);
		when "0111010011100000" => data_out <= rom_array(29920);
		when "0111010011100001" => data_out <= rom_array(29921);
		when "0111010011100010" => data_out <= rom_array(29922);
		when "0111010011100011" => data_out <= rom_array(29923);
		when "0111010011100100" => data_out <= rom_array(29924);
		when "0111010011100101" => data_out <= rom_array(29925);
		when "0111010011100110" => data_out <= rom_array(29926);
		when "0111010011100111" => data_out <= rom_array(29927);
		when "0111010011101000" => data_out <= rom_array(29928);
		when "0111010011101001" => data_out <= rom_array(29929);
		when "0111010011101010" => data_out <= rom_array(29930);
		when "0111010011101011" => data_out <= rom_array(29931);
		when "0111010011101100" => data_out <= rom_array(29932);
		when "0111010011101101" => data_out <= rom_array(29933);
		when "0111010011101110" => data_out <= rom_array(29934);
		when "0111010011101111" => data_out <= rom_array(29935);
		when "0111010011110000" => data_out <= rom_array(29936);
		when "0111010011110001" => data_out <= rom_array(29937);
		when "0111010011110010" => data_out <= rom_array(29938);
		when "0111010011110011" => data_out <= rom_array(29939);
		when "0111010011110100" => data_out <= rom_array(29940);
		when "0111010011110101" => data_out <= rom_array(29941);
		when "0111010011110110" => data_out <= rom_array(29942);
		when "0111010011110111" => data_out <= rom_array(29943);
		when "0111010011111000" => data_out <= rom_array(29944);
		when "0111010011111001" => data_out <= rom_array(29945);
		when "0111010011111010" => data_out <= rom_array(29946);
		when "0111010011111011" => data_out <= rom_array(29947);
		when "0111010011111100" => data_out <= rom_array(29948);
		when "0111010011111101" => data_out <= rom_array(29949);
		when "0111010011111110" => data_out <= rom_array(29950);
		when "0111010011111111" => data_out <= rom_array(29951);
		when "0111010100000000" => data_out <= rom_array(29952);
		when "0111010100000001" => data_out <= rom_array(29953);
		when "0111010100000010" => data_out <= rom_array(29954);
		when "0111010100000011" => data_out <= rom_array(29955);
		when "0111010100000100" => data_out <= rom_array(29956);
		when "0111010100000101" => data_out <= rom_array(29957);
		when "0111010100000110" => data_out <= rom_array(29958);
		when "0111010100000111" => data_out <= rom_array(29959);
		when "0111010100001000" => data_out <= rom_array(29960);
		when "0111010100001001" => data_out <= rom_array(29961);
		when "0111010100001010" => data_out <= rom_array(29962);
		when "0111010100001011" => data_out <= rom_array(29963);
		when "0111010100001100" => data_out <= rom_array(29964);
		when "0111010100001101" => data_out <= rom_array(29965);
		when "0111010100001110" => data_out <= rom_array(29966);
		when "0111010100001111" => data_out <= rom_array(29967);
		when "0111010100010000" => data_out <= rom_array(29968);
		when "0111010100010001" => data_out <= rom_array(29969);
		when "0111010100010010" => data_out <= rom_array(29970);
		when "0111010100010011" => data_out <= rom_array(29971);
		when "0111010100010100" => data_out <= rom_array(29972);
		when "0111010100010101" => data_out <= rom_array(29973);
		when "0111010100010110" => data_out <= rom_array(29974);
		when "0111010100010111" => data_out <= rom_array(29975);
		when "0111010100011000" => data_out <= rom_array(29976);
		when "0111010100011001" => data_out <= rom_array(29977);
		when "0111010100011010" => data_out <= rom_array(29978);
		when "0111010100011011" => data_out <= rom_array(29979);
		when "0111010100011100" => data_out <= rom_array(29980);
		when "0111010100011101" => data_out <= rom_array(29981);
		when "0111010100011110" => data_out <= rom_array(29982);
		when "0111010100011111" => data_out <= rom_array(29983);
		when "0111010100100000" => data_out <= rom_array(29984);
		when "0111010100100001" => data_out <= rom_array(29985);
		when "0111010100100010" => data_out <= rom_array(29986);
		when "0111010100100011" => data_out <= rom_array(29987);
		when "0111010100100100" => data_out <= rom_array(29988);
		when "0111010100100101" => data_out <= rom_array(29989);
		when "0111010100100110" => data_out <= rom_array(29990);
		when "0111010100100111" => data_out <= rom_array(29991);
		when "0111010100101000" => data_out <= rom_array(29992);
		when "0111010100101001" => data_out <= rom_array(29993);
		when "0111010100101010" => data_out <= rom_array(29994);
		when "0111010100101011" => data_out <= rom_array(29995);
		when "0111010100101100" => data_out <= rom_array(29996);
		when "0111010100101101" => data_out <= rom_array(29997);
		when "0111010100101110" => data_out <= rom_array(29998);
		when "0111010100101111" => data_out <= rom_array(29999);
		when "0111010100110000" => data_out <= rom_array(30000);
		when "0111010100110001" => data_out <= rom_array(30001);
		when "0111010100110010" => data_out <= rom_array(30002);
		when "0111010100110011" => data_out <= rom_array(30003);
		when "0111010100110100" => data_out <= rom_array(30004);
		when "0111010100110101" => data_out <= rom_array(30005);
		when "0111010100110110" => data_out <= rom_array(30006);
		when "0111010100110111" => data_out <= rom_array(30007);
		when "0111010100111000" => data_out <= rom_array(30008);
		when "0111010100111001" => data_out <= rom_array(30009);
		when "0111010100111010" => data_out <= rom_array(30010);
		when "0111010100111011" => data_out <= rom_array(30011);
		when "0111010100111100" => data_out <= rom_array(30012);
		when "0111010100111101" => data_out <= rom_array(30013);
		when "0111010100111110" => data_out <= rom_array(30014);
		when "0111010100111111" => data_out <= rom_array(30015);
		when "0111010101000000" => data_out <= rom_array(30016);
		when "0111010101000001" => data_out <= rom_array(30017);
		when "0111010101000010" => data_out <= rom_array(30018);
		when "0111010101000011" => data_out <= rom_array(30019);
		when "0111010101000100" => data_out <= rom_array(30020);
		when "0111010101000101" => data_out <= rom_array(30021);
		when "0111010101000110" => data_out <= rom_array(30022);
		when "0111010101000111" => data_out <= rom_array(30023);
		when "0111010101001000" => data_out <= rom_array(30024);
		when "0111010101001001" => data_out <= rom_array(30025);
		when "0111010101001010" => data_out <= rom_array(30026);
		when "0111010101001011" => data_out <= rom_array(30027);
		when "0111010101001100" => data_out <= rom_array(30028);
		when "0111010101001101" => data_out <= rom_array(30029);
		when "0111010101001110" => data_out <= rom_array(30030);
		when "0111010101001111" => data_out <= rom_array(30031);
		when "0111010101010000" => data_out <= rom_array(30032);
		when "0111010101010001" => data_out <= rom_array(30033);
		when "0111010101010010" => data_out <= rom_array(30034);
		when "0111010101010011" => data_out <= rom_array(30035);
		when "0111010101010100" => data_out <= rom_array(30036);
		when "0111010101010101" => data_out <= rom_array(30037);
		when "0111010101010110" => data_out <= rom_array(30038);
		when "0111010101010111" => data_out <= rom_array(30039);
		when "0111010101011000" => data_out <= rom_array(30040);
		when "0111010101011001" => data_out <= rom_array(30041);
		when "0111010101011010" => data_out <= rom_array(30042);
		when "0111010101011011" => data_out <= rom_array(30043);
		when "0111010101011100" => data_out <= rom_array(30044);
		when "0111010101011101" => data_out <= rom_array(30045);
		when "0111010101011110" => data_out <= rom_array(30046);
		when "0111010101011111" => data_out <= rom_array(30047);
		when "0111010101100000" => data_out <= rom_array(30048);
		when "0111010101100001" => data_out <= rom_array(30049);
		when "0111010101100010" => data_out <= rom_array(30050);
		when "0111010101100011" => data_out <= rom_array(30051);
		when "0111010101100100" => data_out <= rom_array(30052);
		when "0111010101100101" => data_out <= rom_array(30053);
		when "0111010101100110" => data_out <= rom_array(30054);
		when "0111010101100111" => data_out <= rom_array(30055);
		when "0111010101101000" => data_out <= rom_array(30056);
		when "0111010101101001" => data_out <= rom_array(30057);
		when "0111010101101010" => data_out <= rom_array(30058);
		when "0111010101101011" => data_out <= rom_array(30059);
		when "0111010101101100" => data_out <= rom_array(30060);
		when "0111010101101101" => data_out <= rom_array(30061);
		when "0111010101101110" => data_out <= rom_array(30062);
		when "0111010101101111" => data_out <= rom_array(30063);
		when "0111010101110000" => data_out <= rom_array(30064);
		when "0111010101110001" => data_out <= rom_array(30065);
		when "0111010101110010" => data_out <= rom_array(30066);
		when "0111010101110011" => data_out <= rom_array(30067);
		when "0111010101110100" => data_out <= rom_array(30068);
		when "0111010101110101" => data_out <= rom_array(30069);
		when "0111010101110110" => data_out <= rom_array(30070);
		when "0111010101110111" => data_out <= rom_array(30071);
		when "0111010101111000" => data_out <= rom_array(30072);
		when "0111010101111001" => data_out <= rom_array(30073);
		when "0111010101111010" => data_out <= rom_array(30074);
		when "0111010101111011" => data_out <= rom_array(30075);
		when "0111010101111100" => data_out <= rom_array(30076);
		when "0111010101111101" => data_out <= rom_array(30077);
		when "0111010101111110" => data_out <= rom_array(30078);
		when "0111010101111111" => data_out <= rom_array(30079);
		when "0111010110000000" => data_out <= rom_array(30080);
		when "0111010110000001" => data_out <= rom_array(30081);
		when "0111010110000010" => data_out <= rom_array(30082);
		when "0111010110000011" => data_out <= rom_array(30083);
		when "0111010110000100" => data_out <= rom_array(30084);
		when "0111010110000101" => data_out <= rom_array(30085);
		when "0111010110000110" => data_out <= rom_array(30086);
		when "0111010110000111" => data_out <= rom_array(30087);
		when "0111010110001000" => data_out <= rom_array(30088);
		when "0111010110001001" => data_out <= rom_array(30089);
		when "0111010110001010" => data_out <= rom_array(30090);
		when "0111010110001011" => data_out <= rom_array(30091);
		when "0111010110001100" => data_out <= rom_array(30092);
		when "0111010110001101" => data_out <= rom_array(30093);
		when "0111010110001110" => data_out <= rom_array(30094);
		when "0111010110001111" => data_out <= rom_array(30095);
		when "0111010110010000" => data_out <= rom_array(30096);
		when "0111010110010001" => data_out <= rom_array(30097);
		when "0111010110010010" => data_out <= rom_array(30098);
		when "0111010110010011" => data_out <= rom_array(30099);
		when "0111010110010100" => data_out <= rom_array(30100);
		when "0111010110010101" => data_out <= rom_array(30101);
		when "0111010110010110" => data_out <= rom_array(30102);
		when "0111010110010111" => data_out <= rom_array(30103);
		when "0111010110011000" => data_out <= rom_array(30104);
		when "0111010110011001" => data_out <= rom_array(30105);
		when "0111010110011010" => data_out <= rom_array(30106);
		when "0111010110011011" => data_out <= rom_array(30107);
		when "0111010110011100" => data_out <= rom_array(30108);
		when "0111010110011101" => data_out <= rom_array(30109);
		when "0111010110011110" => data_out <= rom_array(30110);
		when "0111010110011111" => data_out <= rom_array(30111);
		when "0111010110100000" => data_out <= rom_array(30112);
		when "0111010110100001" => data_out <= rom_array(30113);
		when "0111010110100010" => data_out <= rom_array(30114);
		when "0111010110100011" => data_out <= rom_array(30115);
		when "0111010110100100" => data_out <= rom_array(30116);
		when "0111010110100101" => data_out <= rom_array(30117);
		when "0111010110100110" => data_out <= rom_array(30118);
		when "0111010110100111" => data_out <= rom_array(30119);
		when "0111010110101000" => data_out <= rom_array(30120);
		when "0111010110101001" => data_out <= rom_array(30121);
		when "0111010110101010" => data_out <= rom_array(30122);
		when "0111010110101011" => data_out <= rom_array(30123);
		when "0111010110101100" => data_out <= rom_array(30124);
		when "0111010110101101" => data_out <= rom_array(30125);
		when "0111010110101110" => data_out <= rom_array(30126);
		when "0111010110101111" => data_out <= rom_array(30127);
		when "0111010110110000" => data_out <= rom_array(30128);
		when "0111010110110001" => data_out <= rom_array(30129);
		when "0111010110110010" => data_out <= rom_array(30130);
		when "0111010110110011" => data_out <= rom_array(30131);
		when "0111010110110100" => data_out <= rom_array(30132);
		when "0111010110110101" => data_out <= rom_array(30133);
		when "0111010110110110" => data_out <= rom_array(30134);
		when "0111010110110111" => data_out <= rom_array(30135);
		when "0111010110111000" => data_out <= rom_array(30136);
		when "0111010110111001" => data_out <= rom_array(30137);
		when "0111010110111010" => data_out <= rom_array(30138);
		when "0111010110111011" => data_out <= rom_array(30139);
		when "0111010110111100" => data_out <= rom_array(30140);
		when "0111010110111101" => data_out <= rom_array(30141);
		when "0111010110111110" => data_out <= rom_array(30142);
		when "0111010110111111" => data_out <= rom_array(30143);
		when "0111010111000000" => data_out <= rom_array(30144);
		when "0111010111000001" => data_out <= rom_array(30145);
		when "0111010111000010" => data_out <= rom_array(30146);
		when "0111010111000011" => data_out <= rom_array(30147);
		when "0111010111000100" => data_out <= rom_array(30148);
		when "0111010111000101" => data_out <= rom_array(30149);
		when "0111010111000110" => data_out <= rom_array(30150);
		when "0111010111000111" => data_out <= rom_array(30151);
		when "0111010111001000" => data_out <= rom_array(30152);
		when "0111010111001001" => data_out <= rom_array(30153);
		when "0111010111001010" => data_out <= rom_array(30154);
		when "0111010111001011" => data_out <= rom_array(30155);
		when "0111010111001100" => data_out <= rom_array(30156);
		when "0111010111001101" => data_out <= rom_array(30157);
		when "0111010111001110" => data_out <= rom_array(30158);
		when "0111010111001111" => data_out <= rom_array(30159);
		when "0111010111010000" => data_out <= rom_array(30160);
		when "0111010111010001" => data_out <= rom_array(30161);
		when "0111010111010010" => data_out <= rom_array(30162);
		when "0111010111010011" => data_out <= rom_array(30163);
		when "0111010111010100" => data_out <= rom_array(30164);
		when "0111010111010101" => data_out <= rom_array(30165);
		when "0111010111010110" => data_out <= rom_array(30166);
		when "0111010111010111" => data_out <= rom_array(30167);
		when "0111010111011000" => data_out <= rom_array(30168);
		when "0111010111011001" => data_out <= rom_array(30169);
		when "0111010111011010" => data_out <= rom_array(30170);
		when "0111010111011011" => data_out <= rom_array(30171);
		when "0111010111011100" => data_out <= rom_array(30172);
		when "0111010111011101" => data_out <= rom_array(30173);
		when "0111010111011110" => data_out <= rom_array(30174);
		when "0111010111011111" => data_out <= rom_array(30175);
		when "0111010111100000" => data_out <= rom_array(30176);
		when "0111010111100001" => data_out <= rom_array(30177);
		when "0111010111100010" => data_out <= rom_array(30178);
		when "0111010111100011" => data_out <= rom_array(30179);
		when "0111010111100100" => data_out <= rom_array(30180);
		when "0111010111100101" => data_out <= rom_array(30181);
		when "0111010111100110" => data_out <= rom_array(30182);
		when "0111010111100111" => data_out <= rom_array(30183);
		when "0111010111101000" => data_out <= rom_array(30184);
		when "0111010111101001" => data_out <= rom_array(30185);
		when "0111010111101010" => data_out <= rom_array(30186);
		when "0111010111101011" => data_out <= rom_array(30187);
		when "0111010111101100" => data_out <= rom_array(30188);
		when "0111010111101101" => data_out <= rom_array(30189);
		when "0111010111101110" => data_out <= rom_array(30190);
		when "0111010111101111" => data_out <= rom_array(30191);
		when "0111010111110000" => data_out <= rom_array(30192);
		when "0111010111110001" => data_out <= rom_array(30193);
		when "0111010111110010" => data_out <= rom_array(30194);
		when "0111010111110011" => data_out <= rom_array(30195);
		when "0111010111110100" => data_out <= rom_array(30196);
		when "0111010111110101" => data_out <= rom_array(30197);
		when "0111010111110110" => data_out <= rom_array(30198);
		when "0111010111110111" => data_out <= rom_array(30199);
		when "0111010111111000" => data_out <= rom_array(30200);
		when "0111010111111001" => data_out <= rom_array(30201);
		when "0111010111111010" => data_out <= rom_array(30202);
		when "0111010111111011" => data_out <= rom_array(30203);
		when "0111010111111100" => data_out <= rom_array(30204);
		when "0111010111111101" => data_out <= rom_array(30205);
		when "0111010111111110" => data_out <= rom_array(30206);
		when "0111010111111111" => data_out <= rom_array(30207);
		when "0111011000000000" => data_out <= rom_array(30208);
		when "0111011000000001" => data_out <= rom_array(30209);
		when "0111011000000010" => data_out <= rom_array(30210);
		when "0111011000000011" => data_out <= rom_array(30211);
		when "0111011000000100" => data_out <= rom_array(30212);
		when "0111011000000101" => data_out <= rom_array(30213);
		when "0111011000000110" => data_out <= rom_array(30214);
		when "0111011000000111" => data_out <= rom_array(30215);
		when "0111011000001000" => data_out <= rom_array(30216);
		when "0111011000001001" => data_out <= rom_array(30217);
		when "0111011000001010" => data_out <= rom_array(30218);
		when "0111011000001011" => data_out <= rom_array(30219);
		when "0111011000001100" => data_out <= rom_array(30220);
		when "0111011000001101" => data_out <= rom_array(30221);
		when "0111011000001110" => data_out <= rom_array(30222);
		when "0111011000001111" => data_out <= rom_array(30223);
		when "0111011000010000" => data_out <= rom_array(30224);
		when "0111011000010001" => data_out <= rom_array(30225);
		when "0111011000010010" => data_out <= rom_array(30226);
		when "0111011000010011" => data_out <= rom_array(30227);
		when "0111011000010100" => data_out <= rom_array(30228);
		when "0111011000010101" => data_out <= rom_array(30229);
		when "0111011000010110" => data_out <= rom_array(30230);
		when "0111011000010111" => data_out <= rom_array(30231);
		when "0111011000011000" => data_out <= rom_array(30232);
		when "0111011000011001" => data_out <= rom_array(30233);
		when "0111011000011010" => data_out <= rom_array(30234);
		when "0111011000011011" => data_out <= rom_array(30235);
		when "0111011000011100" => data_out <= rom_array(30236);
		when "0111011000011101" => data_out <= rom_array(30237);
		when "0111011000011110" => data_out <= rom_array(30238);
		when "0111011000011111" => data_out <= rom_array(30239);
		when "0111011000100000" => data_out <= rom_array(30240);
		when "0111011000100001" => data_out <= rom_array(30241);
		when "0111011000100010" => data_out <= rom_array(30242);
		when "0111011000100011" => data_out <= rom_array(30243);
		when "0111011000100100" => data_out <= rom_array(30244);
		when "0111011000100101" => data_out <= rom_array(30245);
		when "0111011000100110" => data_out <= rom_array(30246);
		when "0111011000100111" => data_out <= rom_array(30247);
		when "0111011000101000" => data_out <= rom_array(30248);
		when "0111011000101001" => data_out <= rom_array(30249);
		when "0111011000101010" => data_out <= rom_array(30250);
		when "0111011000101011" => data_out <= rom_array(30251);
		when "0111011000101100" => data_out <= rom_array(30252);
		when "0111011000101101" => data_out <= rom_array(30253);
		when "0111011000101110" => data_out <= rom_array(30254);
		when "0111011000101111" => data_out <= rom_array(30255);
		when "0111011000110000" => data_out <= rom_array(30256);
		when "0111011000110001" => data_out <= rom_array(30257);
		when "0111011000110010" => data_out <= rom_array(30258);
		when "0111011000110011" => data_out <= rom_array(30259);
		when "0111011000110100" => data_out <= rom_array(30260);
		when "0111011000110101" => data_out <= rom_array(30261);
		when "0111011000110110" => data_out <= rom_array(30262);
		when "0111011000110111" => data_out <= rom_array(30263);
		when "0111011000111000" => data_out <= rom_array(30264);
		when "0111011000111001" => data_out <= rom_array(30265);
		when "0111011000111010" => data_out <= rom_array(30266);
		when "0111011000111011" => data_out <= rom_array(30267);
		when "0111011000111100" => data_out <= rom_array(30268);
		when "0111011000111101" => data_out <= rom_array(30269);
		when "0111011000111110" => data_out <= rom_array(30270);
		when "0111011000111111" => data_out <= rom_array(30271);
		when "0111011001000000" => data_out <= rom_array(30272);
		when "0111011001000001" => data_out <= rom_array(30273);
		when "0111011001000010" => data_out <= rom_array(30274);
		when "0111011001000011" => data_out <= rom_array(30275);
		when "0111011001000100" => data_out <= rom_array(30276);
		when "0111011001000101" => data_out <= rom_array(30277);
		when "0111011001000110" => data_out <= rom_array(30278);
		when "0111011001000111" => data_out <= rom_array(30279);
		when "0111011001001000" => data_out <= rom_array(30280);
		when "0111011001001001" => data_out <= rom_array(30281);
		when "0111011001001010" => data_out <= rom_array(30282);
		when "0111011001001011" => data_out <= rom_array(30283);
		when "0111011001001100" => data_out <= rom_array(30284);
		when "0111011001001101" => data_out <= rom_array(30285);
		when "0111011001001110" => data_out <= rom_array(30286);
		when "0111011001001111" => data_out <= rom_array(30287);
		when "0111011001010000" => data_out <= rom_array(30288);
		when "0111011001010001" => data_out <= rom_array(30289);
		when "0111011001010010" => data_out <= rom_array(30290);
		when "0111011001010011" => data_out <= rom_array(30291);
		when "0111011001010100" => data_out <= rom_array(30292);
		when "0111011001010101" => data_out <= rom_array(30293);
		when "0111011001010110" => data_out <= rom_array(30294);
		when "0111011001010111" => data_out <= rom_array(30295);
		when "0111011001011000" => data_out <= rom_array(30296);
		when "0111011001011001" => data_out <= rom_array(30297);
		when "0111011001011010" => data_out <= rom_array(30298);
		when "0111011001011011" => data_out <= rom_array(30299);
		when "0111011001011100" => data_out <= rom_array(30300);
		when "0111011001011101" => data_out <= rom_array(30301);
		when "0111011001011110" => data_out <= rom_array(30302);
		when "0111011001011111" => data_out <= rom_array(30303);
		when "0111011001100000" => data_out <= rom_array(30304);
		when "0111011001100001" => data_out <= rom_array(30305);
		when "0111011001100010" => data_out <= rom_array(30306);
		when "0111011001100011" => data_out <= rom_array(30307);
		when "0111011001100100" => data_out <= rom_array(30308);
		when "0111011001100101" => data_out <= rom_array(30309);
		when "0111011001100110" => data_out <= rom_array(30310);
		when "0111011001100111" => data_out <= rom_array(30311);
		when "0111011001101000" => data_out <= rom_array(30312);
		when "0111011001101001" => data_out <= rom_array(30313);
		when "0111011001101010" => data_out <= rom_array(30314);
		when "0111011001101011" => data_out <= rom_array(30315);
		when "0111011001101100" => data_out <= rom_array(30316);
		when "0111011001101101" => data_out <= rom_array(30317);
		when "0111011001101110" => data_out <= rom_array(30318);
		when "0111011001101111" => data_out <= rom_array(30319);
		when "0111011001110000" => data_out <= rom_array(30320);
		when "0111011001110001" => data_out <= rom_array(30321);
		when "0111011001110010" => data_out <= rom_array(30322);
		when "0111011001110011" => data_out <= rom_array(30323);
		when "0111011001110100" => data_out <= rom_array(30324);
		when "0111011001110101" => data_out <= rom_array(30325);
		when "0111011001110110" => data_out <= rom_array(30326);
		when "0111011001110111" => data_out <= rom_array(30327);
		when "0111011001111000" => data_out <= rom_array(30328);
		when "0111011001111001" => data_out <= rom_array(30329);
		when "0111011001111010" => data_out <= rom_array(30330);
		when "0111011001111011" => data_out <= rom_array(30331);
		when "0111011001111100" => data_out <= rom_array(30332);
		when "0111011001111101" => data_out <= rom_array(30333);
		when "0111011001111110" => data_out <= rom_array(30334);
		when "0111011001111111" => data_out <= rom_array(30335);
		when "0111011010000000" => data_out <= rom_array(30336);
		when "0111011010000001" => data_out <= rom_array(30337);
		when "0111011010000010" => data_out <= rom_array(30338);
		when "0111011010000011" => data_out <= rom_array(30339);
		when "0111011010000100" => data_out <= rom_array(30340);
		when "0111011010000101" => data_out <= rom_array(30341);
		when "0111011010000110" => data_out <= rom_array(30342);
		when "0111011010000111" => data_out <= rom_array(30343);
		when "0111011010001000" => data_out <= rom_array(30344);
		when "0111011010001001" => data_out <= rom_array(30345);
		when "0111011010001010" => data_out <= rom_array(30346);
		when "0111011010001011" => data_out <= rom_array(30347);
		when "0111011010001100" => data_out <= rom_array(30348);
		when "0111011010001101" => data_out <= rom_array(30349);
		when "0111011010001110" => data_out <= rom_array(30350);
		when "0111011010001111" => data_out <= rom_array(30351);
		when "0111011010010000" => data_out <= rom_array(30352);
		when "0111011010010001" => data_out <= rom_array(30353);
		when "0111011010010010" => data_out <= rom_array(30354);
		when "0111011010010011" => data_out <= rom_array(30355);
		when "0111011010010100" => data_out <= rom_array(30356);
		when "0111011010010101" => data_out <= rom_array(30357);
		when "0111011010010110" => data_out <= rom_array(30358);
		when "0111011010010111" => data_out <= rom_array(30359);
		when "0111011010011000" => data_out <= rom_array(30360);
		when "0111011010011001" => data_out <= rom_array(30361);
		when "0111011010011010" => data_out <= rom_array(30362);
		when "0111011010011011" => data_out <= rom_array(30363);
		when "0111011010011100" => data_out <= rom_array(30364);
		when "0111011010011101" => data_out <= rom_array(30365);
		when "0111011010011110" => data_out <= rom_array(30366);
		when "0111011010011111" => data_out <= rom_array(30367);
		when "0111011010100000" => data_out <= rom_array(30368);
		when "0111011010100001" => data_out <= rom_array(30369);
		when "0111011010100010" => data_out <= rom_array(30370);
		when "0111011010100011" => data_out <= rom_array(30371);
		when "0111011010100100" => data_out <= rom_array(30372);
		when "0111011010100101" => data_out <= rom_array(30373);
		when "0111011010100110" => data_out <= rom_array(30374);
		when "0111011010100111" => data_out <= rom_array(30375);
		when "0111011010101000" => data_out <= rom_array(30376);
		when "0111011010101001" => data_out <= rom_array(30377);
		when "0111011010101010" => data_out <= rom_array(30378);
		when "0111011010101011" => data_out <= rom_array(30379);
		when "0111011010101100" => data_out <= rom_array(30380);
		when "0111011010101101" => data_out <= rom_array(30381);
		when "0111011010101110" => data_out <= rom_array(30382);
		when "0111011010101111" => data_out <= rom_array(30383);
		when "0111011010110000" => data_out <= rom_array(30384);
		when "0111011010110001" => data_out <= rom_array(30385);
		when "0111011010110010" => data_out <= rom_array(30386);
		when "0111011010110011" => data_out <= rom_array(30387);
		when "0111011010110100" => data_out <= rom_array(30388);
		when "0111011010110101" => data_out <= rom_array(30389);
		when "0111011010110110" => data_out <= rom_array(30390);
		when "0111011010110111" => data_out <= rom_array(30391);
		when "0111011010111000" => data_out <= rom_array(30392);
		when "0111011010111001" => data_out <= rom_array(30393);
		when "0111011010111010" => data_out <= rom_array(30394);
		when "0111011010111011" => data_out <= rom_array(30395);
		when "0111011010111100" => data_out <= rom_array(30396);
		when "0111011010111101" => data_out <= rom_array(30397);
		when "0111011010111110" => data_out <= rom_array(30398);
		when "0111011010111111" => data_out <= rom_array(30399);
		when "0111011011000000" => data_out <= rom_array(30400);
		when "0111011011000001" => data_out <= rom_array(30401);
		when "0111011011000010" => data_out <= rom_array(30402);
		when "0111011011000011" => data_out <= rom_array(30403);
		when "0111011011000100" => data_out <= rom_array(30404);
		when "0111011011000101" => data_out <= rom_array(30405);
		when "0111011011000110" => data_out <= rom_array(30406);
		when "0111011011000111" => data_out <= rom_array(30407);
		when "0111011011001000" => data_out <= rom_array(30408);
		when "0111011011001001" => data_out <= rom_array(30409);
		when "0111011011001010" => data_out <= rom_array(30410);
		when "0111011011001011" => data_out <= rom_array(30411);
		when "0111011011001100" => data_out <= rom_array(30412);
		when "0111011011001101" => data_out <= rom_array(30413);
		when "0111011011001110" => data_out <= rom_array(30414);
		when "0111011011001111" => data_out <= rom_array(30415);
		when "0111011011010000" => data_out <= rom_array(30416);
		when "0111011011010001" => data_out <= rom_array(30417);
		when "0111011011010010" => data_out <= rom_array(30418);
		when "0111011011010011" => data_out <= rom_array(30419);
		when "0111011011010100" => data_out <= rom_array(30420);
		when "0111011011010101" => data_out <= rom_array(30421);
		when "0111011011010110" => data_out <= rom_array(30422);
		when "0111011011010111" => data_out <= rom_array(30423);
		when "0111011011011000" => data_out <= rom_array(30424);
		when "0111011011011001" => data_out <= rom_array(30425);
		when "0111011011011010" => data_out <= rom_array(30426);
		when "0111011011011011" => data_out <= rom_array(30427);
		when "0111011011011100" => data_out <= rom_array(30428);
		when "0111011011011101" => data_out <= rom_array(30429);
		when "0111011011011110" => data_out <= rom_array(30430);
		when "0111011011011111" => data_out <= rom_array(30431);
		when "0111011011100000" => data_out <= rom_array(30432);
		when "0111011011100001" => data_out <= rom_array(30433);
		when "0111011011100010" => data_out <= rom_array(30434);
		when "0111011011100011" => data_out <= rom_array(30435);
		when "0111011011100100" => data_out <= rom_array(30436);
		when "0111011011100101" => data_out <= rom_array(30437);
		when "0111011011100110" => data_out <= rom_array(30438);
		when "0111011011100111" => data_out <= rom_array(30439);
		when "0111011011101000" => data_out <= rom_array(30440);
		when "0111011011101001" => data_out <= rom_array(30441);
		when "0111011011101010" => data_out <= rom_array(30442);
		when "0111011011101011" => data_out <= rom_array(30443);
		when "0111011011101100" => data_out <= rom_array(30444);
		when "0111011011101101" => data_out <= rom_array(30445);
		when "0111011011101110" => data_out <= rom_array(30446);
		when "0111011011101111" => data_out <= rom_array(30447);
		when "0111011011110000" => data_out <= rom_array(30448);
		when "0111011011110001" => data_out <= rom_array(30449);
		when "0111011011110010" => data_out <= rom_array(30450);
		when "0111011011110011" => data_out <= rom_array(30451);
		when "0111011011110100" => data_out <= rom_array(30452);
		when "0111011011110101" => data_out <= rom_array(30453);
		when "0111011011110110" => data_out <= rom_array(30454);
		when "0111011011110111" => data_out <= rom_array(30455);
		when "0111011011111000" => data_out <= rom_array(30456);
		when "0111011011111001" => data_out <= rom_array(30457);
		when "0111011011111010" => data_out <= rom_array(30458);
		when "0111011011111011" => data_out <= rom_array(30459);
		when "0111011011111100" => data_out <= rom_array(30460);
		when "0111011011111101" => data_out <= rom_array(30461);
		when "0111011011111110" => data_out <= rom_array(30462);
		when "0111011011111111" => data_out <= rom_array(30463);
		when "0111011100000000" => data_out <= rom_array(30464);
		when "0111011100000001" => data_out <= rom_array(30465);
		when "0111011100000010" => data_out <= rom_array(30466);
		when "0111011100000011" => data_out <= rom_array(30467);
		when "0111011100000100" => data_out <= rom_array(30468);
		when "0111011100000101" => data_out <= rom_array(30469);
		when "0111011100000110" => data_out <= rom_array(30470);
		when "0111011100000111" => data_out <= rom_array(30471);
		when "0111011100001000" => data_out <= rom_array(30472);
		when "0111011100001001" => data_out <= rom_array(30473);
		when "0111011100001010" => data_out <= rom_array(30474);
		when "0111011100001011" => data_out <= rom_array(30475);
		when "0111011100001100" => data_out <= rom_array(30476);
		when "0111011100001101" => data_out <= rom_array(30477);
		when "0111011100001110" => data_out <= rom_array(30478);
		when "0111011100001111" => data_out <= rom_array(30479);
		when "0111011100010000" => data_out <= rom_array(30480);
		when "0111011100010001" => data_out <= rom_array(30481);
		when "0111011100010010" => data_out <= rom_array(30482);
		when "0111011100010011" => data_out <= rom_array(30483);
		when "0111011100010100" => data_out <= rom_array(30484);
		when "0111011100010101" => data_out <= rom_array(30485);
		when "0111011100010110" => data_out <= rom_array(30486);
		when "0111011100010111" => data_out <= rom_array(30487);
		when "0111011100011000" => data_out <= rom_array(30488);
		when "0111011100011001" => data_out <= rom_array(30489);
		when "0111011100011010" => data_out <= rom_array(30490);
		when "0111011100011011" => data_out <= rom_array(30491);
		when "0111011100011100" => data_out <= rom_array(30492);
		when "0111011100011101" => data_out <= rom_array(30493);
		when "0111011100011110" => data_out <= rom_array(30494);
		when "0111011100011111" => data_out <= rom_array(30495);
		when "0111011100100000" => data_out <= rom_array(30496);
		when "0111011100100001" => data_out <= rom_array(30497);
		when "0111011100100010" => data_out <= rom_array(30498);
		when "0111011100100011" => data_out <= rom_array(30499);
		when "0111011100100100" => data_out <= rom_array(30500);
		when "0111011100100101" => data_out <= rom_array(30501);
		when "0111011100100110" => data_out <= rom_array(30502);
		when "0111011100100111" => data_out <= rom_array(30503);
		when "0111011100101000" => data_out <= rom_array(30504);
		when "0111011100101001" => data_out <= rom_array(30505);
		when "0111011100101010" => data_out <= rom_array(30506);
		when "0111011100101011" => data_out <= rom_array(30507);
		when "0111011100101100" => data_out <= rom_array(30508);
		when "0111011100101101" => data_out <= rom_array(30509);
		when "0111011100101110" => data_out <= rom_array(30510);
		when "0111011100101111" => data_out <= rom_array(30511);
		when "0111011100110000" => data_out <= rom_array(30512);
		when "0111011100110001" => data_out <= rom_array(30513);
		when "0111011100110010" => data_out <= rom_array(30514);
		when "0111011100110011" => data_out <= rom_array(30515);
		when "0111011100110100" => data_out <= rom_array(30516);
		when "0111011100110101" => data_out <= rom_array(30517);
		when "0111011100110110" => data_out <= rom_array(30518);
		when "0111011100110111" => data_out <= rom_array(30519);
		when "0111011100111000" => data_out <= rom_array(30520);
		when "0111011100111001" => data_out <= rom_array(30521);
		when "0111011100111010" => data_out <= rom_array(30522);
		when "0111011100111011" => data_out <= rom_array(30523);
		when "0111011100111100" => data_out <= rom_array(30524);
		when "0111011100111101" => data_out <= rom_array(30525);
		when "0111011100111110" => data_out <= rom_array(30526);
		when "0111011100111111" => data_out <= rom_array(30527);
		when "0111011101000000" => data_out <= rom_array(30528);
		when "0111011101000001" => data_out <= rom_array(30529);
		when "0111011101000010" => data_out <= rom_array(30530);
		when "0111011101000011" => data_out <= rom_array(30531);
		when "0111011101000100" => data_out <= rom_array(30532);
		when "0111011101000101" => data_out <= rom_array(30533);
		when "0111011101000110" => data_out <= rom_array(30534);
		when "0111011101000111" => data_out <= rom_array(30535);
		when "0111011101001000" => data_out <= rom_array(30536);
		when "0111011101001001" => data_out <= rom_array(30537);
		when "0111011101001010" => data_out <= rom_array(30538);
		when "0111011101001011" => data_out <= rom_array(30539);
		when "0111011101001100" => data_out <= rom_array(30540);
		when "0111011101001101" => data_out <= rom_array(30541);
		when "0111011101001110" => data_out <= rom_array(30542);
		when "0111011101001111" => data_out <= rom_array(30543);
		when "0111011101010000" => data_out <= rom_array(30544);
		when "0111011101010001" => data_out <= rom_array(30545);
		when "0111011101010010" => data_out <= rom_array(30546);
		when "0111011101010011" => data_out <= rom_array(30547);
		when "0111011101010100" => data_out <= rom_array(30548);
		when "0111011101010101" => data_out <= rom_array(30549);
		when "0111011101010110" => data_out <= rom_array(30550);
		when "0111011101010111" => data_out <= rom_array(30551);
		when "0111011101011000" => data_out <= rom_array(30552);
		when "0111011101011001" => data_out <= rom_array(30553);
		when "0111011101011010" => data_out <= rom_array(30554);
		when "0111011101011011" => data_out <= rom_array(30555);
		when "0111011101011100" => data_out <= rom_array(30556);
		when "0111011101011101" => data_out <= rom_array(30557);
		when "0111011101011110" => data_out <= rom_array(30558);
		when "0111011101011111" => data_out <= rom_array(30559);
		when "0111011101100000" => data_out <= rom_array(30560);
		when "0111011101100001" => data_out <= rom_array(30561);
		when "0111011101100010" => data_out <= rom_array(30562);
		when "0111011101100011" => data_out <= rom_array(30563);
		when "0111011101100100" => data_out <= rom_array(30564);
		when "0111011101100101" => data_out <= rom_array(30565);
		when "0111011101100110" => data_out <= rom_array(30566);
		when "0111011101100111" => data_out <= rom_array(30567);
		when "0111011101101000" => data_out <= rom_array(30568);
		when "0111011101101001" => data_out <= rom_array(30569);
		when "0111011101101010" => data_out <= rom_array(30570);
		when "0111011101101011" => data_out <= rom_array(30571);
		when "0111011101101100" => data_out <= rom_array(30572);
		when "0111011101101101" => data_out <= rom_array(30573);
		when "0111011101101110" => data_out <= rom_array(30574);
		when "0111011101101111" => data_out <= rom_array(30575);
		when "0111011101110000" => data_out <= rom_array(30576);
		when "0111011101110001" => data_out <= rom_array(30577);
		when "0111011101110010" => data_out <= rom_array(30578);
		when "0111011101110011" => data_out <= rom_array(30579);
		when "0111011101110100" => data_out <= rom_array(30580);
		when "0111011101110101" => data_out <= rom_array(30581);
		when "0111011101110110" => data_out <= rom_array(30582);
		when "0111011101110111" => data_out <= rom_array(30583);
		when "0111011101111000" => data_out <= rom_array(30584);
		when "0111011101111001" => data_out <= rom_array(30585);
		when "0111011101111010" => data_out <= rom_array(30586);
		when "0111011101111011" => data_out <= rom_array(30587);
		when "0111011101111100" => data_out <= rom_array(30588);
		when "0111011101111101" => data_out <= rom_array(30589);
		when "0111011101111110" => data_out <= rom_array(30590);
		when "0111011101111111" => data_out <= rom_array(30591);
		when "0111011110000000" => data_out <= rom_array(30592);
		when "0111011110000001" => data_out <= rom_array(30593);
		when "0111011110000010" => data_out <= rom_array(30594);
		when "0111011110000011" => data_out <= rom_array(30595);
		when "0111011110000100" => data_out <= rom_array(30596);
		when "0111011110000101" => data_out <= rom_array(30597);
		when "0111011110000110" => data_out <= rom_array(30598);
		when "0111011110000111" => data_out <= rom_array(30599);
		when "0111011110001000" => data_out <= rom_array(30600);
		when "0111011110001001" => data_out <= rom_array(30601);
		when "0111011110001010" => data_out <= rom_array(30602);
		when "0111011110001011" => data_out <= rom_array(30603);
		when "0111011110001100" => data_out <= rom_array(30604);
		when "0111011110001101" => data_out <= rom_array(30605);
		when "0111011110001110" => data_out <= rom_array(30606);
		when "0111011110001111" => data_out <= rom_array(30607);
		when "0111011110010000" => data_out <= rom_array(30608);
		when "0111011110010001" => data_out <= rom_array(30609);
		when "0111011110010010" => data_out <= rom_array(30610);
		when "0111011110010011" => data_out <= rom_array(30611);
		when "0111011110010100" => data_out <= rom_array(30612);
		when "0111011110010101" => data_out <= rom_array(30613);
		when "0111011110010110" => data_out <= rom_array(30614);
		when "0111011110010111" => data_out <= rom_array(30615);
		when "0111011110011000" => data_out <= rom_array(30616);
		when "0111011110011001" => data_out <= rom_array(30617);
		when "0111011110011010" => data_out <= rom_array(30618);
		when "0111011110011011" => data_out <= rom_array(30619);
		when "0111011110011100" => data_out <= rom_array(30620);
		when "0111011110011101" => data_out <= rom_array(30621);
		when "0111011110011110" => data_out <= rom_array(30622);
		when "0111011110011111" => data_out <= rom_array(30623);
		when "0111011110100000" => data_out <= rom_array(30624);
		when "0111011110100001" => data_out <= rom_array(30625);
		when "0111011110100010" => data_out <= rom_array(30626);
		when "0111011110100011" => data_out <= rom_array(30627);
		when "0111011110100100" => data_out <= rom_array(30628);
		when "0111011110100101" => data_out <= rom_array(30629);
		when "0111011110100110" => data_out <= rom_array(30630);
		when "0111011110100111" => data_out <= rom_array(30631);
		when "0111011110101000" => data_out <= rom_array(30632);
		when "0111011110101001" => data_out <= rom_array(30633);
		when "0111011110101010" => data_out <= rom_array(30634);
		when "0111011110101011" => data_out <= rom_array(30635);
		when "0111011110101100" => data_out <= rom_array(30636);
		when "0111011110101101" => data_out <= rom_array(30637);
		when "0111011110101110" => data_out <= rom_array(30638);
		when "0111011110101111" => data_out <= rom_array(30639);
		when "0111011110110000" => data_out <= rom_array(30640);
		when "0111011110110001" => data_out <= rom_array(30641);
		when "0111011110110010" => data_out <= rom_array(30642);
		when "0111011110110011" => data_out <= rom_array(30643);
		when "0111011110110100" => data_out <= rom_array(30644);
		when "0111011110110101" => data_out <= rom_array(30645);
		when "0111011110110110" => data_out <= rom_array(30646);
		when "0111011110110111" => data_out <= rom_array(30647);
		when "0111011110111000" => data_out <= rom_array(30648);
		when "0111011110111001" => data_out <= rom_array(30649);
		when "0111011110111010" => data_out <= rom_array(30650);
		when "0111011110111011" => data_out <= rom_array(30651);
		when "0111011110111100" => data_out <= rom_array(30652);
		when "0111011110111101" => data_out <= rom_array(30653);
		when "0111011110111110" => data_out <= rom_array(30654);
		when "0111011110111111" => data_out <= rom_array(30655);
		when "0111011111000000" => data_out <= rom_array(30656);
		when "0111011111000001" => data_out <= rom_array(30657);
		when "0111011111000010" => data_out <= rom_array(30658);
		when "0111011111000011" => data_out <= rom_array(30659);
		when "0111011111000100" => data_out <= rom_array(30660);
		when "0111011111000101" => data_out <= rom_array(30661);
		when "0111011111000110" => data_out <= rom_array(30662);
		when "0111011111000111" => data_out <= rom_array(30663);
		when "0111011111001000" => data_out <= rom_array(30664);
		when "0111011111001001" => data_out <= rom_array(30665);
		when "0111011111001010" => data_out <= rom_array(30666);
		when "0111011111001011" => data_out <= rom_array(30667);
		when "0111011111001100" => data_out <= rom_array(30668);
		when "0111011111001101" => data_out <= rom_array(30669);
		when "0111011111001110" => data_out <= rom_array(30670);
		when "0111011111001111" => data_out <= rom_array(30671);
		when "0111011111010000" => data_out <= rom_array(30672);
		when "0111011111010001" => data_out <= rom_array(30673);
		when "0111011111010010" => data_out <= rom_array(30674);
		when "0111011111010011" => data_out <= rom_array(30675);
		when "0111011111010100" => data_out <= rom_array(30676);
		when "0111011111010101" => data_out <= rom_array(30677);
		when "0111011111010110" => data_out <= rom_array(30678);
		when "0111011111010111" => data_out <= rom_array(30679);
		when "0111011111011000" => data_out <= rom_array(30680);
		when "0111011111011001" => data_out <= rom_array(30681);
		when "0111011111011010" => data_out <= rom_array(30682);
		when "0111011111011011" => data_out <= rom_array(30683);
		when "0111011111011100" => data_out <= rom_array(30684);
		when "0111011111011101" => data_out <= rom_array(30685);
		when "0111011111011110" => data_out <= rom_array(30686);
		when "0111011111011111" => data_out <= rom_array(30687);
		when "0111011111100000" => data_out <= rom_array(30688);
		when "0111011111100001" => data_out <= rom_array(30689);
		when "0111011111100010" => data_out <= rom_array(30690);
		when "0111011111100011" => data_out <= rom_array(30691);
		when "0111011111100100" => data_out <= rom_array(30692);
		when "0111011111100101" => data_out <= rom_array(30693);
		when "0111011111100110" => data_out <= rom_array(30694);
		when "0111011111100111" => data_out <= rom_array(30695);
		when "0111011111101000" => data_out <= rom_array(30696);
		when "0111011111101001" => data_out <= rom_array(30697);
		when "0111011111101010" => data_out <= rom_array(30698);
		when "0111011111101011" => data_out <= rom_array(30699);
		when "0111011111101100" => data_out <= rom_array(30700);
		when "0111011111101101" => data_out <= rom_array(30701);
		when "0111011111101110" => data_out <= rom_array(30702);
		when "0111011111101111" => data_out <= rom_array(30703);
		when "0111011111110000" => data_out <= rom_array(30704);
		when "0111011111110001" => data_out <= rom_array(30705);
		when "0111011111110010" => data_out <= rom_array(30706);
		when "0111011111110011" => data_out <= rom_array(30707);
		when "0111011111110100" => data_out <= rom_array(30708);
		when "0111011111110101" => data_out <= rom_array(30709);
		when "0111011111110110" => data_out <= rom_array(30710);
		when "0111011111110111" => data_out <= rom_array(30711);
		when "0111011111111000" => data_out <= rom_array(30712);
		when "0111011111111001" => data_out <= rom_array(30713);
		when "0111011111111010" => data_out <= rom_array(30714);
		when "0111011111111011" => data_out <= rom_array(30715);
		when "0111011111111100" => data_out <= rom_array(30716);
		when "0111011111111101" => data_out <= rom_array(30717);
		when "0111011111111110" => data_out <= rom_array(30718);
		when "0111011111111111" => data_out <= rom_array(30719);
		when "0111100000000000" => data_out <= rom_array(30720);
		when "0111100000000001" => data_out <= rom_array(30721);
		when "0111100000000010" => data_out <= rom_array(30722);
		when "0111100000000011" => data_out <= rom_array(30723);
		when "0111100000000100" => data_out <= rom_array(30724);
		when "0111100000000101" => data_out <= rom_array(30725);
		when "0111100000000110" => data_out <= rom_array(30726);
		when "0111100000000111" => data_out <= rom_array(30727);
		when "0111100000001000" => data_out <= rom_array(30728);
		when "0111100000001001" => data_out <= rom_array(30729);
		when "0111100000001010" => data_out <= rom_array(30730);
		when "0111100000001011" => data_out <= rom_array(30731);
		when "0111100000001100" => data_out <= rom_array(30732);
		when "0111100000001101" => data_out <= rom_array(30733);
		when "0111100000001110" => data_out <= rom_array(30734);
		when "0111100000001111" => data_out <= rom_array(30735);
		when "0111100000010000" => data_out <= rom_array(30736);
		when "0111100000010001" => data_out <= rom_array(30737);
		when "0111100000010010" => data_out <= rom_array(30738);
		when "0111100000010011" => data_out <= rom_array(30739);
		when "0111100000010100" => data_out <= rom_array(30740);
		when "0111100000010101" => data_out <= rom_array(30741);
		when "0111100000010110" => data_out <= rom_array(30742);
		when "0111100000010111" => data_out <= rom_array(30743);
		when "0111100000011000" => data_out <= rom_array(30744);
		when "0111100000011001" => data_out <= rom_array(30745);
		when "0111100000011010" => data_out <= rom_array(30746);
		when "0111100000011011" => data_out <= rom_array(30747);
		when "0111100000011100" => data_out <= rom_array(30748);
		when "0111100000011101" => data_out <= rom_array(30749);
		when "0111100000011110" => data_out <= rom_array(30750);
		when "0111100000011111" => data_out <= rom_array(30751);
		when "0111100000100000" => data_out <= rom_array(30752);
		when "0111100000100001" => data_out <= rom_array(30753);
		when "0111100000100010" => data_out <= rom_array(30754);
		when "0111100000100011" => data_out <= rom_array(30755);
		when "0111100000100100" => data_out <= rom_array(30756);
		when "0111100000100101" => data_out <= rom_array(30757);
		when "0111100000100110" => data_out <= rom_array(30758);
		when "0111100000100111" => data_out <= rom_array(30759);
		when "0111100000101000" => data_out <= rom_array(30760);
		when "0111100000101001" => data_out <= rom_array(30761);
		when "0111100000101010" => data_out <= rom_array(30762);
		when "0111100000101011" => data_out <= rom_array(30763);
		when "0111100000101100" => data_out <= rom_array(30764);
		when "0111100000101101" => data_out <= rom_array(30765);
		when "0111100000101110" => data_out <= rom_array(30766);
		when "0111100000101111" => data_out <= rom_array(30767);
		when "0111100000110000" => data_out <= rom_array(30768);
		when "0111100000110001" => data_out <= rom_array(30769);
		when "0111100000110010" => data_out <= rom_array(30770);
		when "0111100000110011" => data_out <= rom_array(30771);
		when "0111100000110100" => data_out <= rom_array(30772);
		when "0111100000110101" => data_out <= rom_array(30773);
		when "0111100000110110" => data_out <= rom_array(30774);
		when "0111100000110111" => data_out <= rom_array(30775);
		when "0111100000111000" => data_out <= rom_array(30776);
		when "0111100000111001" => data_out <= rom_array(30777);
		when "0111100000111010" => data_out <= rom_array(30778);
		when "0111100000111011" => data_out <= rom_array(30779);
		when "0111100000111100" => data_out <= rom_array(30780);
		when "0111100000111101" => data_out <= rom_array(30781);
		when "0111100000111110" => data_out <= rom_array(30782);
		when "0111100000111111" => data_out <= rom_array(30783);
		when "0111100001000000" => data_out <= rom_array(30784);
		when "0111100001000001" => data_out <= rom_array(30785);
		when "0111100001000010" => data_out <= rom_array(30786);
		when "0111100001000011" => data_out <= rom_array(30787);
		when "0111100001000100" => data_out <= rom_array(30788);
		when "0111100001000101" => data_out <= rom_array(30789);
		when "0111100001000110" => data_out <= rom_array(30790);
		when "0111100001000111" => data_out <= rom_array(30791);
		when "0111100001001000" => data_out <= rom_array(30792);
		when "0111100001001001" => data_out <= rom_array(30793);
		when "0111100001001010" => data_out <= rom_array(30794);
		when "0111100001001011" => data_out <= rom_array(30795);
		when "0111100001001100" => data_out <= rom_array(30796);
		when "0111100001001101" => data_out <= rom_array(30797);
		when "0111100001001110" => data_out <= rom_array(30798);
		when "0111100001001111" => data_out <= rom_array(30799);
		when "0111100001010000" => data_out <= rom_array(30800);
		when "0111100001010001" => data_out <= rom_array(30801);
		when "0111100001010010" => data_out <= rom_array(30802);
		when "0111100001010011" => data_out <= rom_array(30803);
		when "0111100001010100" => data_out <= rom_array(30804);
		when "0111100001010101" => data_out <= rom_array(30805);
		when "0111100001010110" => data_out <= rom_array(30806);
		when "0111100001010111" => data_out <= rom_array(30807);
		when "0111100001011000" => data_out <= rom_array(30808);
		when "0111100001011001" => data_out <= rom_array(30809);
		when "0111100001011010" => data_out <= rom_array(30810);
		when "0111100001011011" => data_out <= rom_array(30811);
		when "0111100001011100" => data_out <= rom_array(30812);
		when "0111100001011101" => data_out <= rom_array(30813);
		when "0111100001011110" => data_out <= rom_array(30814);
		when "0111100001011111" => data_out <= rom_array(30815);
		when "0111100001100000" => data_out <= rom_array(30816);
		when "0111100001100001" => data_out <= rom_array(30817);
		when "0111100001100010" => data_out <= rom_array(30818);
		when "0111100001100011" => data_out <= rom_array(30819);
		when "0111100001100100" => data_out <= rom_array(30820);
		when "0111100001100101" => data_out <= rom_array(30821);
		when "0111100001100110" => data_out <= rom_array(30822);
		when "0111100001100111" => data_out <= rom_array(30823);
		when "0111100001101000" => data_out <= rom_array(30824);
		when "0111100001101001" => data_out <= rom_array(30825);
		when "0111100001101010" => data_out <= rom_array(30826);
		when "0111100001101011" => data_out <= rom_array(30827);
		when "0111100001101100" => data_out <= rom_array(30828);
		when "0111100001101101" => data_out <= rom_array(30829);
		when "0111100001101110" => data_out <= rom_array(30830);
		when "0111100001101111" => data_out <= rom_array(30831);
		when "0111100001110000" => data_out <= rom_array(30832);
		when "0111100001110001" => data_out <= rom_array(30833);
		when "0111100001110010" => data_out <= rom_array(30834);
		when "0111100001110011" => data_out <= rom_array(30835);
		when "0111100001110100" => data_out <= rom_array(30836);
		when "0111100001110101" => data_out <= rom_array(30837);
		when "0111100001110110" => data_out <= rom_array(30838);
		when "0111100001110111" => data_out <= rom_array(30839);
		when "0111100001111000" => data_out <= rom_array(30840);
		when "0111100001111001" => data_out <= rom_array(30841);
		when "0111100001111010" => data_out <= rom_array(30842);
		when "0111100001111011" => data_out <= rom_array(30843);
		when "0111100001111100" => data_out <= rom_array(30844);
		when "0111100001111101" => data_out <= rom_array(30845);
		when "0111100001111110" => data_out <= rom_array(30846);
		when "0111100001111111" => data_out <= rom_array(30847);
		when "0111100010000000" => data_out <= rom_array(30848);
		when "0111100010000001" => data_out <= rom_array(30849);
		when "0111100010000010" => data_out <= rom_array(30850);
		when "0111100010000011" => data_out <= rom_array(30851);
		when "0111100010000100" => data_out <= rom_array(30852);
		when "0111100010000101" => data_out <= rom_array(30853);
		when "0111100010000110" => data_out <= rom_array(30854);
		when "0111100010000111" => data_out <= rom_array(30855);
		when "0111100010001000" => data_out <= rom_array(30856);
		when "0111100010001001" => data_out <= rom_array(30857);
		when "0111100010001010" => data_out <= rom_array(30858);
		when "0111100010001011" => data_out <= rom_array(30859);
		when "0111100010001100" => data_out <= rom_array(30860);
		when "0111100010001101" => data_out <= rom_array(30861);
		when "0111100010001110" => data_out <= rom_array(30862);
		when "0111100010001111" => data_out <= rom_array(30863);
		when "0111100010010000" => data_out <= rom_array(30864);
		when "0111100010010001" => data_out <= rom_array(30865);
		when "0111100010010010" => data_out <= rom_array(30866);
		when "0111100010010011" => data_out <= rom_array(30867);
		when "0111100010010100" => data_out <= rom_array(30868);
		when "0111100010010101" => data_out <= rom_array(30869);
		when "0111100010010110" => data_out <= rom_array(30870);
		when "0111100010010111" => data_out <= rom_array(30871);
		when "0111100010011000" => data_out <= rom_array(30872);
		when "0111100010011001" => data_out <= rom_array(30873);
		when "0111100010011010" => data_out <= rom_array(30874);
		when "0111100010011011" => data_out <= rom_array(30875);
		when "0111100010011100" => data_out <= rom_array(30876);
		when "0111100010011101" => data_out <= rom_array(30877);
		when "0111100010011110" => data_out <= rom_array(30878);
		when "0111100010011111" => data_out <= rom_array(30879);
		when "0111100010100000" => data_out <= rom_array(30880);
		when "0111100010100001" => data_out <= rom_array(30881);
		when "0111100010100010" => data_out <= rom_array(30882);
		when "0111100010100011" => data_out <= rom_array(30883);
		when "0111100010100100" => data_out <= rom_array(30884);
		when "0111100010100101" => data_out <= rom_array(30885);
		when "0111100010100110" => data_out <= rom_array(30886);
		when "0111100010100111" => data_out <= rom_array(30887);
		when "0111100010101000" => data_out <= rom_array(30888);
		when "0111100010101001" => data_out <= rom_array(30889);
		when "0111100010101010" => data_out <= rom_array(30890);
		when "0111100010101011" => data_out <= rom_array(30891);
		when "0111100010101100" => data_out <= rom_array(30892);
		when "0111100010101101" => data_out <= rom_array(30893);
		when "0111100010101110" => data_out <= rom_array(30894);
		when "0111100010101111" => data_out <= rom_array(30895);
		when "0111100010110000" => data_out <= rom_array(30896);
		when "0111100010110001" => data_out <= rom_array(30897);
		when "0111100010110010" => data_out <= rom_array(30898);
		when "0111100010110011" => data_out <= rom_array(30899);
		when "0111100010110100" => data_out <= rom_array(30900);
		when "0111100010110101" => data_out <= rom_array(30901);
		when "0111100010110110" => data_out <= rom_array(30902);
		when "0111100010110111" => data_out <= rom_array(30903);
		when "0111100010111000" => data_out <= rom_array(30904);
		when "0111100010111001" => data_out <= rom_array(30905);
		when "0111100010111010" => data_out <= rom_array(30906);
		when "0111100010111011" => data_out <= rom_array(30907);
		when "0111100010111100" => data_out <= rom_array(30908);
		when "0111100010111101" => data_out <= rom_array(30909);
		when "0111100010111110" => data_out <= rom_array(30910);
		when "0111100010111111" => data_out <= rom_array(30911);
		when "0111100011000000" => data_out <= rom_array(30912);
		when "0111100011000001" => data_out <= rom_array(30913);
		when "0111100011000010" => data_out <= rom_array(30914);
		when "0111100011000011" => data_out <= rom_array(30915);
		when "0111100011000100" => data_out <= rom_array(30916);
		when "0111100011000101" => data_out <= rom_array(30917);
		when "0111100011000110" => data_out <= rom_array(30918);
		when "0111100011000111" => data_out <= rom_array(30919);
		when "0111100011001000" => data_out <= rom_array(30920);
		when "0111100011001001" => data_out <= rom_array(30921);
		when "0111100011001010" => data_out <= rom_array(30922);
		when "0111100011001011" => data_out <= rom_array(30923);
		when "0111100011001100" => data_out <= rom_array(30924);
		when "0111100011001101" => data_out <= rom_array(30925);
		when "0111100011001110" => data_out <= rom_array(30926);
		when "0111100011001111" => data_out <= rom_array(30927);
		when "0111100011010000" => data_out <= rom_array(30928);
		when "0111100011010001" => data_out <= rom_array(30929);
		when "0111100011010010" => data_out <= rom_array(30930);
		when "0111100011010011" => data_out <= rom_array(30931);
		when "0111100011010100" => data_out <= rom_array(30932);
		when "0111100011010101" => data_out <= rom_array(30933);
		when "0111100011010110" => data_out <= rom_array(30934);
		when "0111100011010111" => data_out <= rom_array(30935);
		when "0111100011011000" => data_out <= rom_array(30936);
		when "0111100011011001" => data_out <= rom_array(30937);
		when "0111100011011010" => data_out <= rom_array(30938);
		when "0111100011011011" => data_out <= rom_array(30939);
		when "0111100011011100" => data_out <= rom_array(30940);
		when "0111100011011101" => data_out <= rom_array(30941);
		when "0111100011011110" => data_out <= rom_array(30942);
		when "0111100011011111" => data_out <= rom_array(30943);
		when "0111100011100000" => data_out <= rom_array(30944);
		when "0111100011100001" => data_out <= rom_array(30945);
		when "0111100011100010" => data_out <= rom_array(30946);
		when "0111100011100011" => data_out <= rom_array(30947);
		when "0111100011100100" => data_out <= rom_array(30948);
		when "0111100011100101" => data_out <= rom_array(30949);
		when "0111100011100110" => data_out <= rom_array(30950);
		when "0111100011100111" => data_out <= rom_array(30951);
		when "0111100011101000" => data_out <= rom_array(30952);
		when "0111100011101001" => data_out <= rom_array(30953);
		when "0111100011101010" => data_out <= rom_array(30954);
		when "0111100011101011" => data_out <= rom_array(30955);
		when "0111100011101100" => data_out <= rom_array(30956);
		when "0111100011101101" => data_out <= rom_array(30957);
		when "0111100011101110" => data_out <= rom_array(30958);
		when "0111100011101111" => data_out <= rom_array(30959);
		when "0111100011110000" => data_out <= rom_array(30960);
		when "0111100011110001" => data_out <= rom_array(30961);
		when "0111100011110010" => data_out <= rom_array(30962);
		when "0111100011110011" => data_out <= rom_array(30963);
		when "0111100011110100" => data_out <= rom_array(30964);
		when "0111100011110101" => data_out <= rom_array(30965);
		when "0111100011110110" => data_out <= rom_array(30966);
		when "0111100011110111" => data_out <= rom_array(30967);
		when "0111100011111000" => data_out <= rom_array(30968);
		when "0111100011111001" => data_out <= rom_array(30969);
		when "0111100011111010" => data_out <= rom_array(30970);
		when "0111100011111011" => data_out <= rom_array(30971);
		when "0111100011111100" => data_out <= rom_array(30972);
		when "0111100011111101" => data_out <= rom_array(30973);
		when "0111100011111110" => data_out <= rom_array(30974);
		when "0111100011111111" => data_out <= rom_array(30975);
		when "0111100100000000" => data_out <= rom_array(30976);
		when "0111100100000001" => data_out <= rom_array(30977);
		when "0111100100000010" => data_out <= rom_array(30978);
		when "0111100100000011" => data_out <= rom_array(30979);
		when "0111100100000100" => data_out <= rom_array(30980);
		when "0111100100000101" => data_out <= rom_array(30981);
		when "0111100100000110" => data_out <= rom_array(30982);
		when "0111100100000111" => data_out <= rom_array(30983);
		when "0111100100001000" => data_out <= rom_array(30984);
		when "0111100100001001" => data_out <= rom_array(30985);
		when "0111100100001010" => data_out <= rom_array(30986);
		when "0111100100001011" => data_out <= rom_array(30987);
		when "0111100100001100" => data_out <= rom_array(30988);
		when "0111100100001101" => data_out <= rom_array(30989);
		when "0111100100001110" => data_out <= rom_array(30990);
		when "0111100100001111" => data_out <= rom_array(30991);
		when "0111100100010000" => data_out <= rom_array(30992);
		when "0111100100010001" => data_out <= rom_array(30993);
		when "0111100100010010" => data_out <= rom_array(30994);
		when "0111100100010011" => data_out <= rom_array(30995);
		when "0111100100010100" => data_out <= rom_array(30996);
		when "0111100100010101" => data_out <= rom_array(30997);
		when "0111100100010110" => data_out <= rom_array(30998);
		when "0111100100010111" => data_out <= rom_array(30999);
		when "0111100100011000" => data_out <= rom_array(31000);
		when "0111100100011001" => data_out <= rom_array(31001);
		when "0111100100011010" => data_out <= rom_array(31002);
		when "0111100100011011" => data_out <= rom_array(31003);
		when "0111100100011100" => data_out <= rom_array(31004);
		when "0111100100011101" => data_out <= rom_array(31005);
		when "0111100100011110" => data_out <= rom_array(31006);
		when "0111100100011111" => data_out <= rom_array(31007);
		when "0111100100100000" => data_out <= rom_array(31008);
		when "0111100100100001" => data_out <= rom_array(31009);
		when "0111100100100010" => data_out <= rom_array(31010);
		when "0111100100100011" => data_out <= rom_array(31011);
		when "0111100100100100" => data_out <= rom_array(31012);
		when "0111100100100101" => data_out <= rom_array(31013);
		when "0111100100100110" => data_out <= rom_array(31014);
		when "0111100100100111" => data_out <= rom_array(31015);
		when "0111100100101000" => data_out <= rom_array(31016);
		when "0111100100101001" => data_out <= rom_array(31017);
		when "0111100100101010" => data_out <= rom_array(31018);
		when "0111100100101011" => data_out <= rom_array(31019);
		when "0111100100101100" => data_out <= rom_array(31020);
		when "0111100100101101" => data_out <= rom_array(31021);
		when "0111100100101110" => data_out <= rom_array(31022);
		when "0111100100101111" => data_out <= rom_array(31023);
		when "0111100100110000" => data_out <= rom_array(31024);
		when "0111100100110001" => data_out <= rom_array(31025);
		when "0111100100110010" => data_out <= rom_array(31026);
		when "0111100100110011" => data_out <= rom_array(31027);
		when "0111100100110100" => data_out <= rom_array(31028);
		when "0111100100110101" => data_out <= rom_array(31029);
		when "0111100100110110" => data_out <= rom_array(31030);
		when "0111100100110111" => data_out <= rom_array(31031);
		when "0111100100111000" => data_out <= rom_array(31032);
		when "0111100100111001" => data_out <= rom_array(31033);
		when "0111100100111010" => data_out <= rom_array(31034);
		when "0111100100111011" => data_out <= rom_array(31035);
		when "0111100100111100" => data_out <= rom_array(31036);
		when "0111100100111101" => data_out <= rom_array(31037);
		when "0111100100111110" => data_out <= rom_array(31038);
		when "0111100100111111" => data_out <= rom_array(31039);
		when "0111100101000000" => data_out <= rom_array(31040);
		when "0111100101000001" => data_out <= rom_array(31041);
		when "0111100101000010" => data_out <= rom_array(31042);
		when "0111100101000011" => data_out <= rom_array(31043);
		when "0111100101000100" => data_out <= rom_array(31044);
		when "0111100101000101" => data_out <= rom_array(31045);
		when "0111100101000110" => data_out <= rom_array(31046);
		when "0111100101000111" => data_out <= rom_array(31047);
		when "0111100101001000" => data_out <= rom_array(31048);
		when "0111100101001001" => data_out <= rom_array(31049);
		when "0111100101001010" => data_out <= rom_array(31050);
		when "0111100101001011" => data_out <= rom_array(31051);
		when "0111100101001100" => data_out <= rom_array(31052);
		when "0111100101001101" => data_out <= rom_array(31053);
		when "0111100101001110" => data_out <= rom_array(31054);
		when "0111100101001111" => data_out <= rom_array(31055);
		when "0111100101010000" => data_out <= rom_array(31056);
		when "0111100101010001" => data_out <= rom_array(31057);
		when "0111100101010010" => data_out <= rom_array(31058);
		when "0111100101010011" => data_out <= rom_array(31059);
		when "0111100101010100" => data_out <= rom_array(31060);
		when "0111100101010101" => data_out <= rom_array(31061);
		when "0111100101010110" => data_out <= rom_array(31062);
		when "0111100101010111" => data_out <= rom_array(31063);
		when "0111100101011000" => data_out <= rom_array(31064);
		when "0111100101011001" => data_out <= rom_array(31065);
		when "0111100101011010" => data_out <= rom_array(31066);
		when "0111100101011011" => data_out <= rom_array(31067);
		when "0111100101011100" => data_out <= rom_array(31068);
		when "0111100101011101" => data_out <= rom_array(31069);
		when "0111100101011110" => data_out <= rom_array(31070);
		when "0111100101011111" => data_out <= rom_array(31071);
		when "0111100101100000" => data_out <= rom_array(31072);
		when "0111100101100001" => data_out <= rom_array(31073);
		when "0111100101100010" => data_out <= rom_array(31074);
		when "0111100101100011" => data_out <= rom_array(31075);
		when "0111100101100100" => data_out <= rom_array(31076);
		when "0111100101100101" => data_out <= rom_array(31077);
		when "0111100101100110" => data_out <= rom_array(31078);
		when "0111100101100111" => data_out <= rom_array(31079);
		when "0111100101101000" => data_out <= rom_array(31080);
		when "0111100101101001" => data_out <= rom_array(31081);
		when "0111100101101010" => data_out <= rom_array(31082);
		when "0111100101101011" => data_out <= rom_array(31083);
		when "0111100101101100" => data_out <= rom_array(31084);
		when "0111100101101101" => data_out <= rom_array(31085);
		when "0111100101101110" => data_out <= rom_array(31086);
		when "0111100101101111" => data_out <= rom_array(31087);
		when "0111100101110000" => data_out <= rom_array(31088);
		when "0111100101110001" => data_out <= rom_array(31089);
		when "0111100101110010" => data_out <= rom_array(31090);
		when "0111100101110011" => data_out <= rom_array(31091);
		when "0111100101110100" => data_out <= rom_array(31092);
		when "0111100101110101" => data_out <= rom_array(31093);
		when "0111100101110110" => data_out <= rom_array(31094);
		when "0111100101110111" => data_out <= rom_array(31095);
		when "0111100101111000" => data_out <= rom_array(31096);
		when "0111100101111001" => data_out <= rom_array(31097);
		when "0111100101111010" => data_out <= rom_array(31098);
		when "0111100101111011" => data_out <= rom_array(31099);
		when "0111100101111100" => data_out <= rom_array(31100);
		when "0111100101111101" => data_out <= rom_array(31101);
		when "0111100101111110" => data_out <= rom_array(31102);
		when "0111100101111111" => data_out <= rom_array(31103);
		when "0111100110000000" => data_out <= rom_array(31104);
		when "0111100110000001" => data_out <= rom_array(31105);
		when "0111100110000010" => data_out <= rom_array(31106);
		when "0111100110000011" => data_out <= rom_array(31107);
		when "0111100110000100" => data_out <= rom_array(31108);
		when "0111100110000101" => data_out <= rom_array(31109);
		when "0111100110000110" => data_out <= rom_array(31110);
		when "0111100110000111" => data_out <= rom_array(31111);
		when "0111100110001000" => data_out <= rom_array(31112);
		when "0111100110001001" => data_out <= rom_array(31113);
		when "0111100110001010" => data_out <= rom_array(31114);
		when "0111100110001011" => data_out <= rom_array(31115);
		when "0111100110001100" => data_out <= rom_array(31116);
		when "0111100110001101" => data_out <= rom_array(31117);
		when "0111100110001110" => data_out <= rom_array(31118);
		when "0111100110001111" => data_out <= rom_array(31119);
		when "0111100110010000" => data_out <= rom_array(31120);
		when "0111100110010001" => data_out <= rom_array(31121);
		when "0111100110010010" => data_out <= rom_array(31122);
		when "0111100110010011" => data_out <= rom_array(31123);
		when "0111100110010100" => data_out <= rom_array(31124);
		when "0111100110010101" => data_out <= rom_array(31125);
		when "0111100110010110" => data_out <= rom_array(31126);
		when "0111100110010111" => data_out <= rom_array(31127);
		when "0111100110011000" => data_out <= rom_array(31128);
		when "0111100110011001" => data_out <= rom_array(31129);
		when "0111100110011010" => data_out <= rom_array(31130);
		when "0111100110011011" => data_out <= rom_array(31131);
		when "0111100110011100" => data_out <= rom_array(31132);
		when "0111100110011101" => data_out <= rom_array(31133);
		when "0111100110011110" => data_out <= rom_array(31134);
		when "0111100110011111" => data_out <= rom_array(31135);
		when "0111100110100000" => data_out <= rom_array(31136);
		when "0111100110100001" => data_out <= rom_array(31137);
		when "0111100110100010" => data_out <= rom_array(31138);
		when "0111100110100011" => data_out <= rom_array(31139);
		when "0111100110100100" => data_out <= rom_array(31140);
		when "0111100110100101" => data_out <= rom_array(31141);
		when "0111100110100110" => data_out <= rom_array(31142);
		when "0111100110100111" => data_out <= rom_array(31143);
		when "0111100110101000" => data_out <= rom_array(31144);
		when "0111100110101001" => data_out <= rom_array(31145);
		when "0111100110101010" => data_out <= rom_array(31146);
		when "0111100110101011" => data_out <= rom_array(31147);
		when "0111100110101100" => data_out <= rom_array(31148);
		when "0111100110101101" => data_out <= rom_array(31149);
		when "0111100110101110" => data_out <= rom_array(31150);
		when "0111100110101111" => data_out <= rom_array(31151);
		when "0111100110110000" => data_out <= rom_array(31152);
		when "0111100110110001" => data_out <= rom_array(31153);
		when "0111100110110010" => data_out <= rom_array(31154);
		when "0111100110110011" => data_out <= rom_array(31155);
		when "0111100110110100" => data_out <= rom_array(31156);
		when "0111100110110101" => data_out <= rom_array(31157);
		when "0111100110110110" => data_out <= rom_array(31158);
		when "0111100110110111" => data_out <= rom_array(31159);
		when "0111100110111000" => data_out <= rom_array(31160);
		when "0111100110111001" => data_out <= rom_array(31161);
		when "0111100110111010" => data_out <= rom_array(31162);
		when "0111100110111011" => data_out <= rom_array(31163);
		when "0111100110111100" => data_out <= rom_array(31164);
		when "0111100110111101" => data_out <= rom_array(31165);
		when "0111100110111110" => data_out <= rom_array(31166);
		when "0111100110111111" => data_out <= rom_array(31167);
		when "0111100111000000" => data_out <= rom_array(31168);
		when "0111100111000001" => data_out <= rom_array(31169);
		when "0111100111000010" => data_out <= rom_array(31170);
		when "0111100111000011" => data_out <= rom_array(31171);
		when "0111100111000100" => data_out <= rom_array(31172);
		when "0111100111000101" => data_out <= rom_array(31173);
		when "0111100111000110" => data_out <= rom_array(31174);
		when "0111100111000111" => data_out <= rom_array(31175);
		when "0111100111001000" => data_out <= rom_array(31176);
		when "0111100111001001" => data_out <= rom_array(31177);
		when "0111100111001010" => data_out <= rom_array(31178);
		when "0111100111001011" => data_out <= rom_array(31179);
		when "0111100111001100" => data_out <= rom_array(31180);
		when "0111100111001101" => data_out <= rom_array(31181);
		when "0111100111001110" => data_out <= rom_array(31182);
		when "0111100111001111" => data_out <= rom_array(31183);
		when "0111100111010000" => data_out <= rom_array(31184);
		when "0111100111010001" => data_out <= rom_array(31185);
		when "0111100111010010" => data_out <= rom_array(31186);
		when "0111100111010011" => data_out <= rom_array(31187);
		when "0111100111010100" => data_out <= rom_array(31188);
		when "0111100111010101" => data_out <= rom_array(31189);
		when "0111100111010110" => data_out <= rom_array(31190);
		when "0111100111010111" => data_out <= rom_array(31191);
		when "0111100111011000" => data_out <= rom_array(31192);
		when "0111100111011001" => data_out <= rom_array(31193);
		when "0111100111011010" => data_out <= rom_array(31194);
		when "0111100111011011" => data_out <= rom_array(31195);
		when "0111100111011100" => data_out <= rom_array(31196);
		when "0111100111011101" => data_out <= rom_array(31197);
		when "0111100111011110" => data_out <= rom_array(31198);
		when "0111100111011111" => data_out <= rom_array(31199);
		when "0111100111100000" => data_out <= rom_array(31200);
		when "0111100111100001" => data_out <= rom_array(31201);
		when "0111100111100010" => data_out <= rom_array(31202);
		when "0111100111100011" => data_out <= rom_array(31203);
		when "0111100111100100" => data_out <= rom_array(31204);
		when "0111100111100101" => data_out <= rom_array(31205);
		when "0111100111100110" => data_out <= rom_array(31206);
		when "0111100111100111" => data_out <= rom_array(31207);
		when "0111100111101000" => data_out <= rom_array(31208);
		when "0111100111101001" => data_out <= rom_array(31209);
		when "0111100111101010" => data_out <= rom_array(31210);
		when "0111100111101011" => data_out <= rom_array(31211);
		when "0111100111101100" => data_out <= rom_array(31212);
		when "0111100111101101" => data_out <= rom_array(31213);
		when "0111100111101110" => data_out <= rom_array(31214);
		when "0111100111101111" => data_out <= rom_array(31215);
		when "0111100111110000" => data_out <= rom_array(31216);
		when "0111100111110001" => data_out <= rom_array(31217);
		when "0111100111110010" => data_out <= rom_array(31218);
		when "0111100111110011" => data_out <= rom_array(31219);
		when "0111100111110100" => data_out <= rom_array(31220);
		when "0111100111110101" => data_out <= rom_array(31221);
		when "0111100111110110" => data_out <= rom_array(31222);
		when "0111100111110111" => data_out <= rom_array(31223);
		when "0111100111111000" => data_out <= rom_array(31224);
		when "0111100111111001" => data_out <= rom_array(31225);
		when "0111100111111010" => data_out <= rom_array(31226);
		when "0111100111111011" => data_out <= rom_array(31227);
		when "0111100111111100" => data_out <= rom_array(31228);
		when "0111100111111101" => data_out <= rom_array(31229);
		when "0111100111111110" => data_out <= rom_array(31230);
		when "0111100111111111" => data_out <= rom_array(31231);
		when "0111101000000000" => data_out <= rom_array(31232);
		when "0111101000000001" => data_out <= rom_array(31233);
		when "0111101000000010" => data_out <= rom_array(31234);
		when "0111101000000011" => data_out <= rom_array(31235);
		when "0111101000000100" => data_out <= rom_array(31236);
		when "0111101000000101" => data_out <= rom_array(31237);
		when "0111101000000110" => data_out <= rom_array(31238);
		when "0111101000000111" => data_out <= rom_array(31239);
		when "0111101000001000" => data_out <= rom_array(31240);
		when "0111101000001001" => data_out <= rom_array(31241);
		when "0111101000001010" => data_out <= rom_array(31242);
		when "0111101000001011" => data_out <= rom_array(31243);
		when "0111101000001100" => data_out <= rom_array(31244);
		when "0111101000001101" => data_out <= rom_array(31245);
		when "0111101000001110" => data_out <= rom_array(31246);
		when "0111101000001111" => data_out <= rom_array(31247);
		when "0111101000010000" => data_out <= rom_array(31248);
		when "0111101000010001" => data_out <= rom_array(31249);
		when "0111101000010010" => data_out <= rom_array(31250);
		when "0111101000010011" => data_out <= rom_array(31251);
		when "0111101000010100" => data_out <= rom_array(31252);
		when "0111101000010101" => data_out <= rom_array(31253);
		when "0111101000010110" => data_out <= rom_array(31254);
		when "0111101000010111" => data_out <= rom_array(31255);
		when "0111101000011000" => data_out <= rom_array(31256);
		when "0111101000011001" => data_out <= rom_array(31257);
		when "0111101000011010" => data_out <= rom_array(31258);
		when "0111101000011011" => data_out <= rom_array(31259);
		when "0111101000011100" => data_out <= rom_array(31260);
		when "0111101000011101" => data_out <= rom_array(31261);
		when "0111101000011110" => data_out <= rom_array(31262);
		when "0111101000011111" => data_out <= rom_array(31263);
		when "0111101000100000" => data_out <= rom_array(31264);
		when "0111101000100001" => data_out <= rom_array(31265);
		when "0111101000100010" => data_out <= rom_array(31266);
		when "0111101000100011" => data_out <= rom_array(31267);
		when "0111101000100100" => data_out <= rom_array(31268);
		when "0111101000100101" => data_out <= rom_array(31269);
		when "0111101000100110" => data_out <= rom_array(31270);
		when "0111101000100111" => data_out <= rom_array(31271);
		when "0111101000101000" => data_out <= rom_array(31272);
		when "0111101000101001" => data_out <= rom_array(31273);
		when "0111101000101010" => data_out <= rom_array(31274);
		when "0111101000101011" => data_out <= rom_array(31275);
		when "0111101000101100" => data_out <= rom_array(31276);
		when "0111101000101101" => data_out <= rom_array(31277);
		when "0111101000101110" => data_out <= rom_array(31278);
		when "0111101000101111" => data_out <= rom_array(31279);
		when "0111101000110000" => data_out <= rom_array(31280);
		when "0111101000110001" => data_out <= rom_array(31281);
		when "0111101000110010" => data_out <= rom_array(31282);
		when "0111101000110011" => data_out <= rom_array(31283);
		when "0111101000110100" => data_out <= rom_array(31284);
		when "0111101000110101" => data_out <= rom_array(31285);
		when "0111101000110110" => data_out <= rom_array(31286);
		when "0111101000110111" => data_out <= rom_array(31287);
		when "0111101000111000" => data_out <= rom_array(31288);
		when "0111101000111001" => data_out <= rom_array(31289);
		when "0111101000111010" => data_out <= rom_array(31290);
		when "0111101000111011" => data_out <= rom_array(31291);
		when "0111101000111100" => data_out <= rom_array(31292);
		when "0111101000111101" => data_out <= rom_array(31293);
		when "0111101000111110" => data_out <= rom_array(31294);
		when "0111101000111111" => data_out <= rom_array(31295);
		when "0111101001000000" => data_out <= rom_array(31296);
		when "0111101001000001" => data_out <= rom_array(31297);
		when "0111101001000010" => data_out <= rom_array(31298);
		when "0111101001000011" => data_out <= rom_array(31299);
		when "0111101001000100" => data_out <= rom_array(31300);
		when "0111101001000101" => data_out <= rom_array(31301);
		when "0111101001000110" => data_out <= rom_array(31302);
		when "0111101001000111" => data_out <= rom_array(31303);
		when "0111101001001000" => data_out <= rom_array(31304);
		when "0111101001001001" => data_out <= rom_array(31305);
		when "0111101001001010" => data_out <= rom_array(31306);
		when "0111101001001011" => data_out <= rom_array(31307);
		when "0111101001001100" => data_out <= rom_array(31308);
		when "0111101001001101" => data_out <= rom_array(31309);
		when "0111101001001110" => data_out <= rom_array(31310);
		when "0111101001001111" => data_out <= rom_array(31311);
		when "0111101001010000" => data_out <= rom_array(31312);
		when "0111101001010001" => data_out <= rom_array(31313);
		when "0111101001010010" => data_out <= rom_array(31314);
		when "0111101001010011" => data_out <= rom_array(31315);
		when "0111101001010100" => data_out <= rom_array(31316);
		when "0111101001010101" => data_out <= rom_array(31317);
		when "0111101001010110" => data_out <= rom_array(31318);
		when "0111101001010111" => data_out <= rom_array(31319);
		when "0111101001011000" => data_out <= rom_array(31320);
		when "0111101001011001" => data_out <= rom_array(31321);
		when "0111101001011010" => data_out <= rom_array(31322);
		when "0111101001011011" => data_out <= rom_array(31323);
		when "0111101001011100" => data_out <= rom_array(31324);
		when "0111101001011101" => data_out <= rom_array(31325);
		when "0111101001011110" => data_out <= rom_array(31326);
		when "0111101001011111" => data_out <= rom_array(31327);
		when "0111101001100000" => data_out <= rom_array(31328);
		when "0111101001100001" => data_out <= rom_array(31329);
		when "0111101001100010" => data_out <= rom_array(31330);
		when "0111101001100011" => data_out <= rom_array(31331);
		when "0111101001100100" => data_out <= rom_array(31332);
		when "0111101001100101" => data_out <= rom_array(31333);
		when "0111101001100110" => data_out <= rom_array(31334);
		when "0111101001100111" => data_out <= rom_array(31335);
		when "0111101001101000" => data_out <= rom_array(31336);
		when "0111101001101001" => data_out <= rom_array(31337);
		when "0111101001101010" => data_out <= rom_array(31338);
		when "0111101001101011" => data_out <= rom_array(31339);
		when "0111101001101100" => data_out <= rom_array(31340);
		when "0111101001101101" => data_out <= rom_array(31341);
		when "0111101001101110" => data_out <= rom_array(31342);
		when "0111101001101111" => data_out <= rom_array(31343);
		when "0111101001110000" => data_out <= rom_array(31344);
		when "0111101001110001" => data_out <= rom_array(31345);
		when "0111101001110010" => data_out <= rom_array(31346);
		when "0111101001110011" => data_out <= rom_array(31347);
		when "0111101001110100" => data_out <= rom_array(31348);
		when "0111101001110101" => data_out <= rom_array(31349);
		when "0111101001110110" => data_out <= rom_array(31350);
		when "0111101001110111" => data_out <= rom_array(31351);
		when "0111101001111000" => data_out <= rom_array(31352);
		when "0111101001111001" => data_out <= rom_array(31353);
		when "0111101001111010" => data_out <= rom_array(31354);
		when "0111101001111011" => data_out <= rom_array(31355);
		when "0111101001111100" => data_out <= rom_array(31356);
		when "0111101001111101" => data_out <= rom_array(31357);
		when "0111101001111110" => data_out <= rom_array(31358);
		when "0111101001111111" => data_out <= rom_array(31359);
		when "0111101010000000" => data_out <= rom_array(31360);
		when "0111101010000001" => data_out <= rom_array(31361);
		when "0111101010000010" => data_out <= rom_array(31362);
		when "0111101010000011" => data_out <= rom_array(31363);
		when "0111101010000100" => data_out <= rom_array(31364);
		when "0111101010000101" => data_out <= rom_array(31365);
		when "0111101010000110" => data_out <= rom_array(31366);
		when "0111101010000111" => data_out <= rom_array(31367);
		when "0111101010001000" => data_out <= rom_array(31368);
		when "0111101010001001" => data_out <= rom_array(31369);
		when "0111101010001010" => data_out <= rom_array(31370);
		when "0111101010001011" => data_out <= rom_array(31371);
		when "0111101010001100" => data_out <= rom_array(31372);
		when "0111101010001101" => data_out <= rom_array(31373);
		when "0111101010001110" => data_out <= rom_array(31374);
		when "0111101010001111" => data_out <= rom_array(31375);
		when "0111101010010000" => data_out <= rom_array(31376);
		when "0111101010010001" => data_out <= rom_array(31377);
		when "0111101010010010" => data_out <= rom_array(31378);
		when "0111101010010011" => data_out <= rom_array(31379);
		when "0111101010010100" => data_out <= rom_array(31380);
		when "0111101010010101" => data_out <= rom_array(31381);
		when "0111101010010110" => data_out <= rom_array(31382);
		when "0111101010010111" => data_out <= rom_array(31383);
		when "0111101010011000" => data_out <= rom_array(31384);
		when "0111101010011001" => data_out <= rom_array(31385);
		when "0111101010011010" => data_out <= rom_array(31386);
		when "0111101010011011" => data_out <= rom_array(31387);
		when "0111101010011100" => data_out <= rom_array(31388);
		when "0111101010011101" => data_out <= rom_array(31389);
		when "0111101010011110" => data_out <= rom_array(31390);
		when "0111101010011111" => data_out <= rom_array(31391);
		when "0111101010100000" => data_out <= rom_array(31392);
		when "0111101010100001" => data_out <= rom_array(31393);
		when "0111101010100010" => data_out <= rom_array(31394);
		when "0111101010100011" => data_out <= rom_array(31395);
		when "0111101010100100" => data_out <= rom_array(31396);
		when "0111101010100101" => data_out <= rom_array(31397);
		when "0111101010100110" => data_out <= rom_array(31398);
		when "0111101010100111" => data_out <= rom_array(31399);
		when "0111101010101000" => data_out <= rom_array(31400);
		when "0111101010101001" => data_out <= rom_array(31401);
		when "0111101010101010" => data_out <= rom_array(31402);
		when "0111101010101011" => data_out <= rom_array(31403);
		when "0111101010101100" => data_out <= rom_array(31404);
		when "0111101010101101" => data_out <= rom_array(31405);
		when "0111101010101110" => data_out <= rom_array(31406);
		when "0111101010101111" => data_out <= rom_array(31407);
		when "0111101010110000" => data_out <= rom_array(31408);
		when "0111101010110001" => data_out <= rom_array(31409);
		when "0111101010110010" => data_out <= rom_array(31410);
		when "0111101010110011" => data_out <= rom_array(31411);
		when "0111101010110100" => data_out <= rom_array(31412);
		when "0111101010110101" => data_out <= rom_array(31413);
		when "0111101010110110" => data_out <= rom_array(31414);
		when "0111101010110111" => data_out <= rom_array(31415);
		when "0111101010111000" => data_out <= rom_array(31416);
		when "0111101010111001" => data_out <= rom_array(31417);
		when "0111101010111010" => data_out <= rom_array(31418);
		when "0111101010111011" => data_out <= rom_array(31419);
		when "0111101010111100" => data_out <= rom_array(31420);
		when "0111101010111101" => data_out <= rom_array(31421);
		when "0111101010111110" => data_out <= rom_array(31422);
		when "0111101010111111" => data_out <= rom_array(31423);
		when "0111101011000000" => data_out <= rom_array(31424);
		when "0111101011000001" => data_out <= rom_array(31425);
		when "0111101011000010" => data_out <= rom_array(31426);
		when "0111101011000011" => data_out <= rom_array(31427);
		when "0111101011000100" => data_out <= rom_array(31428);
		when "0111101011000101" => data_out <= rom_array(31429);
		when "0111101011000110" => data_out <= rom_array(31430);
		when "0111101011000111" => data_out <= rom_array(31431);
		when "0111101011001000" => data_out <= rom_array(31432);
		when "0111101011001001" => data_out <= rom_array(31433);
		when "0111101011001010" => data_out <= rom_array(31434);
		when "0111101011001011" => data_out <= rom_array(31435);
		when "0111101011001100" => data_out <= rom_array(31436);
		when "0111101011001101" => data_out <= rom_array(31437);
		when "0111101011001110" => data_out <= rom_array(31438);
		when "0111101011001111" => data_out <= rom_array(31439);
		when "0111101011010000" => data_out <= rom_array(31440);
		when "0111101011010001" => data_out <= rom_array(31441);
		when "0111101011010010" => data_out <= rom_array(31442);
		when "0111101011010011" => data_out <= rom_array(31443);
		when "0111101011010100" => data_out <= rom_array(31444);
		when "0111101011010101" => data_out <= rom_array(31445);
		when "0111101011010110" => data_out <= rom_array(31446);
		when "0111101011010111" => data_out <= rom_array(31447);
		when "0111101011011000" => data_out <= rom_array(31448);
		when "0111101011011001" => data_out <= rom_array(31449);
		when "0111101011011010" => data_out <= rom_array(31450);
		when "0111101011011011" => data_out <= rom_array(31451);
		when "0111101011011100" => data_out <= rom_array(31452);
		when "0111101011011101" => data_out <= rom_array(31453);
		when "0111101011011110" => data_out <= rom_array(31454);
		when "0111101011011111" => data_out <= rom_array(31455);
		when "0111101011100000" => data_out <= rom_array(31456);
		when "0111101011100001" => data_out <= rom_array(31457);
		when "0111101011100010" => data_out <= rom_array(31458);
		when "0111101011100011" => data_out <= rom_array(31459);
		when "0111101011100100" => data_out <= rom_array(31460);
		when "0111101011100101" => data_out <= rom_array(31461);
		when "0111101011100110" => data_out <= rom_array(31462);
		when "0111101011100111" => data_out <= rom_array(31463);
		when "0111101011101000" => data_out <= rom_array(31464);
		when "0111101011101001" => data_out <= rom_array(31465);
		when "0111101011101010" => data_out <= rom_array(31466);
		when "0111101011101011" => data_out <= rom_array(31467);
		when "0111101011101100" => data_out <= rom_array(31468);
		when "0111101011101101" => data_out <= rom_array(31469);
		when "0111101011101110" => data_out <= rom_array(31470);
		when "0111101011101111" => data_out <= rom_array(31471);
		when "0111101011110000" => data_out <= rom_array(31472);
		when "0111101011110001" => data_out <= rom_array(31473);
		when "0111101011110010" => data_out <= rom_array(31474);
		when "0111101011110011" => data_out <= rom_array(31475);
		when "0111101011110100" => data_out <= rom_array(31476);
		when "0111101011110101" => data_out <= rom_array(31477);
		when "0111101011110110" => data_out <= rom_array(31478);
		when "0111101011110111" => data_out <= rom_array(31479);
		when "0111101011111000" => data_out <= rom_array(31480);
		when "0111101011111001" => data_out <= rom_array(31481);
		when "0111101011111010" => data_out <= rom_array(31482);
		when "0111101011111011" => data_out <= rom_array(31483);
		when "0111101011111100" => data_out <= rom_array(31484);
		when "0111101011111101" => data_out <= rom_array(31485);
		when "0111101011111110" => data_out <= rom_array(31486);
		when "0111101011111111" => data_out <= rom_array(31487);
		when "0111101100000000" => data_out <= rom_array(31488);
		when "0111101100000001" => data_out <= rom_array(31489);
		when "0111101100000010" => data_out <= rom_array(31490);
		when "0111101100000011" => data_out <= rom_array(31491);
		when "0111101100000100" => data_out <= rom_array(31492);
		when "0111101100000101" => data_out <= rom_array(31493);
		when "0111101100000110" => data_out <= rom_array(31494);
		when "0111101100000111" => data_out <= rom_array(31495);
		when "0111101100001000" => data_out <= rom_array(31496);
		when "0111101100001001" => data_out <= rom_array(31497);
		when "0111101100001010" => data_out <= rom_array(31498);
		when "0111101100001011" => data_out <= rom_array(31499);
		when "0111101100001100" => data_out <= rom_array(31500);
		when "0111101100001101" => data_out <= rom_array(31501);
		when "0111101100001110" => data_out <= rom_array(31502);
		when "0111101100001111" => data_out <= rom_array(31503);
		when "0111101100010000" => data_out <= rom_array(31504);
		when "0111101100010001" => data_out <= rom_array(31505);
		when "0111101100010010" => data_out <= rom_array(31506);
		when "0111101100010011" => data_out <= rom_array(31507);
		when "0111101100010100" => data_out <= rom_array(31508);
		when "0111101100010101" => data_out <= rom_array(31509);
		when "0111101100010110" => data_out <= rom_array(31510);
		when "0111101100010111" => data_out <= rom_array(31511);
		when "0111101100011000" => data_out <= rom_array(31512);
		when "0111101100011001" => data_out <= rom_array(31513);
		when "0111101100011010" => data_out <= rom_array(31514);
		when "0111101100011011" => data_out <= rom_array(31515);
		when "0111101100011100" => data_out <= rom_array(31516);
		when "0111101100011101" => data_out <= rom_array(31517);
		when "0111101100011110" => data_out <= rom_array(31518);
		when "0111101100011111" => data_out <= rom_array(31519);
		when "0111101100100000" => data_out <= rom_array(31520);
		when "0111101100100001" => data_out <= rom_array(31521);
		when "0111101100100010" => data_out <= rom_array(31522);
		when "0111101100100011" => data_out <= rom_array(31523);
		when "0111101100100100" => data_out <= rom_array(31524);
		when "0111101100100101" => data_out <= rom_array(31525);
		when "0111101100100110" => data_out <= rom_array(31526);
		when "0111101100100111" => data_out <= rom_array(31527);
		when "0111101100101000" => data_out <= rom_array(31528);
		when "0111101100101001" => data_out <= rom_array(31529);
		when "0111101100101010" => data_out <= rom_array(31530);
		when "0111101100101011" => data_out <= rom_array(31531);
		when "0111101100101100" => data_out <= rom_array(31532);
		when "0111101100101101" => data_out <= rom_array(31533);
		when "0111101100101110" => data_out <= rom_array(31534);
		when "0111101100101111" => data_out <= rom_array(31535);
		when "0111101100110000" => data_out <= rom_array(31536);
		when "0111101100110001" => data_out <= rom_array(31537);
		when "0111101100110010" => data_out <= rom_array(31538);
		when "0111101100110011" => data_out <= rom_array(31539);
		when "0111101100110100" => data_out <= rom_array(31540);
		when "0111101100110101" => data_out <= rom_array(31541);
		when "0111101100110110" => data_out <= rom_array(31542);
		when "0111101100110111" => data_out <= rom_array(31543);
		when "0111101100111000" => data_out <= rom_array(31544);
		when "0111101100111001" => data_out <= rom_array(31545);
		when "0111101100111010" => data_out <= rom_array(31546);
		when "0111101100111011" => data_out <= rom_array(31547);
		when "0111101100111100" => data_out <= rom_array(31548);
		when "0111101100111101" => data_out <= rom_array(31549);
		when "0111101100111110" => data_out <= rom_array(31550);
		when "0111101100111111" => data_out <= rom_array(31551);
		when "0111101101000000" => data_out <= rom_array(31552);
		when "0111101101000001" => data_out <= rom_array(31553);
		when "0111101101000010" => data_out <= rom_array(31554);
		when "0111101101000011" => data_out <= rom_array(31555);
		when "0111101101000100" => data_out <= rom_array(31556);
		when "0111101101000101" => data_out <= rom_array(31557);
		when "0111101101000110" => data_out <= rom_array(31558);
		when "0111101101000111" => data_out <= rom_array(31559);
		when "0111101101001000" => data_out <= rom_array(31560);
		when "0111101101001001" => data_out <= rom_array(31561);
		when "0111101101001010" => data_out <= rom_array(31562);
		when "0111101101001011" => data_out <= rom_array(31563);
		when "0111101101001100" => data_out <= rom_array(31564);
		when "0111101101001101" => data_out <= rom_array(31565);
		when "0111101101001110" => data_out <= rom_array(31566);
		when "0111101101001111" => data_out <= rom_array(31567);
		when "0111101101010000" => data_out <= rom_array(31568);
		when "0111101101010001" => data_out <= rom_array(31569);
		when "0111101101010010" => data_out <= rom_array(31570);
		when "0111101101010011" => data_out <= rom_array(31571);
		when "0111101101010100" => data_out <= rom_array(31572);
		when "0111101101010101" => data_out <= rom_array(31573);
		when "0111101101010110" => data_out <= rom_array(31574);
		when "0111101101010111" => data_out <= rom_array(31575);
		when "0111101101011000" => data_out <= rom_array(31576);
		when "0111101101011001" => data_out <= rom_array(31577);
		when "0111101101011010" => data_out <= rom_array(31578);
		when "0111101101011011" => data_out <= rom_array(31579);
		when "0111101101011100" => data_out <= rom_array(31580);
		when "0111101101011101" => data_out <= rom_array(31581);
		when "0111101101011110" => data_out <= rom_array(31582);
		when "0111101101011111" => data_out <= rom_array(31583);
		when "0111101101100000" => data_out <= rom_array(31584);
		when "0111101101100001" => data_out <= rom_array(31585);
		when "0111101101100010" => data_out <= rom_array(31586);
		when "0111101101100011" => data_out <= rom_array(31587);
		when "0111101101100100" => data_out <= rom_array(31588);
		when "0111101101100101" => data_out <= rom_array(31589);
		when "0111101101100110" => data_out <= rom_array(31590);
		when "0111101101100111" => data_out <= rom_array(31591);
		when "0111101101101000" => data_out <= rom_array(31592);
		when "0111101101101001" => data_out <= rom_array(31593);
		when "0111101101101010" => data_out <= rom_array(31594);
		when "0111101101101011" => data_out <= rom_array(31595);
		when "0111101101101100" => data_out <= rom_array(31596);
		when "0111101101101101" => data_out <= rom_array(31597);
		when "0111101101101110" => data_out <= rom_array(31598);
		when "0111101101101111" => data_out <= rom_array(31599);
		when "0111101101110000" => data_out <= rom_array(31600);
		when "0111101101110001" => data_out <= rom_array(31601);
		when "0111101101110010" => data_out <= rom_array(31602);
		when "0111101101110011" => data_out <= rom_array(31603);
		when "0111101101110100" => data_out <= rom_array(31604);
		when "0111101101110101" => data_out <= rom_array(31605);
		when "0111101101110110" => data_out <= rom_array(31606);
		when "0111101101110111" => data_out <= rom_array(31607);
		when "0111101101111000" => data_out <= rom_array(31608);
		when "0111101101111001" => data_out <= rom_array(31609);
		when "0111101101111010" => data_out <= rom_array(31610);
		when "0111101101111011" => data_out <= rom_array(31611);
		when "0111101101111100" => data_out <= rom_array(31612);
		when "0111101101111101" => data_out <= rom_array(31613);
		when "0111101101111110" => data_out <= rom_array(31614);
		when "0111101101111111" => data_out <= rom_array(31615);
		when "0111101110000000" => data_out <= rom_array(31616);
		when "0111101110000001" => data_out <= rom_array(31617);
		when "0111101110000010" => data_out <= rom_array(31618);
		when "0111101110000011" => data_out <= rom_array(31619);
		when "0111101110000100" => data_out <= rom_array(31620);
		when "0111101110000101" => data_out <= rom_array(31621);
		when "0111101110000110" => data_out <= rom_array(31622);
		when "0111101110000111" => data_out <= rom_array(31623);
		when "0111101110001000" => data_out <= rom_array(31624);
		when "0111101110001001" => data_out <= rom_array(31625);
		when "0111101110001010" => data_out <= rom_array(31626);
		when "0111101110001011" => data_out <= rom_array(31627);
		when "0111101110001100" => data_out <= rom_array(31628);
		when "0111101110001101" => data_out <= rom_array(31629);
		when "0111101110001110" => data_out <= rom_array(31630);
		when "0111101110001111" => data_out <= rom_array(31631);
		when "0111101110010000" => data_out <= rom_array(31632);
		when "0111101110010001" => data_out <= rom_array(31633);
		when "0111101110010010" => data_out <= rom_array(31634);
		when "0111101110010011" => data_out <= rom_array(31635);
		when "0111101110010100" => data_out <= rom_array(31636);
		when "0111101110010101" => data_out <= rom_array(31637);
		when "0111101110010110" => data_out <= rom_array(31638);
		when "0111101110010111" => data_out <= rom_array(31639);
		when "0111101110011000" => data_out <= rom_array(31640);
		when "0111101110011001" => data_out <= rom_array(31641);
		when "0111101110011010" => data_out <= rom_array(31642);
		when "0111101110011011" => data_out <= rom_array(31643);
		when "0111101110011100" => data_out <= rom_array(31644);
		when "0111101110011101" => data_out <= rom_array(31645);
		when "0111101110011110" => data_out <= rom_array(31646);
		when "0111101110011111" => data_out <= rom_array(31647);
		when "0111101110100000" => data_out <= rom_array(31648);
		when "0111101110100001" => data_out <= rom_array(31649);
		when "0111101110100010" => data_out <= rom_array(31650);
		when "0111101110100011" => data_out <= rom_array(31651);
		when "0111101110100100" => data_out <= rom_array(31652);
		when "0111101110100101" => data_out <= rom_array(31653);
		when "0111101110100110" => data_out <= rom_array(31654);
		when "0111101110100111" => data_out <= rom_array(31655);
		when "0111101110101000" => data_out <= rom_array(31656);
		when "0111101110101001" => data_out <= rom_array(31657);
		when "0111101110101010" => data_out <= rom_array(31658);
		when "0111101110101011" => data_out <= rom_array(31659);
		when "0111101110101100" => data_out <= rom_array(31660);
		when "0111101110101101" => data_out <= rom_array(31661);
		when "0111101110101110" => data_out <= rom_array(31662);
		when "0111101110101111" => data_out <= rom_array(31663);
		when "0111101110110000" => data_out <= rom_array(31664);
		when "0111101110110001" => data_out <= rom_array(31665);
		when "0111101110110010" => data_out <= rom_array(31666);
		when "0111101110110011" => data_out <= rom_array(31667);
		when "0111101110110100" => data_out <= rom_array(31668);
		when "0111101110110101" => data_out <= rom_array(31669);
		when "0111101110110110" => data_out <= rom_array(31670);
		when "0111101110110111" => data_out <= rom_array(31671);
		when "0111101110111000" => data_out <= rom_array(31672);
		when "0111101110111001" => data_out <= rom_array(31673);
		when "0111101110111010" => data_out <= rom_array(31674);
		when "0111101110111011" => data_out <= rom_array(31675);
		when "0111101110111100" => data_out <= rom_array(31676);
		when "0111101110111101" => data_out <= rom_array(31677);
		when "0111101110111110" => data_out <= rom_array(31678);
		when "0111101110111111" => data_out <= rom_array(31679);
		when "0111101111000000" => data_out <= rom_array(31680);
		when "0111101111000001" => data_out <= rom_array(31681);
		when "0111101111000010" => data_out <= rom_array(31682);
		when "0111101111000011" => data_out <= rom_array(31683);
		when "0111101111000100" => data_out <= rom_array(31684);
		when "0111101111000101" => data_out <= rom_array(31685);
		when "0111101111000110" => data_out <= rom_array(31686);
		when "0111101111000111" => data_out <= rom_array(31687);
		when "0111101111001000" => data_out <= rom_array(31688);
		when "0111101111001001" => data_out <= rom_array(31689);
		when "0111101111001010" => data_out <= rom_array(31690);
		when "0111101111001011" => data_out <= rom_array(31691);
		when "0111101111001100" => data_out <= rom_array(31692);
		when "0111101111001101" => data_out <= rom_array(31693);
		when "0111101111001110" => data_out <= rom_array(31694);
		when "0111101111001111" => data_out <= rom_array(31695);
		when "0111101111010000" => data_out <= rom_array(31696);
		when "0111101111010001" => data_out <= rom_array(31697);
		when "0111101111010010" => data_out <= rom_array(31698);
		when "0111101111010011" => data_out <= rom_array(31699);
		when "0111101111010100" => data_out <= rom_array(31700);
		when "0111101111010101" => data_out <= rom_array(31701);
		when "0111101111010110" => data_out <= rom_array(31702);
		when "0111101111010111" => data_out <= rom_array(31703);
		when "0111101111011000" => data_out <= rom_array(31704);
		when "0111101111011001" => data_out <= rom_array(31705);
		when "0111101111011010" => data_out <= rom_array(31706);
		when "0111101111011011" => data_out <= rom_array(31707);
		when "0111101111011100" => data_out <= rom_array(31708);
		when "0111101111011101" => data_out <= rom_array(31709);
		when "0111101111011110" => data_out <= rom_array(31710);
		when "0111101111011111" => data_out <= rom_array(31711);
		when "0111101111100000" => data_out <= rom_array(31712);
		when "0111101111100001" => data_out <= rom_array(31713);
		when "0111101111100010" => data_out <= rom_array(31714);
		when "0111101111100011" => data_out <= rom_array(31715);
		when "0111101111100100" => data_out <= rom_array(31716);
		when "0111101111100101" => data_out <= rom_array(31717);
		when "0111101111100110" => data_out <= rom_array(31718);
		when "0111101111100111" => data_out <= rom_array(31719);
		when "0111101111101000" => data_out <= rom_array(31720);
		when "0111101111101001" => data_out <= rom_array(31721);
		when "0111101111101010" => data_out <= rom_array(31722);
		when "0111101111101011" => data_out <= rom_array(31723);
		when "0111101111101100" => data_out <= rom_array(31724);
		when "0111101111101101" => data_out <= rom_array(31725);
		when "0111101111101110" => data_out <= rom_array(31726);
		when "0111101111101111" => data_out <= rom_array(31727);
		when "0111101111110000" => data_out <= rom_array(31728);
		when "0111101111110001" => data_out <= rom_array(31729);
		when "0111101111110010" => data_out <= rom_array(31730);
		when "0111101111110011" => data_out <= rom_array(31731);
		when "0111101111110100" => data_out <= rom_array(31732);
		when "0111101111110101" => data_out <= rom_array(31733);
		when "0111101111110110" => data_out <= rom_array(31734);
		when "0111101111110111" => data_out <= rom_array(31735);
		when "0111101111111000" => data_out <= rom_array(31736);
		when "0111101111111001" => data_out <= rom_array(31737);
		when "0111101111111010" => data_out <= rom_array(31738);
		when "0111101111111011" => data_out <= rom_array(31739);
		when "0111101111111100" => data_out <= rom_array(31740);
		when "0111101111111101" => data_out <= rom_array(31741);
		when "0111101111111110" => data_out <= rom_array(31742);
		when "0111101111111111" => data_out <= rom_array(31743);
		when "0111110000000000" => data_out <= rom_array(31744);
		when "0111110000000001" => data_out <= rom_array(31745);
		when "0111110000000010" => data_out <= rom_array(31746);
		when "0111110000000011" => data_out <= rom_array(31747);
		when "0111110000000100" => data_out <= rom_array(31748);
		when "0111110000000101" => data_out <= rom_array(31749);
		when "0111110000000110" => data_out <= rom_array(31750);
		when "0111110000000111" => data_out <= rom_array(31751);
		when "0111110000001000" => data_out <= rom_array(31752);
		when "0111110000001001" => data_out <= rom_array(31753);
		when "0111110000001010" => data_out <= rom_array(31754);
		when "0111110000001011" => data_out <= rom_array(31755);
		when "0111110000001100" => data_out <= rom_array(31756);
		when "0111110000001101" => data_out <= rom_array(31757);
		when "0111110000001110" => data_out <= rom_array(31758);
		when "0111110000001111" => data_out <= rom_array(31759);
		when "0111110000010000" => data_out <= rom_array(31760);
		when "0111110000010001" => data_out <= rom_array(31761);
		when "0111110000010010" => data_out <= rom_array(31762);
		when "0111110000010011" => data_out <= rom_array(31763);
		when "0111110000010100" => data_out <= rom_array(31764);
		when "0111110000010101" => data_out <= rom_array(31765);
		when "0111110000010110" => data_out <= rom_array(31766);
		when "0111110000010111" => data_out <= rom_array(31767);
		when "0111110000011000" => data_out <= rom_array(31768);
		when "0111110000011001" => data_out <= rom_array(31769);
		when "0111110000011010" => data_out <= rom_array(31770);
		when "0111110000011011" => data_out <= rom_array(31771);
		when "0111110000011100" => data_out <= rom_array(31772);
		when "0111110000011101" => data_out <= rom_array(31773);
		when "0111110000011110" => data_out <= rom_array(31774);
		when "0111110000011111" => data_out <= rom_array(31775);
		when "0111110000100000" => data_out <= rom_array(31776);
		when "0111110000100001" => data_out <= rom_array(31777);
		when "0111110000100010" => data_out <= rom_array(31778);
		when "0111110000100011" => data_out <= rom_array(31779);
		when "0111110000100100" => data_out <= rom_array(31780);
		when "0111110000100101" => data_out <= rom_array(31781);
		when "0111110000100110" => data_out <= rom_array(31782);
		when "0111110000100111" => data_out <= rom_array(31783);
		when "0111110000101000" => data_out <= rom_array(31784);
		when "0111110000101001" => data_out <= rom_array(31785);
		when "0111110000101010" => data_out <= rom_array(31786);
		when "0111110000101011" => data_out <= rom_array(31787);
		when "0111110000101100" => data_out <= rom_array(31788);
		when "0111110000101101" => data_out <= rom_array(31789);
		when "0111110000101110" => data_out <= rom_array(31790);
		when "0111110000101111" => data_out <= rom_array(31791);
		when "0111110000110000" => data_out <= rom_array(31792);
		when "0111110000110001" => data_out <= rom_array(31793);
		when "0111110000110010" => data_out <= rom_array(31794);
		when "0111110000110011" => data_out <= rom_array(31795);
		when "0111110000110100" => data_out <= rom_array(31796);
		when "0111110000110101" => data_out <= rom_array(31797);
		when "0111110000110110" => data_out <= rom_array(31798);
		when "0111110000110111" => data_out <= rom_array(31799);
		when "0111110000111000" => data_out <= rom_array(31800);
		when "0111110000111001" => data_out <= rom_array(31801);
		when "0111110000111010" => data_out <= rom_array(31802);
		when "0111110000111011" => data_out <= rom_array(31803);
		when "0111110000111100" => data_out <= rom_array(31804);
		when "0111110000111101" => data_out <= rom_array(31805);
		when "0111110000111110" => data_out <= rom_array(31806);
		when "0111110000111111" => data_out <= rom_array(31807);
		when "0111110001000000" => data_out <= rom_array(31808);
		when "0111110001000001" => data_out <= rom_array(31809);
		when "0111110001000010" => data_out <= rom_array(31810);
		when "0111110001000011" => data_out <= rom_array(31811);
		when "0111110001000100" => data_out <= rom_array(31812);
		when "0111110001000101" => data_out <= rom_array(31813);
		when "0111110001000110" => data_out <= rom_array(31814);
		when "0111110001000111" => data_out <= rom_array(31815);
		when "0111110001001000" => data_out <= rom_array(31816);
		when "0111110001001001" => data_out <= rom_array(31817);
		when "0111110001001010" => data_out <= rom_array(31818);
		when "0111110001001011" => data_out <= rom_array(31819);
		when "0111110001001100" => data_out <= rom_array(31820);
		when "0111110001001101" => data_out <= rom_array(31821);
		when "0111110001001110" => data_out <= rom_array(31822);
		when "0111110001001111" => data_out <= rom_array(31823);
		when "0111110001010000" => data_out <= rom_array(31824);
		when "0111110001010001" => data_out <= rom_array(31825);
		when "0111110001010010" => data_out <= rom_array(31826);
		when "0111110001010011" => data_out <= rom_array(31827);
		when "0111110001010100" => data_out <= rom_array(31828);
		when "0111110001010101" => data_out <= rom_array(31829);
		when "0111110001010110" => data_out <= rom_array(31830);
		when "0111110001010111" => data_out <= rom_array(31831);
		when "0111110001011000" => data_out <= rom_array(31832);
		when "0111110001011001" => data_out <= rom_array(31833);
		when "0111110001011010" => data_out <= rom_array(31834);
		when "0111110001011011" => data_out <= rom_array(31835);
		when "0111110001011100" => data_out <= rom_array(31836);
		when "0111110001011101" => data_out <= rom_array(31837);
		when "0111110001011110" => data_out <= rom_array(31838);
		when "0111110001011111" => data_out <= rom_array(31839);
		when "0111110001100000" => data_out <= rom_array(31840);
		when "0111110001100001" => data_out <= rom_array(31841);
		when "0111110001100010" => data_out <= rom_array(31842);
		when "0111110001100011" => data_out <= rom_array(31843);
		when "0111110001100100" => data_out <= rom_array(31844);
		when "0111110001100101" => data_out <= rom_array(31845);
		when "0111110001100110" => data_out <= rom_array(31846);
		when "0111110001100111" => data_out <= rom_array(31847);
		when "0111110001101000" => data_out <= rom_array(31848);
		when "0111110001101001" => data_out <= rom_array(31849);
		when "0111110001101010" => data_out <= rom_array(31850);
		when "0111110001101011" => data_out <= rom_array(31851);
		when "0111110001101100" => data_out <= rom_array(31852);
		when "0111110001101101" => data_out <= rom_array(31853);
		when "0111110001101110" => data_out <= rom_array(31854);
		when "0111110001101111" => data_out <= rom_array(31855);
		when "0111110001110000" => data_out <= rom_array(31856);
		when "0111110001110001" => data_out <= rom_array(31857);
		when "0111110001110010" => data_out <= rom_array(31858);
		when "0111110001110011" => data_out <= rom_array(31859);
		when "0111110001110100" => data_out <= rom_array(31860);
		when "0111110001110101" => data_out <= rom_array(31861);
		when "0111110001110110" => data_out <= rom_array(31862);
		when "0111110001110111" => data_out <= rom_array(31863);
		when "0111110001111000" => data_out <= rom_array(31864);
		when "0111110001111001" => data_out <= rom_array(31865);
		when "0111110001111010" => data_out <= rom_array(31866);
		when "0111110001111011" => data_out <= rom_array(31867);
		when "0111110001111100" => data_out <= rom_array(31868);
		when "0111110001111101" => data_out <= rom_array(31869);
		when "0111110001111110" => data_out <= rom_array(31870);
		when "0111110001111111" => data_out <= rom_array(31871);
		when "0111110010000000" => data_out <= rom_array(31872);
		when "0111110010000001" => data_out <= rom_array(31873);
		when "0111110010000010" => data_out <= rom_array(31874);
		when "0111110010000011" => data_out <= rom_array(31875);
		when "0111110010000100" => data_out <= rom_array(31876);
		when "0111110010000101" => data_out <= rom_array(31877);
		when "0111110010000110" => data_out <= rom_array(31878);
		when "0111110010000111" => data_out <= rom_array(31879);
		when "0111110010001000" => data_out <= rom_array(31880);
		when "0111110010001001" => data_out <= rom_array(31881);
		when "0111110010001010" => data_out <= rom_array(31882);
		when "0111110010001011" => data_out <= rom_array(31883);
		when "0111110010001100" => data_out <= rom_array(31884);
		when "0111110010001101" => data_out <= rom_array(31885);
		when "0111110010001110" => data_out <= rom_array(31886);
		when "0111110010001111" => data_out <= rom_array(31887);
		when "0111110010010000" => data_out <= rom_array(31888);
		when "0111110010010001" => data_out <= rom_array(31889);
		when "0111110010010010" => data_out <= rom_array(31890);
		when "0111110010010011" => data_out <= rom_array(31891);
		when "0111110010010100" => data_out <= rom_array(31892);
		when "0111110010010101" => data_out <= rom_array(31893);
		when "0111110010010110" => data_out <= rom_array(31894);
		when "0111110010010111" => data_out <= rom_array(31895);
		when "0111110010011000" => data_out <= rom_array(31896);
		when "0111110010011001" => data_out <= rom_array(31897);
		when "0111110010011010" => data_out <= rom_array(31898);
		when "0111110010011011" => data_out <= rom_array(31899);
		when "0111110010011100" => data_out <= rom_array(31900);
		when "0111110010011101" => data_out <= rom_array(31901);
		when "0111110010011110" => data_out <= rom_array(31902);
		when "0111110010011111" => data_out <= rom_array(31903);
		when "0111110010100000" => data_out <= rom_array(31904);
		when "0111110010100001" => data_out <= rom_array(31905);
		when "0111110010100010" => data_out <= rom_array(31906);
		when "0111110010100011" => data_out <= rom_array(31907);
		when "0111110010100100" => data_out <= rom_array(31908);
		when "0111110010100101" => data_out <= rom_array(31909);
		when "0111110010100110" => data_out <= rom_array(31910);
		when "0111110010100111" => data_out <= rom_array(31911);
		when "0111110010101000" => data_out <= rom_array(31912);
		when "0111110010101001" => data_out <= rom_array(31913);
		when "0111110010101010" => data_out <= rom_array(31914);
		when "0111110010101011" => data_out <= rom_array(31915);
		when "0111110010101100" => data_out <= rom_array(31916);
		when "0111110010101101" => data_out <= rom_array(31917);
		when "0111110010101110" => data_out <= rom_array(31918);
		when "0111110010101111" => data_out <= rom_array(31919);
		when "0111110010110000" => data_out <= rom_array(31920);
		when "0111110010110001" => data_out <= rom_array(31921);
		when "0111110010110010" => data_out <= rom_array(31922);
		when "0111110010110011" => data_out <= rom_array(31923);
		when "0111110010110100" => data_out <= rom_array(31924);
		when "0111110010110101" => data_out <= rom_array(31925);
		when "0111110010110110" => data_out <= rom_array(31926);
		when "0111110010110111" => data_out <= rom_array(31927);
		when "0111110010111000" => data_out <= rom_array(31928);
		when "0111110010111001" => data_out <= rom_array(31929);
		when "0111110010111010" => data_out <= rom_array(31930);
		when "0111110010111011" => data_out <= rom_array(31931);
		when "0111110010111100" => data_out <= rom_array(31932);
		when "0111110010111101" => data_out <= rom_array(31933);
		when "0111110010111110" => data_out <= rom_array(31934);
		when "0111110010111111" => data_out <= rom_array(31935);
		when "0111110011000000" => data_out <= rom_array(31936);
		when "0111110011000001" => data_out <= rom_array(31937);
		when "0111110011000010" => data_out <= rom_array(31938);
		when "0111110011000011" => data_out <= rom_array(31939);
		when "0111110011000100" => data_out <= rom_array(31940);
		when "0111110011000101" => data_out <= rom_array(31941);
		when "0111110011000110" => data_out <= rom_array(31942);
		when "0111110011000111" => data_out <= rom_array(31943);
		when "0111110011001000" => data_out <= rom_array(31944);
		when "0111110011001001" => data_out <= rom_array(31945);
		when "0111110011001010" => data_out <= rom_array(31946);
		when "0111110011001011" => data_out <= rom_array(31947);
		when "0111110011001100" => data_out <= rom_array(31948);
		when "0111110011001101" => data_out <= rom_array(31949);
		when "0111110011001110" => data_out <= rom_array(31950);
		when "0111110011001111" => data_out <= rom_array(31951);
		when "0111110011010000" => data_out <= rom_array(31952);
		when "0111110011010001" => data_out <= rom_array(31953);
		when "0111110011010010" => data_out <= rom_array(31954);
		when "0111110011010011" => data_out <= rom_array(31955);
		when "0111110011010100" => data_out <= rom_array(31956);
		when "0111110011010101" => data_out <= rom_array(31957);
		when "0111110011010110" => data_out <= rom_array(31958);
		when "0111110011010111" => data_out <= rom_array(31959);
		when "0111110011011000" => data_out <= rom_array(31960);
		when "0111110011011001" => data_out <= rom_array(31961);
		when "0111110011011010" => data_out <= rom_array(31962);
		when "0111110011011011" => data_out <= rom_array(31963);
		when "0111110011011100" => data_out <= rom_array(31964);
		when "0111110011011101" => data_out <= rom_array(31965);
		when "0111110011011110" => data_out <= rom_array(31966);
		when "0111110011011111" => data_out <= rom_array(31967);
		when "0111110011100000" => data_out <= rom_array(31968);
		when "0111110011100001" => data_out <= rom_array(31969);
		when "0111110011100010" => data_out <= rom_array(31970);
		when "0111110011100011" => data_out <= rom_array(31971);
		when "0111110011100100" => data_out <= rom_array(31972);
		when "0111110011100101" => data_out <= rom_array(31973);
		when "0111110011100110" => data_out <= rom_array(31974);
		when "0111110011100111" => data_out <= rom_array(31975);
		when "0111110011101000" => data_out <= rom_array(31976);
		when "0111110011101001" => data_out <= rom_array(31977);
		when "0111110011101010" => data_out <= rom_array(31978);
		when "0111110011101011" => data_out <= rom_array(31979);
		when "0111110011101100" => data_out <= rom_array(31980);
		when "0111110011101101" => data_out <= rom_array(31981);
		when "0111110011101110" => data_out <= rom_array(31982);
		when "0111110011101111" => data_out <= rom_array(31983);
		when "0111110011110000" => data_out <= rom_array(31984);
		when "0111110011110001" => data_out <= rom_array(31985);
		when "0111110011110010" => data_out <= rom_array(31986);
		when "0111110011110011" => data_out <= rom_array(31987);
		when "0111110011110100" => data_out <= rom_array(31988);
		when "0111110011110101" => data_out <= rom_array(31989);
		when "0111110011110110" => data_out <= rom_array(31990);
		when "0111110011110111" => data_out <= rom_array(31991);
		when "0111110011111000" => data_out <= rom_array(31992);
		when "0111110011111001" => data_out <= rom_array(31993);
		when "0111110011111010" => data_out <= rom_array(31994);
		when "0111110011111011" => data_out <= rom_array(31995);
		when "0111110011111100" => data_out <= rom_array(31996);
		when "0111110011111101" => data_out <= rom_array(31997);
		when "0111110011111110" => data_out <= rom_array(31998);
		when "0111110011111111" => data_out <= rom_array(31999);
		when "0111110100000000" => data_out <= rom_array(32000);
		when "0111110100000001" => data_out <= rom_array(32001);
		when "0111110100000010" => data_out <= rom_array(32002);
		when "0111110100000011" => data_out <= rom_array(32003);
		when "0111110100000100" => data_out <= rom_array(32004);
		when "0111110100000101" => data_out <= rom_array(32005);
		when "0111110100000110" => data_out <= rom_array(32006);
		when "0111110100000111" => data_out <= rom_array(32007);
		when "0111110100001000" => data_out <= rom_array(32008);
		when "0111110100001001" => data_out <= rom_array(32009);
		when "0111110100001010" => data_out <= rom_array(32010);
		when "0111110100001011" => data_out <= rom_array(32011);
		when "0111110100001100" => data_out <= rom_array(32012);
		when "0111110100001101" => data_out <= rom_array(32013);
		when "0111110100001110" => data_out <= rom_array(32014);
		when "0111110100001111" => data_out <= rom_array(32015);
		when "0111110100010000" => data_out <= rom_array(32016);
		when "0111110100010001" => data_out <= rom_array(32017);
		when "0111110100010010" => data_out <= rom_array(32018);
		when "0111110100010011" => data_out <= rom_array(32019);
		when "0111110100010100" => data_out <= rom_array(32020);
		when "0111110100010101" => data_out <= rom_array(32021);
		when "0111110100010110" => data_out <= rom_array(32022);
		when "0111110100010111" => data_out <= rom_array(32023);
		when "0111110100011000" => data_out <= rom_array(32024);
		when "0111110100011001" => data_out <= rom_array(32025);
		when "0111110100011010" => data_out <= rom_array(32026);
		when "0111110100011011" => data_out <= rom_array(32027);
		when "0111110100011100" => data_out <= rom_array(32028);
		when "0111110100011101" => data_out <= rom_array(32029);
		when "0111110100011110" => data_out <= rom_array(32030);
		when "0111110100011111" => data_out <= rom_array(32031);
		when "0111110100100000" => data_out <= rom_array(32032);
		when "0111110100100001" => data_out <= rom_array(32033);
		when "0111110100100010" => data_out <= rom_array(32034);
		when "0111110100100011" => data_out <= rom_array(32035);
		when "0111110100100100" => data_out <= rom_array(32036);
		when "0111110100100101" => data_out <= rom_array(32037);
		when "0111110100100110" => data_out <= rom_array(32038);
		when "0111110100100111" => data_out <= rom_array(32039);
		when "0111110100101000" => data_out <= rom_array(32040);
		when "0111110100101001" => data_out <= rom_array(32041);
		when "0111110100101010" => data_out <= rom_array(32042);
		when "0111110100101011" => data_out <= rom_array(32043);
		when "0111110100101100" => data_out <= rom_array(32044);
		when "0111110100101101" => data_out <= rom_array(32045);
		when "0111110100101110" => data_out <= rom_array(32046);
		when "0111110100101111" => data_out <= rom_array(32047);
		when "0111110100110000" => data_out <= rom_array(32048);
		when "0111110100110001" => data_out <= rom_array(32049);
		when "0111110100110010" => data_out <= rom_array(32050);
		when "0111110100110011" => data_out <= rom_array(32051);
		when "0111110100110100" => data_out <= rom_array(32052);
		when "0111110100110101" => data_out <= rom_array(32053);
		when "0111110100110110" => data_out <= rom_array(32054);
		when "0111110100110111" => data_out <= rom_array(32055);
		when "0111110100111000" => data_out <= rom_array(32056);
		when "0111110100111001" => data_out <= rom_array(32057);
		when "0111110100111010" => data_out <= rom_array(32058);
		when "0111110100111011" => data_out <= rom_array(32059);
		when "0111110100111100" => data_out <= rom_array(32060);
		when "0111110100111101" => data_out <= rom_array(32061);
		when "0111110100111110" => data_out <= rom_array(32062);
		when "0111110100111111" => data_out <= rom_array(32063);
		when "0111110101000000" => data_out <= rom_array(32064);
		when "0111110101000001" => data_out <= rom_array(32065);
		when "0111110101000010" => data_out <= rom_array(32066);
		when "0111110101000011" => data_out <= rom_array(32067);
		when "0111110101000100" => data_out <= rom_array(32068);
		when "0111110101000101" => data_out <= rom_array(32069);
		when "0111110101000110" => data_out <= rom_array(32070);
		when "0111110101000111" => data_out <= rom_array(32071);
		when "0111110101001000" => data_out <= rom_array(32072);
		when "0111110101001001" => data_out <= rom_array(32073);
		when "0111110101001010" => data_out <= rom_array(32074);
		when "0111110101001011" => data_out <= rom_array(32075);
		when "0111110101001100" => data_out <= rom_array(32076);
		when "0111110101001101" => data_out <= rom_array(32077);
		when "0111110101001110" => data_out <= rom_array(32078);
		when "0111110101001111" => data_out <= rom_array(32079);
		when "0111110101010000" => data_out <= rom_array(32080);
		when "0111110101010001" => data_out <= rom_array(32081);
		when "0111110101010010" => data_out <= rom_array(32082);
		when "0111110101010011" => data_out <= rom_array(32083);
		when "0111110101010100" => data_out <= rom_array(32084);
		when "0111110101010101" => data_out <= rom_array(32085);
		when "0111110101010110" => data_out <= rom_array(32086);
		when "0111110101010111" => data_out <= rom_array(32087);
		when "0111110101011000" => data_out <= rom_array(32088);
		when "0111110101011001" => data_out <= rom_array(32089);
		when "0111110101011010" => data_out <= rom_array(32090);
		when "0111110101011011" => data_out <= rom_array(32091);
		when "0111110101011100" => data_out <= rom_array(32092);
		when "0111110101011101" => data_out <= rom_array(32093);
		when "0111110101011110" => data_out <= rom_array(32094);
		when "0111110101011111" => data_out <= rom_array(32095);
		when "0111110101100000" => data_out <= rom_array(32096);
		when "0111110101100001" => data_out <= rom_array(32097);
		when "0111110101100010" => data_out <= rom_array(32098);
		when "0111110101100011" => data_out <= rom_array(32099);
		when "0111110101100100" => data_out <= rom_array(32100);
		when "0111110101100101" => data_out <= rom_array(32101);
		when "0111110101100110" => data_out <= rom_array(32102);
		when "0111110101100111" => data_out <= rom_array(32103);
		when "0111110101101000" => data_out <= rom_array(32104);
		when "0111110101101001" => data_out <= rom_array(32105);
		when "0111110101101010" => data_out <= rom_array(32106);
		when "0111110101101011" => data_out <= rom_array(32107);
		when "0111110101101100" => data_out <= rom_array(32108);
		when "0111110101101101" => data_out <= rom_array(32109);
		when "0111110101101110" => data_out <= rom_array(32110);
		when "0111110101101111" => data_out <= rom_array(32111);
		when "0111110101110000" => data_out <= rom_array(32112);
		when "0111110101110001" => data_out <= rom_array(32113);
		when "0111110101110010" => data_out <= rom_array(32114);
		when "0111110101110011" => data_out <= rom_array(32115);
		when "0111110101110100" => data_out <= rom_array(32116);
		when "0111110101110101" => data_out <= rom_array(32117);
		when "0111110101110110" => data_out <= rom_array(32118);
		when "0111110101110111" => data_out <= rom_array(32119);
		when "0111110101111000" => data_out <= rom_array(32120);
		when "0111110101111001" => data_out <= rom_array(32121);
		when "0111110101111010" => data_out <= rom_array(32122);
		when "0111110101111011" => data_out <= rom_array(32123);
		when "0111110101111100" => data_out <= rom_array(32124);
		when "0111110101111101" => data_out <= rom_array(32125);
		when "0111110101111110" => data_out <= rom_array(32126);
		when "0111110101111111" => data_out <= rom_array(32127);
		when "0111110110000000" => data_out <= rom_array(32128);
		when "0111110110000001" => data_out <= rom_array(32129);
		when "0111110110000010" => data_out <= rom_array(32130);
		when "0111110110000011" => data_out <= rom_array(32131);
		when "0111110110000100" => data_out <= rom_array(32132);
		when "0111110110000101" => data_out <= rom_array(32133);
		when "0111110110000110" => data_out <= rom_array(32134);
		when "0111110110000111" => data_out <= rom_array(32135);
		when "0111110110001000" => data_out <= rom_array(32136);
		when "0111110110001001" => data_out <= rom_array(32137);
		when "0111110110001010" => data_out <= rom_array(32138);
		when "0111110110001011" => data_out <= rom_array(32139);
		when "0111110110001100" => data_out <= rom_array(32140);
		when "0111110110001101" => data_out <= rom_array(32141);
		when "0111110110001110" => data_out <= rom_array(32142);
		when "0111110110001111" => data_out <= rom_array(32143);
		when "0111110110010000" => data_out <= rom_array(32144);
		when "0111110110010001" => data_out <= rom_array(32145);
		when "0111110110010010" => data_out <= rom_array(32146);
		when "0111110110010011" => data_out <= rom_array(32147);
		when "0111110110010100" => data_out <= rom_array(32148);
		when "0111110110010101" => data_out <= rom_array(32149);
		when "0111110110010110" => data_out <= rom_array(32150);
		when "0111110110010111" => data_out <= rom_array(32151);
		when "0111110110011000" => data_out <= rom_array(32152);
		when "0111110110011001" => data_out <= rom_array(32153);
		when "0111110110011010" => data_out <= rom_array(32154);
		when "0111110110011011" => data_out <= rom_array(32155);
		when "0111110110011100" => data_out <= rom_array(32156);
		when "0111110110011101" => data_out <= rom_array(32157);
		when "0111110110011110" => data_out <= rom_array(32158);
		when "0111110110011111" => data_out <= rom_array(32159);
		when "0111110110100000" => data_out <= rom_array(32160);
		when "0111110110100001" => data_out <= rom_array(32161);
		when "0111110110100010" => data_out <= rom_array(32162);
		when "0111110110100011" => data_out <= rom_array(32163);
		when "0111110110100100" => data_out <= rom_array(32164);
		when "0111110110100101" => data_out <= rom_array(32165);
		when "0111110110100110" => data_out <= rom_array(32166);
		when "0111110110100111" => data_out <= rom_array(32167);
		when "0111110110101000" => data_out <= rom_array(32168);
		when "0111110110101001" => data_out <= rom_array(32169);
		when "0111110110101010" => data_out <= rom_array(32170);
		when "0111110110101011" => data_out <= rom_array(32171);
		when "0111110110101100" => data_out <= rom_array(32172);
		when "0111110110101101" => data_out <= rom_array(32173);
		when "0111110110101110" => data_out <= rom_array(32174);
		when "0111110110101111" => data_out <= rom_array(32175);
		when "0111110110110000" => data_out <= rom_array(32176);
		when "0111110110110001" => data_out <= rom_array(32177);
		when "0111110110110010" => data_out <= rom_array(32178);
		when "0111110110110011" => data_out <= rom_array(32179);
		when "0111110110110100" => data_out <= rom_array(32180);
		when "0111110110110101" => data_out <= rom_array(32181);
		when "0111110110110110" => data_out <= rom_array(32182);
		when "0111110110110111" => data_out <= rom_array(32183);
		when "0111110110111000" => data_out <= rom_array(32184);
		when "0111110110111001" => data_out <= rom_array(32185);
		when "0111110110111010" => data_out <= rom_array(32186);
		when "0111110110111011" => data_out <= rom_array(32187);
		when "0111110110111100" => data_out <= rom_array(32188);
		when "0111110110111101" => data_out <= rom_array(32189);
		when "0111110110111110" => data_out <= rom_array(32190);
		when "0111110110111111" => data_out <= rom_array(32191);
		when "0111110111000000" => data_out <= rom_array(32192);
		when "0111110111000001" => data_out <= rom_array(32193);
		when "0111110111000010" => data_out <= rom_array(32194);
		when "0111110111000011" => data_out <= rom_array(32195);
		when "0111110111000100" => data_out <= rom_array(32196);
		when "0111110111000101" => data_out <= rom_array(32197);
		when "0111110111000110" => data_out <= rom_array(32198);
		when "0111110111000111" => data_out <= rom_array(32199);
		when "0111110111001000" => data_out <= rom_array(32200);
		when "0111110111001001" => data_out <= rom_array(32201);
		when "0111110111001010" => data_out <= rom_array(32202);
		when "0111110111001011" => data_out <= rom_array(32203);
		when "0111110111001100" => data_out <= rom_array(32204);
		when "0111110111001101" => data_out <= rom_array(32205);
		when "0111110111001110" => data_out <= rom_array(32206);
		when "0111110111001111" => data_out <= rom_array(32207);
		when "0111110111010000" => data_out <= rom_array(32208);
		when "0111110111010001" => data_out <= rom_array(32209);
		when "0111110111010010" => data_out <= rom_array(32210);
		when "0111110111010011" => data_out <= rom_array(32211);
		when "0111110111010100" => data_out <= rom_array(32212);
		when "0111110111010101" => data_out <= rom_array(32213);
		when "0111110111010110" => data_out <= rom_array(32214);
		when "0111110111010111" => data_out <= rom_array(32215);
		when "0111110111011000" => data_out <= rom_array(32216);
		when "0111110111011001" => data_out <= rom_array(32217);
		when "0111110111011010" => data_out <= rom_array(32218);
		when "0111110111011011" => data_out <= rom_array(32219);
		when "0111110111011100" => data_out <= rom_array(32220);
		when "0111110111011101" => data_out <= rom_array(32221);
		when "0111110111011110" => data_out <= rom_array(32222);
		when "0111110111011111" => data_out <= rom_array(32223);
		when "0111110111100000" => data_out <= rom_array(32224);
		when "0111110111100001" => data_out <= rom_array(32225);
		when "0111110111100010" => data_out <= rom_array(32226);
		when "0111110111100011" => data_out <= rom_array(32227);
		when "0111110111100100" => data_out <= rom_array(32228);
		when "0111110111100101" => data_out <= rom_array(32229);
		when "0111110111100110" => data_out <= rom_array(32230);
		when "0111110111100111" => data_out <= rom_array(32231);
		when "0111110111101000" => data_out <= rom_array(32232);
		when "0111110111101001" => data_out <= rom_array(32233);
		when "0111110111101010" => data_out <= rom_array(32234);
		when "0111110111101011" => data_out <= rom_array(32235);
		when "0111110111101100" => data_out <= rom_array(32236);
		when "0111110111101101" => data_out <= rom_array(32237);
		when "0111110111101110" => data_out <= rom_array(32238);
		when "0111110111101111" => data_out <= rom_array(32239);
		when "0111110111110000" => data_out <= rom_array(32240);
		when "0111110111110001" => data_out <= rom_array(32241);
		when "0111110111110010" => data_out <= rom_array(32242);
		when "0111110111110011" => data_out <= rom_array(32243);
		when "0111110111110100" => data_out <= rom_array(32244);
		when "0111110111110101" => data_out <= rom_array(32245);
		when "0111110111110110" => data_out <= rom_array(32246);
		when "0111110111110111" => data_out <= rom_array(32247);
		when "0111110111111000" => data_out <= rom_array(32248);
		when "0111110111111001" => data_out <= rom_array(32249);
		when "0111110111111010" => data_out <= rom_array(32250);
		when "0111110111111011" => data_out <= rom_array(32251);
		when "0111110111111100" => data_out <= rom_array(32252);
		when "0111110111111101" => data_out <= rom_array(32253);
		when "0111110111111110" => data_out <= rom_array(32254);
		when "0111110111111111" => data_out <= rom_array(32255);
		when "0111111000000000" => data_out <= rom_array(32256);
		when "0111111000000001" => data_out <= rom_array(32257);
		when "0111111000000010" => data_out <= rom_array(32258);
		when "0111111000000011" => data_out <= rom_array(32259);
		when "0111111000000100" => data_out <= rom_array(32260);
		when "0111111000000101" => data_out <= rom_array(32261);
		when "0111111000000110" => data_out <= rom_array(32262);
		when "0111111000000111" => data_out <= rom_array(32263);
		when "0111111000001000" => data_out <= rom_array(32264);
		when "0111111000001001" => data_out <= rom_array(32265);
		when "0111111000001010" => data_out <= rom_array(32266);
		when "0111111000001011" => data_out <= rom_array(32267);
		when "0111111000001100" => data_out <= rom_array(32268);
		when "0111111000001101" => data_out <= rom_array(32269);
		when "0111111000001110" => data_out <= rom_array(32270);
		when "0111111000001111" => data_out <= rom_array(32271);
		when "0111111000010000" => data_out <= rom_array(32272);
		when "0111111000010001" => data_out <= rom_array(32273);
		when "0111111000010010" => data_out <= rom_array(32274);
		when "0111111000010011" => data_out <= rom_array(32275);
		when "0111111000010100" => data_out <= rom_array(32276);
		when "0111111000010101" => data_out <= rom_array(32277);
		when "0111111000010110" => data_out <= rom_array(32278);
		when "0111111000010111" => data_out <= rom_array(32279);
		when "0111111000011000" => data_out <= rom_array(32280);
		when "0111111000011001" => data_out <= rom_array(32281);
		when "0111111000011010" => data_out <= rom_array(32282);
		when "0111111000011011" => data_out <= rom_array(32283);
		when "0111111000011100" => data_out <= rom_array(32284);
		when "0111111000011101" => data_out <= rom_array(32285);
		when "0111111000011110" => data_out <= rom_array(32286);
		when "0111111000011111" => data_out <= rom_array(32287);
		when "0111111000100000" => data_out <= rom_array(32288);
		when "0111111000100001" => data_out <= rom_array(32289);
		when "0111111000100010" => data_out <= rom_array(32290);
		when "0111111000100011" => data_out <= rom_array(32291);
		when "0111111000100100" => data_out <= rom_array(32292);
		when "0111111000100101" => data_out <= rom_array(32293);
		when "0111111000100110" => data_out <= rom_array(32294);
		when "0111111000100111" => data_out <= rom_array(32295);
		when "0111111000101000" => data_out <= rom_array(32296);
		when "0111111000101001" => data_out <= rom_array(32297);
		when "0111111000101010" => data_out <= rom_array(32298);
		when "0111111000101011" => data_out <= rom_array(32299);
		when "0111111000101100" => data_out <= rom_array(32300);
		when "0111111000101101" => data_out <= rom_array(32301);
		when "0111111000101110" => data_out <= rom_array(32302);
		when "0111111000101111" => data_out <= rom_array(32303);
		when "0111111000110000" => data_out <= rom_array(32304);
		when "0111111000110001" => data_out <= rom_array(32305);
		when "0111111000110010" => data_out <= rom_array(32306);
		when "0111111000110011" => data_out <= rom_array(32307);
		when "0111111000110100" => data_out <= rom_array(32308);
		when "0111111000110101" => data_out <= rom_array(32309);
		when "0111111000110110" => data_out <= rom_array(32310);
		when "0111111000110111" => data_out <= rom_array(32311);
		when "0111111000111000" => data_out <= rom_array(32312);
		when "0111111000111001" => data_out <= rom_array(32313);
		when "0111111000111010" => data_out <= rom_array(32314);
		when "0111111000111011" => data_out <= rom_array(32315);
		when "0111111000111100" => data_out <= rom_array(32316);
		when "0111111000111101" => data_out <= rom_array(32317);
		when "0111111000111110" => data_out <= rom_array(32318);
		when "0111111000111111" => data_out <= rom_array(32319);
		when "0111111001000000" => data_out <= rom_array(32320);
		when "0111111001000001" => data_out <= rom_array(32321);
		when "0111111001000010" => data_out <= rom_array(32322);
		when "0111111001000011" => data_out <= rom_array(32323);
		when "0111111001000100" => data_out <= rom_array(32324);
		when "0111111001000101" => data_out <= rom_array(32325);
		when "0111111001000110" => data_out <= rom_array(32326);
		when "0111111001000111" => data_out <= rom_array(32327);
		when "0111111001001000" => data_out <= rom_array(32328);
		when "0111111001001001" => data_out <= rom_array(32329);
		when "0111111001001010" => data_out <= rom_array(32330);
		when "0111111001001011" => data_out <= rom_array(32331);
		when "0111111001001100" => data_out <= rom_array(32332);
		when "0111111001001101" => data_out <= rom_array(32333);
		when "0111111001001110" => data_out <= rom_array(32334);
		when "0111111001001111" => data_out <= rom_array(32335);
		when "0111111001010000" => data_out <= rom_array(32336);
		when "0111111001010001" => data_out <= rom_array(32337);
		when "0111111001010010" => data_out <= rom_array(32338);
		when "0111111001010011" => data_out <= rom_array(32339);
		when "0111111001010100" => data_out <= rom_array(32340);
		when "0111111001010101" => data_out <= rom_array(32341);
		when "0111111001010110" => data_out <= rom_array(32342);
		when "0111111001010111" => data_out <= rom_array(32343);
		when "0111111001011000" => data_out <= rom_array(32344);
		when "0111111001011001" => data_out <= rom_array(32345);
		when "0111111001011010" => data_out <= rom_array(32346);
		when "0111111001011011" => data_out <= rom_array(32347);
		when "0111111001011100" => data_out <= rom_array(32348);
		when "0111111001011101" => data_out <= rom_array(32349);
		when "0111111001011110" => data_out <= rom_array(32350);
		when "0111111001011111" => data_out <= rom_array(32351);
		when "0111111001100000" => data_out <= rom_array(32352);
		when "0111111001100001" => data_out <= rom_array(32353);
		when "0111111001100010" => data_out <= rom_array(32354);
		when "0111111001100011" => data_out <= rom_array(32355);
		when "0111111001100100" => data_out <= rom_array(32356);
		when "0111111001100101" => data_out <= rom_array(32357);
		when "0111111001100110" => data_out <= rom_array(32358);
		when "0111111001100111" => data_out <= rom_array(32359);
		when "0111111001101000" => data_out <= rom_array(32360);
		when "0111111001101001" => data_out <= rom_array(32361);
		when "0111111001101010" => data_out <= rom_array(32362);
		when "0111111001101011" => data_out <= rom_array(32363);
		when "0111111001101100" => data_out <= rom_array(32364);
		when "0111111001101101" => data_out <= rom_array(32365);
		when "0111111001101110" => data_out <= rom_array(32366);
		when "0111111001101111" => data_out <= rom_array(32367);
		when "0111111001110000" => data_out <= rom_array(32368);
		when "0111111001110001" => data_out <= rom_array(32369);
		when "0111111001110010" => data_out <= rom_array(32370);
		when "0111111001110011" => data_out <= rom_array(32371);
		when "0111111001110100" => data_out <= rom_array(32372);
		when "0111111001110101" => data_out <= rom_array(32373);
		when "0111111001110110" => data_out <= rom_array(32374);
		when "0111111001110111" => data_out <= rom_array(32375);
		when "0111111001111000" => data_out <= rom_array(32376);
		when "0111111001111001" => data_out <= rom_array(32377);
		when "0111111001111010" => data_out <= rom_array(32378);
		when "0111111001111011" => data_out <= rom_array(32379);
		when "0111111001111100" => data_out <= rom_array(32380);
		when "0111111001111101" => data_out <= rom_array(32381);
		when "0111111001111110" => data_out <= rom_array(32382);
		when "0111111001111111" => data_out <= rom_array(32383);
		when "0111111010000000" => data_out <= rom_array(32384);
		when "0111111010000001" => data_out <= rom_array(32385);
		when "0111111010000010" => data_out <= rom_array(32386);
		when "0111111010000011" => data_out <= rom_array(32387);
		when "0111111010000100" => data_out <= rom_array(32388);
		when "0111111010000101" => data_out <= rom_array(32389);
		when "0111111010000110" => data_out <= rom_array(32390);
		when "0111111010000111" => data_out <= rom_array(32391);
		when "0111111010001000" => data_out <= rom_array(32392);
		when "0111111010001001" => data_out <= rom_array(32393);
		when "0111111010001010" => data_out <= rom_array(32394);
		when "0111111010001011" => data_out <= rom_array(32395);
		when "0111111010001100" => data_out <= rom_array(32396);
		when "0111111010001101" => data_out <= rom_array(32397);
		when "0111111010001110" => data_out <= rom_array(32398);
		when "0111111010001111" => data_out <= rom_array(32399);
		when "0111111010010000" => data_out <= rom_array(32400);
		when "0111111010010001" => data_out <= rom_array(32401);
		when "0111111010010010" => data_out <= rom_array(32402);
		when "0111111010010011" => data_out <= rom_array(32403);
		when "0111111010010100" => data_out <= rom_array(32404);
		when "0111111010010101" => data_out <= rom_array(32405);
		when "0111111010010110" => data_out <= rom_array(32406);
		when "0111111010010111" => data_out <= rom_array(32407);
		when "0111111010011000" => data_out <= rom_array(32408);
		when "0111111010011001" => data_out <= rom_array(32409);
		when "0111111010011010" => data_out <= rom_array(32410);
		when "0111111010011011" => data_out <= rom_array(32411);
		when "0111111010011100" => data_out <= rom_array(32412);
		when "0111111010011101" => data_out <= rom_array(32413);
		when "0111111010011110" => data_out <= rom_array(32414);
		when "0111111010011111" => data_out <= rom_array(32415);
		when "0111111010100000" => data_out <= rom_array(32416);
		when "0111111010100001" => data_out <= rom_array(32417);
		when "0111111010100010" => data_out <= rom_array(32418);
		when "0111111010100011" => data_out <= rom_array(32419);
		when "0111111010100100" => data_out <= rom_array(32420);
		when "0111111010100101" => data_out <= rom_array(32421);
		when "0111111010100110" => data_out <= rom_array(32422);
		when "0111111010100111" => data_out <= rom_array(32423);
		when "0111111010101000" => data_out <= rom_array(32424);
		when "0111111010101001" => data_out <= rom_array(32425);
		when "0111111010101010" => data_out <= rom_array(32426);
		when "0111111010101011" => data_out <= rom_array(32427);
		when "0111111010101100" => data_out <= rom_array(32428);
		when "0111111010101101" => data_out <= rom_array(32429);
		when "0111111010101110" => data_out <= rom_array(32430);
		when "0111111010101111" => data_out <= rom_array(32431);
		when "0111111010110000" => data_out <= rom_array(32432);
		when "0111111010110001" => data_out <= rom_array(32433);
		when "0111111010110010" => data_out <= rom_array(32434);
		when "0111111010110011" => data_out <= rom_array(32435);
		when "0111111010110100" => data_out <= rom_array(32436);
		when "0111111010110101" => data_out <= rom_array(32437);
		when "0111111010110110" => data_out <= rom_array(32438);
		when "0111111010110111" => data_out <= rom_array(32439);
		when "0111111010111000" => data_out <= rom_array(32440);
		when "0111111010111001" => data_out <= rom_array(32441);
		when "0111111010111010" => data_out <= rom_array(32442);
		when "0111111010111011" => data_out <= rom_array(32443);
		when "0111111010111100" => data_out <= rom_array(32444);
		when "0111111010111101" => data_out <= rom_array(32445);
		when "0111111010111110" => data_out <= rom_array(32446);
		when "0111111010111111" => data_out <= rom_array(32447);
		when "0111111011000000" => data_out <= rom_array(32448);
		when "0111111011000001" => data_out <= rom_array(32449);
		when "0111111011000010" => data_out <= rom_array(32450);
		when "0111111011000011" => data_out <= rom_array(32451);
		when "0111111011000100" => data_out <= rom_array(32452);
		when "0111111011000101" => data_out <= rom_array(32453);
		when "0111111011000110" => data_out <= rom_array(32454);
		when "0111111011000111" => data_out <= rom_array(32455);
		when "0111111011001000" => data_out <= rom_array(32456);
		when "0111111011001001" => data_out <= rom_array(32457);
		when "0111111011001010" => data_out <= rom_array(32458);
		when "0111111011001011" => data_out <= rom_array(32459);
		when "0111111011001100" => data_out <= rom_array(32460);
		when "0111111011001101" => data_out <= rom_array(32461);
		when "0111111011001110" => data_out <= rom_array(32462);
		when "0111111011001111" => data_out <= rom_array(32463);
		when "0111111011010000" => data_out <= rom_array(32464);
		when "0111111011010001" => data_out <= rom_array(32465);
		when "0111111011010010" => data_out <= rom_array(32466);
		when "0111111011010011" => data_out <= rom_array(32467);
		when "0111111011010100" => data_out <= rom_array(32468);
		when "0111111011010101" => data_out <= rom_array(32469);
		when "0111111011010110" => data_out <= rom_array(32470);
		when "0111111011010111" => data_out <= rom_array(32471);
		when "0111111011011000" => data_out <= rom_array(32472);
		when "0111111011011001" => data_out <= rom_array(32473);
		when "0111111011011010" => data_out <= rom_array(32474);
		when "0111111011011011" => data_out <= rom_array(32475);
		when "0111111011011100" => data_out <= rom_array(32476);
		when "0111111011011101" => data_out <= rom_array(32477);
		when "0111111011011110" => data_out <= rom_array(32478);
		when "0111111011011111" => data_out <= rom_array(32479);
		when "0111111011100000" => data_out <= rom_array(32480);
		when "0111111011100001" => data_out <= rom_array(32481);
		when "0111111011100010" => data_out <= rom_array(32482);
		when "0111111011100011" => data_out <= rom_array(32483);
		when "0111111011100100" => data_out <= rom_array(32484);
		when "0111111011100101" => data_out <= rom_array(32485);
		when "0111111011100110" => data_out <= rom_array(32486);
		when "0111111011100111" => data_out <= rom_array(32487);
		when "0111111011101000" => data_out <= rom_array(32488);
		when "0111111011101001" => data_out <= rom_array(32489);
		when "0111111011101010" => data_out <= rom_array(32490);
		when "0111111011101011" => data_out <= rom_array(32491);
		when "0111111011101100" => data_out <= rom_array(32492);
		when "0111111011101101" => data_out <= rom_array(32493);
		when "0111111011101110" => data_out <= rom_array(32494);
		when "0111111011101111" => data_out <= rom_array(32495);
		when "0111111011110000" => data_out <= rom_array(32496);
		when "0111111011110001" => data_out <= rom_array(32497);
		when "0111111011110010" => data_out <= rom_array(32498);
		when "0111111011110011" => data_out <= rom_array(32499);
		when "0111111011110100" => data_out <= rom_array(32500);
		when "0111111011110101" => data_out <= rom_array(32501);
		when "0111111011110110" => data_out <= rom_array(32502);
		when "0111111011110111" => data_out <= rom_array(32503);
		when "0111111011111000" => data_out <= rom_array(32504);
		when "0111111011111001" => data_out <= rom_array(32505);
		when "0111111011111010" => data_out <= rom_array(32506);
		when "0111111011111011" => data_out <= rom_array(32507);
		when "0111111011111100" => data_out <= rom_array(32508);
		when "0111111011111101" => data_out <= rom_array(32509);
		when "0111111011111110" => data_out <= rom_array(32510);
		when "0111111011111111" => data_out <= rom_array(32511);
		when "0111111100000000" => data_out <= rom_array(32512);
		when "0111111100000001" => data_out <= rom_array(32513);
		when "0111111100000010" => data_out <= rom_array(32514);
		when "0111111100000011" => data_out <= rom_array(32515);
		when "0111111100000100" => data_out <= rom_array(32516);
		when "0111111100000101" => data_out <= rom_array(32517);
		when "0111111100000110" => data_out <= rom_array(32518);
		when "0111111100000111" => data_out <= rom_array(32519);
		when "0111111100001000" => data_out <= rom_array(32520);
		when "0111111100001001" => data_out <= rom_array(32521);
		when "0111111100001010" => data_out <= rom_array(32522);
		when "0111111100001011" => data_out <= rom_array(32523);
		when "0111111100001100" => data_out <= rom_array(32524);
		when "0111111100001101" => data_out <= rom_array(32525);
		when "0111111100001110" => data_out <= rom_array(32526);
		when "0111111100001111" => data_out <= rom_array(32527);
		when "0111111100010000" => data_out <= rom_array(32528);
		when "0111111100010001" => data_out <= rom_array(32529);
		when "0111111100010010" => data_out <= rom_array(32530);
		when "0111111100010011" => data_out <= rom_array(32531);
		when "0111111100010100" => data_out <= rom_array(32532);
		when "0111111100010101" => data_out <= rom_array(32533);
		when "0111111100010110" => data_out <= rom_array(32534);
		when "0111111100010111" => data_out <= rom_array(32535);
		when "0111111100011000" => data_out <= rom_array(32536);
		when "0111111100011001" => data_out <= rom_array(32537);
		when "0111111100011010" => data_out <= rom_array(32538);
		when "0111111100011011" => data_out <= rom_array(32539);
		when "0111111100011100" => data_out <= rom_array(32540);
		when "0111111100011101" => data_out <= rom_array(32541);
		when "0111111100011110" => data_out <= rom_array(32542);
		when "0111111100011111" => data_out <= rom_array(32543);
		when "0111111100100000" => data_out <= rom_array(32544);
		when "0111111100100001" => data_out <= rom_array(32545);
		when "0111111100100010" => data_out <= rom_array(32546);
		when "0111111100100011" => data_out <= rom_array(32547);
		when "0111111100100100" => data_out <= rom_array(32548);
		when "0111111100100101" => data_out <= rom_array(32549);
		when "0111111100100110" => data_out <= rom_array(32550);
		when "0111111100100111" => data_out <= rom_array(32551);
		when "0111111100101000" => data_out <= rom_array(32552);
		when "0111111100101001" => data_out <= rom_array(32553);
		when "0111111100101010" => data_out <= rom_array(32554);
		when "0111111100101011" => data_out <= rom_array(32555);
		when "0111111100101100" => data_out <= rom_array(32556);
		when "0111111100101101" => data_out <= rom_array(32557);
		when "0111111100101110" => data_out <= rom_array(32558);
		when "0111111100101111" => data_out <= rom_array(32559);
		when "0111111100110000" => data_out <= rom_array(32560);
		when "0111111100110001" => data_out <= rom_array(32561);
		when "0111111100110010" => data_out <= rom_array(32562);
		when "0111111100110011" => data_out <= rom_array(32563);
		when "0111111100110100" => data_out <= rom_array(32564);
		when "0111111100110101" => data_out <= rom_array(32565);
		when "0111111100110110" => data_out <= rom_array(32566);
		when "0111111100110111" => data_out <= rom_array(32567);
		when "0111111100111000" => data_out <= rom_array(32568);
		when "0111111100111001" => data_out <= rom_array(32569);
		when "0111111100111010" => data_out <= rom_array(32570);
		when "0111111100111011" => data_out <= rom_array(32571);
		when "0111111100111100" => data_out <= rom_array(32572);
		when "0111111100111101" => data_out <= rom_array(32573);
		when "0111111100111110" => data_out <= rom_array(32574);
		when "0111111100111111" => data_out <= rom_array(32575);
		when "0111111101000000" => data_out <= rom_array(32576);
		when "0111111101000001" => data_out <= rom_array(32577);
		when "0111111101000010" => data_out <= rom_array(32578);
		when "0111111101000011" => data_out <= rom_array(32579);
		when "0111111101000100" => data_out <= rom_array(32580);
		when "0111111101000101" => data_out <= rom_array(32581);
		when "0111111101000110" => data_out <= rom_array(32582);
		when "0111111101000111" => data_out <= rom_array(32583);
		when "0111111101001000" => data_out <= rom_array(32584);
		when "0111111101001001" => data_out <= rom_array(32585);
		when "0111111101001010" => data_out <= rom_array(32586);
		when "0111111101001011" => data_out <= rom_array(32587);
		when "0111111101001100" => data_out <= rom_array(32588);
		when "0111111101001101" => data_out <= rom_array(32589);
		when "0111111101001110" => data_out <= rom_array(32590);
		when "0111111101001111" => data_out <= rom_array(32591);
		when "0111111101010000" => data_out <= rom_array(32592);
		when "0111111101010001" => data_out <= rom_array(32593);
		when "0111111101010010" => data_out <= rom_array(32594);
		when "0111111101010011" => data_out <= rom_array(32595);
		when "0111111101010100" => data_out <= rom_array(32596);
		when "0111111101010101" => data_out <= rom_array(32597);
		when "0111111101010110" => data_out <= rom_array(32598);
		when "0111111101010111" => data_out <= rom_array(32599);
		when "0111111101011000" => data_out <= rom_array(32600);
		when "0111111101011001" => data_out <= rom_array(32601);
		when "0111111101011010" => data_out <= rom_array(32602);
		when "0111111101011011" => data_out <= rom_array(32603);
		when "0111111101011100" => data_out <= rom_array(32604);
		when "0111111101011101" => data_out <= rom_array(32605);
		when "0111111101011110" => data_out <= rom_array(32606);
		when "0111111101011111" => data_out <= rom_array(32607);
		when "0111111101100000" => data_out <= rom_array(32608);
		when "0111111101100001" => data_out <= rom_array(32609);
		when "0111111101100010" => data_out <= rom_array(32610);
		when "0111111101100011" => data_out <= rom_array(32611);
		when "0111111101100100" => data_out <= rom_array(32612);
		when "0111111101100101" => data_out <= rom_array(32613);
		when "0111111101100110" => data_out <= rom_array(32614);
		when "0111111101100111" => data_out <= rom_array(32615);
		when "0111111101101000" => data_out <= rom_array(32616);
		when "0111111101101001" => data_out <= rom_array(32617);
		when "0111111101101010" => data_out <= rom_array(32618);
		when "0111111101101011" => data_out <= rom_array(32619);
		when "0111111101101100" => data_out <= rom_array(32620);
		when "0111111101101101" => data_out <= rom_array(32621);
		when "0111111101101110" => data_out <= rom_array(32622);
		when "0111111101101111" => data_out <= rom_array(32623);
		when "0111111101110000" => data_out <= rom_array(32624);
		when "0111111101110001" => data_out <= rom_array(32625);
		when "0111111101110010" => data_out <= rom_array(32626);
		when "0111111101110011" => data_out <= rom_array(32627);
		when "0111111101110100" => data_out <= rom_array(32628);
		when "0111111101110101" => data_out <= rom_array(32629);
		when "0111111101110110" => data_out <= rom_array(32630);
		when "0111111101110111" => data_out <= rom_array(32631);
		when "0111111101111000" => data_out <= rom_array(32632);
		when "0111111101111001" => data_out <= rom_array(32633);
		when "0111111101111010" => data_out <= rom_array(32634);
		when "0111111101111011" => data_out <= rom_array(32635);
		when "0111111101111100" => data_out <= rom_array(32636);
		when "0111111101111101" => data_out <= rom_array(32637);
		when "0111111101111110" => data_out <= rom_array(32638);
		when "0111111101111111" => data_out <= rom_array(32639);
		when "0111111110000000" => data_out <= rom_array(32640);
		when "0111111110000001" => data_out <= rom_array(32641);
		when "0111111110000010" => data_out <= rom_array(32642);
		when "0111111110000011" => data_out <= rom_array(32643);
		when "0111111110000100" => data_out <= rom_array(32644);
		when "0111111110000101" => data_out <= rom_array(32645);
		when "0111111110000110" => data_out <= rom_array(32646);
		when "0111111110000111" => data_out <= rom_array(32647);
		when "0111111110001000" => data_out <= rom_array(32648);
		when "0111111110001001" => data_out <= rom_array(32649);
		when "0111111110001010" => data_out <= rom_array(32650);
		when "0111111110001011" => data_out <= rom_array(32651);
		when "0111111110001100" => data_out <= rom_array(32652);
		when "0111111110001101" => data_out <= rom_array(32653);
		when "0111111110001110" => data_out <= rom_array(32654);
		when "0111111110001111" => data_out <= rom_array(32655);
		when "0111111110010000" => data_out <= rom_array(32656);
		when "0111111110010001" => data_out <= rom_array(32657);
		when "0111111110010010" => data_out <= rom_array(32658);
		when "0111111110010011" => data_out <= rom_array(32659);
		when "0111111110010100" => data_out <= rom_array(32660);
		when "0111111110010101" => data_out <= rom_array(32661);
		when "0111111110010110" => data_out <= rom_array(32662);
		when "0111111110010111" => data_out <= rom_array(32663);
		when "0111111110011000" => data_out <= rom_array(32664);
		when "0111111110011001" => data_out <= rom_array(32665);
		when "0111111110011010" => data_out <= rom_array(32666);
		when "0111111110011011" => data_out <= rom_array(32667);
		when "0111111110011100" => data_out <= rom_array(32668);
		when "0111111110011101" => data_out <= rom_array(32669);
		when "0111111110011110" => data_out <= rom_array(32670);
		when "0111111110011111" => data_out <= rom_array(32671);
		when "0111111110100000" => data_out <= rom_array(32672);
		when "0111111110100001" => data_out <= rom_array(32673);
		when "0111111110100010" => data_out <= rom_array(32674);
		when "0111111110100011" => data_out <= rom_array(32675);
		when "0111111110100100" => data_out <= rom_array(32676);
		when "0111111110100101" => data_out <= rom_array(32677);
		when "0111111110100110" => data_out <= rom_array(32678);
		when "0111111110100111" => data_out <= rom_array(32679);
		when "0111111110101000" => data_out <= rom_array(32680);
		when "0111111110101001" => data_out <= rom_array(32681);
		when "0111111110101010" => data_out <= rom_array(32682);
		when "0111111110101011" => data_out <= rom_array(32683);
		when "0111111110101100" => data_out <= rom_array(32684);
		when "0111111110101101" => data_out <= rom_array(32685);
		when "0111111110101110" => data_out <= rom_array(32686);
		when "0111111110101111" => data_out <= rom_array(32687);
		when "0111111110110000" => data_out <= rom_array(32688);
		when "0111111110110001" => data_out <= rom_array(32689);
		when "0111111110110010" => data_out <= rom_array(32690);
		when "0111111110110011" => data_out <= rom_array(32691);
		when "0111111110110100" => data_out <= rom_array(32692);
		when "0111111110110101" => data_out <= rom_array(32693);
		when "0111111110110110" => data_out <= rom_array(32694);
		when "0111111110110111" => data_out <= rom_array(32695);
		when "0111111110111000" => data_out <= rom_array(32696);
		when "0111111110111001" => data_out <= rom_array(32697);
		when "0111111110111010" => data_out <= rom_array(32698);
		when "0111111110111011" => data_out <= rom_array(32699);
		when "0111111110111100" => data_out <= rom_array(32700);
		when "0111111110111101" => data_out <= rom_array(32701);
		when "0111111110111110" => data_out <= rom_array(32702);
		when "0111111110111111" => data_out <= rom_array(32703);
		when "0111111111000000" => data_out <= rom_array(32704);
		when "0111111111000001" => data_out <= rom_array(32705);
		when "0111111111000010" => data_out <= rom_array(32706);
		when "0111111111000011" => data_out <= rom_array(32707);
		when "0111111111000100" => data_out <= rom_array(32708);
		when "0111111111000101" => data_out <= rom_array(32709);
		when "0111111111000110" => data_out <= rom_array(32710);
		when "0111111111000111" => data_out <= rom_array(32711);
		when "0111111111001000" => data_out <= rom_array(32712);
		when "0111111111001001" => data_out <= rom_array(32713);
		when "0111111111001010" => data_out <= rom_array(32714);
		when "0111111111001011" => data_out <= rom_array(32715);
		when "0111111111001100" => data_out <= rom_array(32716);
		when "0111111111001101" => data_out <= rom_array(32717);
		when "0111111111001110" => data_out <= rom_array(32718);
		when "0111111111001111" => data_out <= rom_array(32719);
		when "0111111111010000" => data_out <= rom_array(32720);
		when "0111111111010001" => data_out <= rom_array(32721);
		when "0111111111010010" => data_out <= rom_array(32722);
		when "0111111111010011" => data_out <= rom_array(32723);
		when "0111111111010100" => data_out <= rom_array(32724);
		when "0111111111010101" => data_out <= rom_array(32725);
		when "0111111111010110" => data_out <= rom_array(32726);
		when "0111111111010111" => data_out <= rom_array(32727);
		when "0111111111011000" => data_out <= rom_array(32728);
		when "0111111111011001" => data_out <= rom_array(32729);
		when "0111111111011010" => data_out <= rom_array(32730);
		when "0111111111011011" => data_out <= rom_array(32731);
		when "0111111111011100" => data_out <= rom_array(32732);
		when "0111111111011101" => data_out <= rom_array(32733);
		when "0111111111011110" => data_out <= rom_array(32734);
		when "0111111111011111" => data_out <= rom_array(32735);
		when "0111111111100000" => data_out <= rom_array(32736);
		when "0111111111100001" => data_out <= rom_array(32737);
		when "0111111111100010" => data_out <= rom_array(32738);
		when "0111111111100011" => data_out <= rom_array(32739);
		when "0111111111100100" => data_out <= rom_array(32740);
		when "0111111111100101" => data_out <= rom_array(32741);
		when "0111111111100110" => data_out <= rom_array(32742);
		when "0111111111100111" => data_out <= rom_array(32743);
		when "0111111111101000" => data_out <= rom_array(32744);
		when "0111111111101001" => data_out <= rom_array(32745);
		when "0111111111101010" => data_out <= rom_array(32746);
		when "0111111111101011" => data_out <= rom_array(32747);
		when "0111111111101100" => data_out <= rom_array(32748);
		when "0111111111101101" => data_out <= rom_array(32749);
		when "0111111111101110" => data_out <= rom_array(32750);
		when "0111111111101111" => data_out <= rom_array(32751);
		when "0111111111110000" => data_out <= rom_array(32752);
		when "0111111111110001" => data_out <= rom_array(32753);
		when "0111111111110010" => data_out <= rom_array(32754);
		when "0111111111110011" => data_out <= rom_array(32755);
		when "0111111111110100" => data_out <= rom_array(32756);
		when "0111111111110101" => data_out <= rom_array(32757);
		when "0111111111110110" => data_out <= rom_array(32758);
		when "0111111111110111" => data_out <= rom_array(32759);
		when "0111111111111000" => data_out <= rom_array(32760);
		when "0111111111111001" => data_out <= rom_array(32761);
		when "0111111111111010" => data_out <= rom_array(32762);
		when "0111111111111011" => data_out <= rom_array(32763);
		when "0111111111111100" => data_out <= rom_array(32764);
		when "0111111111111101" => data_out <= rom_array(32765);
		when "0111111111111110" => data_out <= rom_array(32766);
		when "0111111111111111" => data_out <= rom_array(32767);
		when "1000000000000000" => data_out <= rom_array(32768);
		when "1000000000000001" => data_out <= rom_array(32769);
		when "1000000000000010" => data_out <= rom_array(32770);
		when "1000000000000011" => data_out <= rom_array(32771);
		when "1000000000000100" => data_out <= rom_array(32772);
		when "1000000000000101" => data_out <= rom_array(32773);
		when "1000000000000110" => data_out <= rom_array(32774);
		when "1000000000000111" => data_out <= rom_array(32775);
		when "1000000000001000" => data_out <= rom_array(32776);
		when "1000000000001001" => data_out <= rom_array(32777);
		when "1000000000001010" => data_out <= rom_array(32778);
		when "1000000000001011" => data_out <= rom_array(32779);
		when "1000000000001100" => data_out <= rom_array(32780);
		when "1000000000001101" => data_out <= rom_array(32781);
		when "1000000000001110" => data_out <= rom_array(32782);
		when "1000000000001111" => data_out <= rom_array(32783);
		when "1000000000010000" => data_out <= rom_array(32784);
		when "1000000000010001" => data_out <= rom_array(32785);
		when "1000000000010010" => data_out <= rom_array(32786);
		when "1000000000010011" => data_out <= rom_array(32787);
		when "1000000000010100" => data_out <= rom_array(32788);
		when "1000000000010101" => data_out <= rom_array(32789);
		when "1000000000010110" => data_out <= rom_array(32790);
		when "1000000000010111" => data_out <= rom_array(32791);
		when "1000000000011000" => data_out <= rom_array(32792);
		when "1000000000011001" => data_out <= rom_array(32793);
		when "1000000000011010" => data_out <= rom_array(32794);
		when "1000000000011011" => data_out <= rom_array(32795);
		when "1000000000011100" => data_out <= rom_array(32796);
		when "1000000000011101" => data_out <= rom_array(32797);
		when "1000000000011110" => data_out <= rom_array(32798);
		when "1000000000011111" => data_out <= rom_array(32799);
		when "1000000000100000" => data_out <= rom_array(32800);
		when "1000000000100001" => data_out <= rom_array(32801);
		when "1000000000100010" => data_out <= rom_array(32802);
		when "1000000000100011" => data_out <= rom_array(32803);
		when "1000000000100100" => data_out <= rom_array(32804);
		when "1000000000100101" => data_out <= rom_array(32805);
		when "1000000000100110" => data_out <= rom_array(32806);
		when "1000000000100111" => data_out <= rom_array(32807);
		when "1000000000101000" => data_out <= rom_array(32808);
		when "1000000000101001" => data_out <= rom_array(32809);
		when "1000000000101010" => data_out <= rom_array(32810);
		when "1000000000101011" => data_out <= rom_array(32811);
		when "1000000000101100" => data_out <= rom_array(32812);
		when "1000000000101101" => data_out <= rom_array(32813);
		when "1000000000101110" => data_out <= rom_array(32814);
		when "1000000000101111" => data_out <= rom_array(32815);
		when "1000000000110000" => data_out <= rom_array(32816);
		when "1000000000110001" => data_out <= rom_array(32817);
		when "1000000000110010" => data_out <= rom_array(32818);
		when "1000000000110011" => data_out <= rom_array(32819);
		when "1000000000110100" => data_out <= rom_array(32820);
		when "1000000000110101" => data_out <= rom_array(32821);
		when "1000000000110110" => data_out <= rom_array(32822);
		when "1000000000110111" => data_out <= rom_array(32823);
		when "1000000000111000" => data_out <= rom_array(32824);
		when "1000000000111001" => data_out <= rom_array(32825);
		when "1000000000111010" => data_out <= rom_array(32826);
		when "1000000000111011" => data_out <= rom_array(32827);
		when "1000000000111100" => data_out <= rom_array(32828);
		when "1000000000111101" => data_out <= rom_array(32829);
		when "1000000000111110" => data_out <= rom_array(32830);
		when "1000000000111111" => data_out <= rom_array(32831);
		when "1000000001000000" => data_out <= rom_array(32832);
		when "1000000001000001" => data_out <= rom_array(32833);
		when "1000000001000010" => data_out <= rom_array(32834);
		when "1000000001000011" => data_out <= rom_array(32835);
		when "1000000001000100" => data_out <= rom_array(32836);
		when "1000000001000101" => data_out <= rom_array(32837);
		when "1000000001000110" => data_out <= rom_array(32838);
		when "1000000001000111" => data_out <= rom_array(32839);
		when "1000000001001000" => data_out <= rom_array(32840);
		when "1000000001001001" => data_out <= rom_array(32841);
		when "1000000001001010" => data_out <= rom_array(32842);
		when "1000000001001011" => data_out <= rom_array(32843);
		when "1000000001001100" => data_out <= rom_array(32844);
		when "1000000001001101" => data_out <= rom_array(32845);
		when "1000000001001110" => data_out <= rom_array(32846);
		when "1000000001001111" => data_out <= rom_array(32847);
		when "1000000001010000" => data_out <= rom_array(32848);
		when "1000000001010001" => data_out <= rom_array(32849);
		when "1000000001010010" => data_out <= rom_array(32850);
		when "1000000001010011" => data_out <= rom_array(32851);
		when "1000000001010100" => data_out <= rom_array(32852);
		when "1000000001010101" => data_out <= rom_array(32853);
		when "1000000001010110" => data_out <= rom_array(32854);
		when "1000000001010111" => data_out <= rom_array(32855);
		when "1000000001011000" => data_out <= rom_array(32856);
		when "1000000001011001" => data_out <= rom_array(32857);
		when "1000000001011010" => data_out <= rom_array(32858);
		when "1000000001011011" => data_out <= rom_array(32859);
		when "1000000001011100" => data_out <= rom_array(32860);
		when "1000000001011101" => data_out <= rom_array(32861);
		when "1000000001011110" => data_out <= rom_array(32862);
		when "1000000001011111" => data_out <= rom_array(32863);
		when "1000000001100000" => data_out <= rom_array(32864);
		when "1000000001100001" => data_out <= rom_array(32865);
		when "1000000001100010" => data_out <= rom_array(32866);
		when "1000000001100011" => data_out <= rom_array(32867);
		when "1000000001100100" => data_out <= rom_array(32868);
		when "1000000001100101" => data_out <= rom_array(32869);
		when "1000000001100110" => data_out <= rom_array(32870);
		when "1000000001100111" => data_out <= rom_array(32871);
		when "1000000001101000" => data_out <= rom_array(32872);
		when "1000000001101001" => data_out <= rom_array(32873);
		when "1000000001101010" => data_out <= rom_array(32874);
		when "1000000001101011" => data_out <= rom_array(32875);
		when "1000000001101100" => data_out <= rom_array(32876);
		when "1000000001101101" => data_out <= rom_array(32877);
		when "1000000001101110" => data_out <= rom_array(32878);
		when "1000000001101111" => data_out <= rom_array(32879);
		when "1000000001110000" => data_out <= rom_array(32880);
		when "1000000001110001" => data_out <= rom_array(32881);
		when "1000000001110010" => data_out <= rom_array(32882);
		when "1000000001110011" => data_out <= rom_array(32883);
		when "1000000001110100" => data_out <= rom_array(32884);
		when "1000000001110101" => data_out <= rom_array(32885);
		when "1000000001110110" => data_out <= rom_array(32886);
		when "1000000001110111" => data_out <= rom_array(32887);
		when "1000000001111000" => data_out <= rom_array(32888);
		when "1000000001111001" => data_out <= rom_array(32889);
		when "1000000001111010" => data_out <= rom_array(32890);
		when "1000000001111011" => data_out <= rom_array(32891);
		when "1000000001111100" => data_out <= rom_array(32892);
		when "1000000001111101" => data_out <= rom_array(32893);
		when "1000000001111110" => data_out <= rom_array(32894);
		when "1000000001111111" => data_out <= rom_array(32895);
		when "1000000010000000" => data_out <= rom_array(32896);
		when "1000000010000001" => data_out <= rom_array(32897);
		when "1000000010000010" => data_out <= rom_array(32898);
		when "1000000010000011" => data_out <= rom_array(32899);
		when "1000000010000100" => data_out <= rom_array(32900);
		when "1000000010000101" => data_out <= rom_array(32901);
		when "1000000010000110" => data_out <= rom_array(32902);
		when "1000000010000111" => data_out <= rom_array(32903);
		when "1000000010001000" => data_out <= rom_array(32904);
		when "1000000010001001" => data_out <= rom_array(32905);
		when "1000000010001010" => data_out <= rom_array(32906);
		when "1000000010001011" => data_out <= rom_array(32907);
		when "1000000010001100" => data_out <= rom_array(32908);
		when "1000000010001101" => data_out <= rom_array(32909);
		when "1000000010001110" => data_out <= rom_array(32910);
		when "1000000010001111" => data_out <= rom_array(32911);
		when "1000000010010000" => data_out <= rom_array(32912);
		when "1000000010010001" => data_out <= rom_array(32913);
		when "1000000010010010" => data_out <= rom_array(32914);
		when "1000000010010011" => data_out <= rom_array(32915);
		when "1000000010010100" => data_out <= rom_array(32916);
		when "1000000010010101" => data_out <= rom_array(32917);
		when "1000000010010110" => data_out <= rom_array(32918);
		when "1000000010010111" => data_out <= rom_array(32919);
		when "1000000010011000" => data_out <= rom_array(32920);
		when "1000000010011001" => data_out <= rom_array(32921);
		when "1000000010011010" => data_out <= rom_array(32922);
		when "1000000010011011" => data_out <= rom_array(32923);
		when "1000000010011100" => data_out <= rom_array(32924);
		when "1000000010011101" => data_out <= rom_array(32925);
		when "1000000010011110" => data_out <= rom_array(32926);
		when "1000000010011111" => data_out <= rom_array(32927);
		when "1000000010100000" => data_out <= rom_array(32928);
		when "1000000010100001" => data_out <= rom_array(32929);
		when "1000000010100010" => data_out <= rom_array(32930);
		when "1000000010100011" => data_out <= rom_array(32931);
		when "1000000010100100" => data_out <= rom_array(32932);
		when "1000000010100101" => data_out <= rom_array(32933);
		when "1000000010100110" => data_out <= rom_array(32934);
		when "1000000010100111" => data_out <= rom_array(32935);
		when "1000000010101000" => data_out <= rom_array(32936);
		when "1000000010101001" => data_out <= rom_array(32937);
		when "1000000010101010" => data_out <= rom_array(32938);
		when "1000000010101011" => data_out <= rom_array(32939);
		when "1000000010101100" => data_out <= rom_array(32940);
		when "1000000010101101" => data_out <= rom_array(32941);
		when "1000000010101110" => data_out <= rom_array(32942);
		when "1000000010101111" => data_out <= rom_array(32943);
		when "1000000010110000" => data_out <= rom_array(32944);
		when "1000000010110001" => data_out <= rom_array(32945);
		when "1000000010110010" => data_out <= rom_array(32946);
		when "1000000010110011" => data_out <= rom_array(32947);
		when "1000000010110100" => data_out <= rom_array(32948);
		when "1000000010110101" => data_out <= rom_array(32949);
		when "1000000010110110" => data_out <= rom_array(32950);
		when "1000000010110111" => data_out <= rom_array(32951);
		when "1000000010111000" => data_out <= rom_array(32952);
		when "1000000010111001" => data_out <= rom_array(32953);
		when "1000000010111010" => data_out <= rom_array(32954);
		when "1000000010111011" => data_out <= rom_array(32955);
		when "1000000010111100" => data_out <= rom_array(32956);
		when "1000000010111101" => data_out <= rom_array(32957);
		when "1000000010111110" => data_out <= rom_array(32958);
		when "1000000010111111" => data_out <= rom_array(32959);
		when "1000000011000000" => data_out <= rom_array(32960);
		when "1000000011000001" => data_out <= rom_array(32961);
		when "1000000011000010" => data_out <= rom_array(32962);
		when "1000000011000011" => data_out <= rom_array(32963);
		when "1000000011000100" => data_out <= rom_array(32964);
		when "1000000011000101" => data_out <= rom_array(32965);
		when "1000000011000110" => data_out <= rom_array(32966);
		when "1000000011000111" => data_out <= rom_array(32967);
		when "1000000011001000" => data_out <= rom_array(32968);
		when "1000000011001001" => data_out <= rom_array(32969);
		when "1000000011001010" => data_out <= rom_array(32970);
		when "1000000011001011" => data_out <= rom_array(32971);
		when "1000000011001100" => data_out <= rom_array(32972);
		when "1000000011001101" => data_out <= rom_array(32973);
		when "1000000011001110" => data_out <= rom_array(32974);
		when "1000000011001111" => data_out <= rom_array(32975);
		when "1000000011010000" => data_out <= rom_array(32976);
		when "1000000011010001" => data_out <= rom_array(32977);
		when "1000000011010010" => data_out <= rom_array(32978);
		when "1000000011010011" => data_out <= rom_array(32979);
		when "1000000011010100" => data_out <= rom_array(32980);
		when "1000000011010101" => data_out <= rom_array(32981);
		when "1000000011010110" => data_out <= rom_array(32982);
		when "1000000011010111" => data_out <= rom_array(32983);
		when "1000000011011000" => data_out <= rom_array(32984);
		when "1000000011011001" => data_out <= rom_array(32985);
		when "1000000011011010" => data_out <= rom_array(32986);
		when "1000000011011011" => data_out <= rom_array(32987);
		when "1000000011011100" => data_out <= rom_array(32988);
		when "1000000011011101" => data_out <= rom_array(32989);
		when "1000000011011110" => data_out <= rom_array(32990);
		when "1000000011011111" => data_out <= rom_array(32991);
		when "1000000011100000" => data_out <= rom_array(32992);
		when "1000000011100001" => data_out <= rom_array(32993);
		when "1000000011100010" => data_out <= rom_array(32994);
		when "1000000011100011" => data_out <= rom_array(32995);
		when "1000000011100100" => data_out <= rom_array(32996);
		when "1000000011100101" => data_out <= rom_array(32997);
		when "1000000011100110" => data_out <= rom_array(32998);
		when "1000000011100111" => data_out <= rom_array(32999);
		when "1000000011101000" => data_out <= rom_array(33000);
		when "1000000011101001" => data_out <= rom_array(33001);
		when "1000000011101010" => data_out <= rom_array(33002);
		when "1000000011101011" => data_out <= rom_array(33003);
		when "1000000011101100" => data_out <= rom_array(33004);
		when "1000000011101101" => data_out <= rom_array(33005);
		when "1000000011101110" => data_out <= rom_array(33006);
		when "1000000011101111" => data_out <= rom_array(33007);
		when "1000000011110000" => data_out <= rom_array(33008);
		when "1000000011110001" => data_out <= rom_array(33009);
		when "1000000011110010" => data_out <= rom_array(33010);
		when "1000000011110011" => data_out <= rom_array(33011);
		when "1000000011110100" => data_out <= rom_array(33012);
		when "1000000011110101" => data_out <= rom_array(33013);
		when "1000000011110110" => data_out <= rom_array(33014);
		when "1000000011110111" => data_out <= rom_array(33015);
		when "1000000011111000" => data_out <= rom_array(33016);
		when "1000000011111001" => data_out <= rom_array(33017);
		when "1000000011111010" => data_out <= rom_array(33018);
		when "1000000011111011" => data_out <= rom_array(33019);
		when "1000000011111100" => data_out <= rom_array(33020);
		when "1000000011111101" => data_out <= rom_array(33021);
		when "1000000011111110" => data_out <= rom_array(33022);
		when "1000000011111111" => data_out <= rom_array(33023);
		when "1000000100000000" => data_out <= rom_array(33024);
		when "1000000100000001" => data_out <= rom_array(33025);
		when "1000000100000010" => data_out <= rom_array(33026);
		when "1000000100000011" => data_out <= rom_array(33027);
		when "1000000100000100" => data_out <= rom_array(33028);
		when "1000000100000101" => data_out <= rom_array(33029);
		when "1000000100000110" => data_out <= rom_array(33030);
		when "1000000100000111" => data_out <= rom_array(33031);
		when "1000000100001000" => data_out <= rom_array(33032);
		when "1000000100001001" => data_out <= rom_array(33033);
		when "1000000100001010" => data_out <= rom_array(33034);
		when "1000000100001011" => data_out <= rom_array(33035);
		when "1000000100001100" => data_out <= rom_array(33036);
		when "1000000100001101" => data_out <= rom_array(33037);
		when "1000000100001110" => data_out <= rom_array(33038);
		when "1000000100001111" => data_out <= rom_array(33039);
		when "1000000100010000" => data_out <= rom_array(33040);
		when "1000000100010001" => data_out <= rom_array(33041);
		when "1000000100010010" => data_out <= rom_array(33042);
		when "1000000100010011" => data_out <= rom_array(33043);
		when "1000000100010100" => data_out <= rom_array(33044);
		when "1000000100010101" => data_out <= rom_array(33045);
		when "1000000100010110" => data_out <= rom_array(33046);
		when "1000000100010111" => data_out <= rom_array(33047);
		when "1000000100011000" => data_out <= rom_array(33048);
		when "1000000100011001" => data_out <= rom_array(33049);
		when "1000000100011010" => data_out <= rom_array(33050);
		when "1000000100011011" => data_out <= rom_array(33051);
		when "1000000100011100" => data_out <= rom_array(33052);
		when "1000000100011101" => data_out <= rom_array(33053);
		when "1000000100011110" => data_out <= rom_array(33054);
		when "1000000100011111" => data_out <= rom_array(33055);
		when "1000000100100000" => data_out <= rom_array(33056);
		when "1000000100100001" => data_out <= rom_array(33057);
		when "1000000100100010" => data_out <= rom_array(33058);
		when "1000000100100011" => data_out <= rom_array(33059);
		when "1000000100100100" => data_out <= rom_array(33060);
		when "1000000100100101" => data_out <= rom_array(33061);
		when "1000000100100110" => data_out <= rom_array(33062);
		when "1000000100100111" => data_out <= rom_array(33063);
		when "1000000100101000" => data_out <= rom_array(33064);
		when "1000000100101001" => data_out <= rom_array(33065);
		when "1000000100101010" => data_out <= rom_array(33066);
		when "1000000100101011" => data_out <= rom_array(33067);
		when "1000000100101100" => data_out <= rom_array(33068);
		when "1000000100101101" => data_out <= rom_array(33069);
		when "1000000100101110" => data_out <= rom_array(33070);
		when "1000000100101111" => data_out <= rom_array(33071);
		when "1000000100110000" => data_out <= rom_array(33072);
		when "1000000100110001" => data_out <= rom_array(33073);
		when "1000000100110010" => data_out <= rom_array(33074);
		when "1000000100110011" => data_out <= rom_array(33075);
		when "1000000100110100" => data_out <= rom_array(33076);
		when "1000000100110101" => data_out <= rom_array(33077);
		when "1000000100110110" => data_out <= rom_array(33078);
		when "1000000100110111" => data_out <= rom_array(33079);
		when "1000000100111000" => data_out <= rom_array(33080);
		when "1000000100111001" => data_out <= rom_array(33081);
		when "1000000100111010" => data_out <= rom_array(33082);
		when "1000000100111011" => data_out <= rom_array(33083);
		when "1000000100111100" => data_out <= rom_array(33084);
		when "1000000100111101" => data_out <= rom_array(33085);
		when "1000000100111110" => data_out <= rom_array(33086);
		when "1000000100111111" => data_out <= rom_array(33087);
		when "1000000101000000" => data_out <= rom_array(33088);
		when "1000000101000001" => data_out <= rom_array(33089);
		when "1000000101000010" => data_out <= rom_array(33090);
		when "1000000101000011" => data_out <= rom_array(33091);
		when "1000000101000100" => data_out <= rom_array(33092);
		when "1000000101000101" => data_out <= rom_array(33093);
		when "1000000101000110" => data_out <= rom_array(33094);
		when "1000000101000111" => data_out <= rom_array(33095);
		when "1000000101001000" => data_out <= rom_array(33096);
		when "1000000101001001" => data_out <= rom_array(33097);
		when "1000000101001010" => data_out <= rom_array(33098);
		when "1000000101001011" => data_out <= rom_array(33099);
		when "1000000101001100" => data_out <= rom_array(33100);
		when "1000000101001101" => data_out <= rom_array(33101);
		when "1000000101001110" => data_out <= rom_array(33102);
		when "1000000101001111" => data_out <= rom_array(33103);
		when "1000000101010000" => data_out <= rom_array(33104);
		when "1000000101010001" => data_out <= rom_array(33105);
		when "1000000101010010" => data_out <= rom_array(33106);
		when "1000000101010011" => data_out <= rom_array(33107);
		when "1000000101010100" => data_out <= rom_array(33108);
		when "1000000101010101" => data_out <= rom_array(33109);
		when "1000000101010110" => data_out <= rom_array(33110);
		when "1000000101010111" => data_out <= rom_array(33111);
		when "1000000101011000" => data_out <= rom_array(33112);
		when "1000000101011001" => data_out <= rom_array(33113);
		when "1000000101011010" => data_out <= rom_array(33114);
		when "1000000101011011" => data_out <= rom_array(33115);
		when "1000000101011100" => data_out <= rom_array(33116);
		when "1000000101011101" => data_out <= rom_array(33117);
		when "1000000101011110" => data_out <= rom_array(33118);
		when "1000000101011111" => data_out <= rom_array(33119);
		when "1000000101100000" => data_out <= rom_array(33120);
		when "1000000101100001" => data_out <= rom_array(33121);
		when "1000000101100010" => data_out <= rom_array(33122);
		when "1000000101100011" => data_out <= rom_array(33123);
		when "1000000101100100" => data_out <= rom_array(33124);
		when "1000000101100101" => data_out <= rom_array(33125);
		when "1000000101100110" => data_out <= rom_array(33126);
		when "1000000101100111" => data_out <= rom_array(33127);
		when "1000000101101000" => data_out <= rom_array(33128);
		when "1000000101101001" => data_out <= rom_array(33129);
		when "1000000101101010" => data_out <= rom_array(33130);
		when "1000000101101011" => data_out <= rom_array(33131);
		when "1000000101101100" => data_out <= rom_array(33132);
		when "1000000101101101" => data_out <= rom_array(33133);
		when "1000000101101110" => data_out <= rom_array(33134);
		when "1000000101101111" => data_out <= rom_array(33135);
		when "1000000101110000" => data_out <= rom_array(33136);
		when "1000000101110001" => data_out <= rom_array(33137);
		when "1000000101110010" => data_out <= rom_array(33138);
		when "1000000101110011" => data_out <= rom_array(33139);
		when "1000000101110100" => data_out <= rom_array(33140);
		when "1000000101110101" => data_out <= rom_array(33141);
		when "1000000101110110" => data_out <= rom_array(33142);
		when "1000000101110111" => data_out <= rom_array(33143);
		when "1000000101111000" => data_out <= rom_array(33144);
		when "1000000101111001" => data_out <= rom_array(33145);
		when "1000000101111010" => data_out <= rom_array(33146);
		when "1000000101111011" => data_out <= rom_array(33147);
		when "1000000101111100" => data_out <= rom_array(33148);
		when "1000000101111101" => data_out <= rom_array(33149);
		when "1000000101111110" => data_out <= rom_array(33150);
		when "1000000101111111" => data_out <= rom_array(33151);
		when "1000000110000000" => data_out <= rom_array(33152);
		when "1000000110000001" => data_out <= rom_array(33153);
		when "1000000110000010" => data_out <= rom_array(33154);
		when "1000000110000011" => data_out <= rom_array(33155);
		when "1000000110000100" => data_out <= rom_array(33156);
		when "1000000110000101" => data_out <= rom_array(33157);
		when "1000000110000110" => data_out <= rom_array(33158);
		when "1000000110000111" => data_out <= rom_array(33159);
		when "1000000110001000" => data_out <= rom_array(33160);
		when "1000000110001001" => data_out <= rom_array(33161);
		when "1000000110001010" => data_out <= rom_array(33162);
		when "1000000110001011" => data_out <= rom_array(33163);
		when "1000000110001100" => data_out <= rom_array(33164);
		when "1000000110001101" => data_out <= rom_array(33165);
		when "1000000110001110" => data_out <= rom_array(33166);
		when "1000000110001111" => data_out <= rom_array(33167);
		when "1000000110010000" => data_out <= rom_array(33168);
		when "1000000110010001" => data_out <= rom_array(33169);
		when "1000000110010010" => data_out <= rom_array(33170);
		when "1000000110010011" => data_out <= rom_array(33171);
		when "1000000110010100" => data_out <= rom_array(33172);
		when "1000000110010101" => data_out <= rom_array(33173);
		when "1000000110010110" => data_out <= rom_array(33174);
		when "1000000110010111" => data_out <= rom_array(33175);
		when "1000000110011000" => data_out <= rom_array(33176);
		when "1000000110011001" => data_out <= rom_array(33177);
		when "1000000110011010" => data_out <= rom_array(33178);
		when "1000000110011011" => data_out <= rom_array(33179);
		when "1000000110011100" => data_out <= rom_array(33180);
		when "1000000110011101" => data_out <= rom_array(33181);
		when "1000000110011110" => data_out <= rom_array(33182);
		when "1000000110011111" => data_out <= rom_array(33183);
		when "1000000110100000" => data_out <= rom_array(33184);
		when "1000000110100001" => data_out <= rom_array(33185);
		when "1000000110100010" => data_out <= rom_array(33186);
		when "1000000110100011" => data_out <= rom_array(33187);
		when "1000000110100100" => data_out <= rom_array(33188);
		when "1000000110100101" => data_out <= rom_array(33189);
		when "1000000110100110" => data_out <= rom_array(33190);
		when "1000000110100111" => data_out <= rom_array(33191);
		when "1000000110101000" => data_out <= rom_array(33192);
		when "1000000110101001" => data_out <= rom_array(33193);
		when "1000000110101010" => data_out <= rom_array(33194);
		when "1000000110101011" => data_out <= rom_array(33195);
		when "1000000110101100" => data_out <= rom_array(33196);
		when "1000000110101101" => data_out <= rom_array(33197);
		when "1000000110101110" => data_out <= rom_array(33198);
		when "1000000110101111" => data_out <= rom_array(33199);
		when "1000000110110000" => data_out <= rom_array(33200);
		when "1000000110110001" => data_out <= rom_array(33201);
		when "1000000110110010" => data_out <= rom_array(33202);
		when "1000000110110011" => data_out <= rom_array(33203);
		when "1000000110110100" => data_out <= rom_array(33204);
		when "1000000110110101" => data_out <= rom_array(33205);
		when "1000000110110110" => data_out <= rom_array(33206);
		when "1000000110110111" => data_out <= rom_array(33207);
		when "1000000110111000" => data_out <= rom_array(33208);
		when "1000000110111001" => data_out <= rom_array(33209);
		when "1000000110111010" => data_out <= rom_array(33210);
		when "1000000110111011" => data_out <= rom_array(33211);
		when "1000000110111100" => data_out <= rom_array(33212);
		when "1000000110111101" => data_out <= rom_array(33213);
		when "1000000110111110" => data_out <= rom_array(33214);
		when "1000000110111111" => data_out <= rom_array(33215);
		when "1000000111000000" => data_out <= rom_array(33216);
		when "1000000111000001" => data_out <= rom_array(33217);
		when "1000000111000010" => data_out <= rom_array(33218);
		when "1000000111000011" => data_out <= rom_array(33219);
		when "1000000111000100" => data_out <= rom_array(33220);
		when "1000000111000101" => data_out <= rom_array(33221);
		when "1000000111000110" => data_out <= rom_array(33222);
		when "1000000111000111" => data_out <= rom_array(33223);
		when "1000000111001000" => data_out <= rom_array(33224);
		when "1000000111001001" => data_out <= rom_array(33225);
		when "1000000111001010" => data_out <= rom_array(33226);
		when "1000000111001011" => data_out <= rom_array(33227);
		when "1000000111001100" => data_out <= rom_array(33228);
		when "1000000111001101" => data_out <= rom_array(33229);
		when "1000000111001110" => data_out <= rom_array(33230);
		when "1000000111001111" => data_out <= rom_array(33231);
		when "1000000111010000" => data_out <= rom_array(33232);
		when "1000000111010001" => data_out <= rom_array(33233);
		when "1000000111010010" => data_out <= rom_array(33234);
		when "1000000111010011" => data_out <= rom_array(33235);
		when "1000000111010100" => data_out <= rom_array(33236);
		when "1000000111010101" => data_out <= rom_array(33237);
		when "1000000111010110" => data_out <= rom_array(33238);
		when "1000000111010111" => data_out <= rom_array(33239);
		when "1000000111011000" => data_out <= rom_array(33240);
		when "1000000111011001" => data_out <= rom_array(33241);
		when "1000000111011010" => data_out <= rom_array(33242);
		when "1000000111011011" => data_out <= rom_array(33243);
		when "1000000111011100" => data_out <= rom_array(33244);
		when "1000000111011101" => data_out <= rom_array(33245);
		when "1000000111011110" => data_out <= rom_array(33246);
		when "1000000111011111" => data_out <= rom_array(33247);
		when "1000000111100000" => data_out <= rom_array(33248);
		when "1000000111100001" => data_out <= rom_array(33249);
		when "1000000111100010" => data_out <= rom_array(33250);
		when "1000000111100011" => data_out <= rom_array(33251);
		when "1000000111100100" => data_out <= rom_array(33252);
		when "1000000111100101" => data_out <= rom_array(33253);
		when "1000000111100110" => data_out <= rom_array(33254);
		when "1000000111100111" => data_out <= rom_array(33255);
		when "1000000111101000" => data_out <= rom_array(33256);
		when "1000000111101001" => data_out <= rom_array(33257);
		when "1000000111101010" => data_out <= rom_array(33258);
		when "1000000111101011" => data_out <= rom_array(33259);
		when "1000000111101100" => data_out <= rom_array(33260);
		when "1000000111101101" => data_out <= rom_array(33261);
		when "1000000111101110" => data_out <= rom_array(33262);
		when "1000000111101111" => data_out <= rom_array(33263);
		when "1000000111110000" => data_out <= rom_array(33264);
		when "1000000111110001" => data_out <= rom_array(33265);
		when "1000000111110010" => data_out <= rom_array(33266);
		when "1000000111110011" => data_out <= rom_array(33267);
		when "1000000111110100" => data_out <= rom_array(33268);
		when "1000000111110101" => data_out <= rom_array(33269);
		when "1000000111110110" => data_out <= rom_array(33270);
		when "1000000111110111" => data_out <= rom_array(33271);
		when "1000000111111000" => data_out <= rom_array(33272);
		when "1000000111111001" => data_out <= rom_array(33273);
		when "1000000111111010" => data_out <= rom_array(33274);
		when "1000000111111011" => data_out <= rom_array(33275);
		when "1000000111111100" => data_out <= rom_array(33276);
		when "1000000111111101" => data_out <= rom_array(33277);
		when "1000000111111110" => data_out <= rom_array(33278);
		when "1000000111111111" => data_out <= rom_array(33279);
		when "1000001000000000" => data_out <= rom_array(33280);
		when "1000001000000001" => data_out <= rom_array(33281);
		when "1000001000000010" => data_out <= rom_array(33282);
		when "1000001000000011" => data_out <= rom_array(33283);
		when "1000001000000100" => data_out <= rom_array(33284);
		when "1000001000000101" => data_out <= rom_array(33285);
		when "1000001000000110" => data_out <= rom_array(33286);
		when "1000001000000111" => data_out <= rom_array(33287);
		when "1000001000001000" => data_out <= rom_array(33288);
		when "1000001000001001" => data_out <= rom_array(33289);
		when "1000001000001010" => data_out <= rom_array(33290);
		when "1000001000001011" => data_out <= rom_array(33291);
		when "1000001000001100" => data_out <= rom_array(33292);
		when "1000001000001101" => data_out <= rom_array(33293);
		when "1000001000001110" => data_out <= rom_array(33294);
		when "1000001000001111" => data_out <= rom_array(33295);
		when "1000001000010000" => data_out <= rom_array(33296);
		when "1000001000010001" => data_out <= rom_array(33297);
		when "1000001000010010" => data_out <= rom_array(33298);
		when "1000001000010011" => data_out <= rom_array(33299);
		when "1000001000010100" => data_out <= rom_array(33300);
		when "1000001000010101" => data_out <= rom_array(33301);
		when "1000001000010110" => data_out <= rom_array(33302);
		when "1000001000010111" => data_out <= rom_array(33303);
		when "1000001000011000" => data_out <= rom_array(33304);
		when "1000001000011001" => data_out <= rom_array(33305);
		when "1000001000011010" => data_out <= rom_array(33306);
		when "1000001000011011" => data_out <= rom_array(33307);
		when "1000001000011100" => data_out <= rom_array(33308);
		when "1000001000011101" => data_out <= rom_array(33309);
		when "1000001000011110" => data_out <= rom_array(33310);
		when "1000001000011111" => data_out <= rom_array(33311);
		when "1000001000100000" => data_out <= rom_array(33312);
		when "1000001000100001" => data_out <= rom_array(33313);
		when "1000001000100010" => data_out <= rom_array(33314);
		when "1000001000100011" => data_out <= rom_array(33315);
		when "1000001000100100" => data_out <= rom_array(33316);
		when "1000001000100101" => data_out <= rom_array(33317);
		when "1000001000100110" => data_out <= rom_array(33318);
		when "1000001000100111" => data_out <= rom_array(33319);
		when "1000001000101000" => data_out <= rom_array(33320);
		when "1000001000101001" => data_out <= rom_array(33321);
		when "1000001000101010" => data_out <= rom_array(33322);
		when "1000001000101011" => data_out <= rom_array(33323);
		when "1000001000101100" => data_out <= rom_array(33324);
		when "1000001000101101" => data_out <= rom_array(33325);
		when "1000001000101110" => data_out <= rom_array(33326);
		when "1000001000101111" => data_out <= rom_array(33327);
		when "1000001000110000" => data_out <= rom_array(33328);
		when "1000001000110001" => data_out <= rom_array(33329);
		when "1000001000110010" => data_out <= rom_array(33330);
		when "1000001000110011" => data_out <= rom_array(33331);
		when "1000001000110100" => data_out <= rom_array(33332);
		when "1000001000110101" => data_out <= rom_array(33333);
		when "1000001000110110" => data_out <= rom_array(33334);
		when "1000001000110111" => data_out <= rom_array(33335);
		when "1000001000111000" => data_out <= rom_array(33336);
		when "1000001000111001" => data_out <= rom_array(33337);
		when "1000001000111010" => data_out <= rom_array(33338);
		when "1000001000111011" => data_out <= rom_array(33339);
		when "1000001000111100" => data_out <= rom_array(33340);
		when "1000001000111101" => data_out <= rom_array(33341);
		when "1000001000111110" => data_out <= rom_array(33342);
		when "1000001000111111" => data_out <= rom_array(33343);
		when "1000001001000000" => data_out <= rom_array(33344);
		when "1000001001000001" => data_out <= rom_array(33345);
		when "1000001001000010" => data_out <= rom_array(33346);
		when "1000001001000011" => data_out <= rom_array(33347);
		when "1000001001000100" => data_out <= rom_array(33348);
		when "1000001001000101" => data_out <= rom_array(33349);
		when "1000001001000110" => data_out <= rom_array(33350);
		when "1000001001000111" => data_out <= rom_array(33351);
		when "1000001001001000" => data_out <= rom_array(33352);
		when "1000001001001001" => data_out <= rom_array(33353);
		when "1000001001001010" => data_out <= rom_array(33354);
		when "1000001001001011" => data_out <= rom_array(33355);
		when "1000001001001100" => data_out <= rom_array(33356);
		when "1000001001001101" => data_out <= rom_array(33357);
		when "1000001001001110" => data_out <= rom_array(33358);
		when "1000001001001111" => data_out <= rom_array(33359);
		when "1000001001010000" => data_out <= rom_array(33360);
		when "1000001001010001" => data_out <= rom_array(33361);
		when "1000001001010010" => data_out <= rom_array(33362);
		when "1000001001010011" => data_out <= rom_array(33363);
		when "1000001001010100" => data_out <= rom_array(33364);
		when "1000001001010101" => data_out <= rom_array(33365);
		when "1000001001010110" => data_out <= rom_array(33366);
		when "1000001001010111" => data_out <= rom_array(33367);
		when "1000001001011000" => data_out <= rom_array(33368);
		when "1000001001011001" => data_out <= rom_array(33369);
		when "1000001001011010" => data_out <= rom_array(33370);
		when "1000001001011011" => data_out <= rom_array(33371);
		when "1000001001011100" => data_out <= rom_array(33372);
		when "1000001001011101" => data_out <= rom_array(33373);
		when "1000001001011110" => data_out <= rom_array(33374);
		when "1000001001011111" => data_out <= rom_array(33375);
		when "1000001001100000" => data_out <= rom_array(33376);
		when "1000001001100001" => data_out <= rom_array(33377);
		when "1000001001100010" => data_out <= rom_array(33378);
		when "1000001001100011" => data_out <= rom_array(33379);
		when "1000001001100100" => data_out <= rom_array(33380);
		when "1000001001100101" => data_out <= rom_array(33381);
		when "1000001001100110" => data_out <= rom_array(33382);
		when "1000001001100111" => data_out <= rom_array(33383);
		when "1000001001101000" => data_out <= rom_array(33384);
		when "1000001001101001" => data_out <= rom_array(33385);
		when "1000001001101010" => data_out <= rom_array(33386);
		when "1000001001101011" => data_out <= rom_array(33387);
		when "1000001001101100" => data_out <= rom_array(33388);
		when "1000001001101101" => data_out <= rom_array(33389);
		when "1000001001101110" => data_out <= rom_array(33390);
		when "1000001001101111" => data_out <= rom_array(33391);
		when "1000001001110000" => data_out <= rom_array(33392);
		when "1000001001110001" => data_out <= rom_array(33393);
		when "1000001001110010" => data_out <= rom_array(33394);
		when "1000001001110011" => data_out <= rom_array(33395);
		when "1000001001110100" => data_out <= rom_array(33396);
		when "1000001001110101" => data_out <= rom_array(33397);
		when "1000001001110110" => data_out <= rom_array(33398);
		when "1000001001110111" => data_out <= rom_array(33399);
		when "1000001001111000" => data_out <= rom_array(33400);
		when "1000001001111001" => data_out <= rom_array(33401);
		when "1000001001111010" => data_out <= rom_array(33402);
		when "1000001001111011" => data_out <= rom_array(33403);
		when "1000001001111100" => data_out <= rom_array(33404);
		when "1000001001111101" => data_out <= rom_array(33405);
		when "1000001001111110" => data_out <= rom_array(33406);
		when "1000001001111111" => data_out <= rom_array(33407);
		when "1000001010000000" => data_out <= rom_array(33408);
		when "1000001010000001" => data_out <= rom_array(33409);
		when "1000001010000010" => data_out <= rom_array(33410);
		when "1000001010000011" => data_out <= rom_array(33411);
		when "1000001010000100" => data_out <= rom_array(33412);
		when "1000001010000101" => data_out <= rom_array(33413);
		when "1000001010000110" => data_out <= rom_array(33414);
		when "1000001010000111" => data_out <= rom_array(33415);
		when "1000001010001000" => data_out <= rom_array(33416);
		when "1000001010001001" => data_out <= rom_array(33417);
		when "1000001010001010" => data_out <= rom_array(33418);
		when "1000001010001011" => data_out <= rom_array(33419);
		when "1000001010001100" => data_out <= rom_array(33420);
		when "1000001010001101" => data_out <= rom_array(33421);
		when "1000001010001110" => data_out <= rom_array(33422);
		when "1000001010001111" => data_out <= rom_array(33423);
		when "1000001010010000" => data_out <= rom_array(33424);
		when "1000001010010001" => data_out <= rom_array(33425);
		when "1000001010010010" => data_out <= rom_array(33426);
		when "1000001010010011" => data_out <= rom_array(33427);
		when "1000001010010100" => data_out <= rom_array(33428);
		when "1000001010010101" => data_out <= rom_array(33429);
		when "1000001010010110" => data_out <= rom_array(33430);
		when "1000001010010111" => data_out <= rom_array(33431);
		when "1000001010011000" => data_out <= rom_array(33432);
		when "1000001010011001" => data_out <= rom_array(33433);
		when "1000001010011010" => data_out <= rom_array(33434);
		when "1000001010011011" => data_out <= rom_array(33435);
		when "1000001010011100" => data_out <= rom_array(33436);
		when "1000001010011101" => data_out <= rom_array(33437);
		when "1000001010011110" => data_out <= rom_array(33438);
		when "1000001010011111" => data_out <= rom_array(33439);
		when "1000001010100000" => data_out <= rom_array(33440);
		when "1000001010100001" => data_out <= rom_array(33441);
		when "1000001010100010" => data_out <= rom_array(33442);
		when "1000001010100011" => data_out <= rom_array(33443);
		when "1000001010100100" => data_out <= rom_array(33444);
		when "1000001010100101" => data_out <= rom_array(33445);
		when "1000001010100110" => data_out <= rom_array(33446);
		when "1000001010100111" => data_out <= rom_array(33447);
		when "1000001010101000" => data_out <= rom_array(33448);
		when "1000001010101001" => data_out <= rom_array(33449);
		when "1000001010101010" => data_out <= rom_array(33450);
		when "1000001010101011" => data_out <= rom_array(33451);
		when "1000001010101100" => data_out <= rom_array(33452);
		when "1000001010101101" => data_out <= rom_array(33453);
		when "1000001010101110" => data_out <= rom_array(33454);
		when "1000001010101111" => data_out <= rom_array(33455);
		when "1000001010110000" => data_out <= rom_array(33456);
		when "1000001010110001" => data_out <= rom_array(33457);
		when "1000001010110010" => data_out <= rom_array(33458);
		when "1000001010110011" => data_out <= rom_array(33459);
		when "1000001010110100" => data_out <= rom_array(33460);
		when "1000001010110101" => data_out <= rom_array(33461);
		when "1000001010110110" => data_out <= rom_array(33462);
		when "1000001010110111" => data_out <= rom_array(33463);
		when "1000001010111000" => data_out <= rom_array(33464);
		when "1000001010111001" => data_out <= rom_array(33465);
		when "1000001010111010" => data_out <= rom_array(33466);
		when "1000001010111011" => data_out <= rom_array(33467);
		when "1000001010111100" => data_out <= rom_array(33468);
		when "1000001010111101" => data_out <= rom_array(33469);
		when "1000001010111110" => data_out <= rom_array(33470);
		when "1000001010111111" => data_out <= rom_array(33471);
		when "1000001011000000" => data_out <= rom_array(33472);
		when "1000001011000001" => data_out <= rom_array(33473);
		when "1000001011000010" => data_out <= rom_array(33474);
		when "1000001011000011" => data_out <= rom_array(33475);
		when "1000001011000100" => data_out <= rom_array(33476);
		when "1000001011000101" => data_out <= rom_array(33477);
		when "1000001011000110" => data_out <= rom_array(33478);
		when "1000001011000111" => data_out <= rom_array(33479);
		when "1000001011001000" => data_out <= rom_array(33480);
		when "1000001011001001" => data_out <= rom_array(33481);
		when "1000001011001010" => data_out <= rom_array(33482);
		when "1000001011001011" => data_out <= rom_array(33483);
		when "1000001011001100" => data_out <= rom_array(33484);
		when "1000001011001101" => data_out <= rom_array(33485);
		when "1000001011001110" => data_out <= rom_array(33486);
		when "1000001011001111" => data_out <= rom_array(33487);
		when "1000001011010000" => data_out <= rom_array(33488);
		when "1000001011010001" => data_out <= rom_array(33489);
		when "1000001011010010" => data_out <= rom_array(33490);
		when "1000001011010011" => data_out <= rom_array(33491);
		when "1000001011010100" => data_out <= rom_array(33492);
		when "1000001011010101" => data_out <= rom_array(33493);
		when "1000001011010110" => data_out <= rom_array(33494);
		when "1000001011010111" => data_out <= rom_array(33495);
		when "1000001011011000" => data_out <= rom_array(33496);
		when "1000001011011001" => data_out <= rom_array(33497);
		when "1000001011011010" => data_out <= rom_array(33498);
		when "1000001011011011" => data_out <= rom_array(33499);
		when "1000001011011100" => data_out <= rom_array(33500);
		when "1000001011011101" => data_out <= rom_array(33501);
		when "1000001011011110" => data_out <= rom_array(33502);
		when "1000001011011111" => data_out <= rom_array(33503);
		when "1000001011100000" => data_out <= rom_array(33504);
		when "1000001011100001" => data_out <= rom_array(33505);
		when "1000001011100010" => data_out <= rom_array(33506);
		when "1000001011100011" => data_out <= rom_array(33507);
		when "1000001011100100" => data_out <= rom_array(33508);
		when "1000001011100101" => data_out <= rom_array(33509);
		when "1000001011100110" => data_out <= rom_array(33510);
		when "1000001011100111" => data_out <= rom_array(33511);
		when "1000001011101000" => data_out <= rom_array(33512);
		when "1000001011101001" => data_out <= rom_array(33513);
		when "1000001011101010" => data_out <= rom_array(33514);
		when "1000001011101011" => data_out <= rom_array(33515);
		when "1000001011101100" => data_out <= rom_array(33516);
		when "1000001011101101" => data_out <= rom_array(33517);
		when "1000001011101110" => data_out <= rom_array(33518);
		when "1000001011101111" => data_out <= rom_array(33519);
		when "1000001011110000" => data_out <= rom_array(33520);
		when "1000001011110001" => data_out <= rom_array(33521);
		when "1000001011110010" => data_out <= rom_array(33522);
		when "1000001011110011" => data_out <= rom_array(33523);
		when "1000001011110100" => data_out <= rom_array(33524);
		when "1000001011110101" => data_out <= rom_array(33525);
		when "1000001011110110" => data_out <= rom_array(33526);
		when "1000001011110111" => data_out <= rom_array(33527);
		when "1000001011111000" => data_out <= rom_array(33528);
		when "1000001011111001" => data_out <= rom_array(33529);
		when "1000001011111010" => data_out <= rom_array(33530);
		when "1000001011111011" => data_out <= rom_array(33531);
		when "1000001011111100" => data_out <= rom_array(33532);
		when "1000001011111101" => data_out <= rom_array(33533);
		when "1000001011111110" => data_out <= rom_array(33534);
		when "1000001011111111" => data_out <= rom_array(33535);
		when "1000001100000000" => data_out <= rom_array(33536);
		when "1000001100000001" => data_out <= rom_array(33537);
		when "1000001100000010" => data_out <= rom_array(33538);
		when "1000001100000011" => data_out <= rom_array(33539);
		when "1000001100000100" => data_out <= rom_array(33540);
		when "1000001100000101" => data_out <= rom_array(33541);
		when "1000001100000110" => data_out <= rom_array(33542);
		when "1000001100000111" => data_out <= rom_array(33543);
		when "1000001100001000" => data_out <= rom_array(33544);
		when "1000001100001001" => data_out <= rom_array(33545);
		when "1000001100001010" => data_out <= rom_array(33546);
		when "1000001100001011" => data_out <= rom_array(33547);
		when "1000001100001100" => data_out <= rom_array(33548);
		when "1000001100001101" => data_out <= rom_array(33549);
		when "1000001100001110" => data_out <= rom_array(33550);
		when "1000001100001111" => data_out <= rom_array(33551);
		when "1000001100010000" => data_out <= rom_array(33552);
		when "1000001100010001" => data_out <= rom_array(33553);
		when "1000001100010010" => data_out <= rom_array(33554);
		when "1000001100010011" => data_out <= rom_array(33555);
		when "1000001100010100" => data_out <= rom_array(33556);
		when "1000001100010101" => data_out <= rom_array(33557);
		when "1000001100010110" => data_out <= rom_array(33558);
		when "1000001100010111" => data_out <= rom_array(33559);
		when "1000001100011000" => data_out <= rom_array(33560);
		when "1000001100011001" => data_out <= rom_array(33561);
		when "1000001100011010" => data_out <= rom_array(33562);
		when "1000001100011011" => data_out <= rom_array(33563);
		when "1000001100011100" => data_out <= rom_array(33564);
		when "1000001100011101" => data_out <= rom_array(33565);
		when "1000001100011110" => data_out <= rom_array(33566);
		when "1000001100011111" => data_out <= rom_array(33567);
		when "1000001100100000" => data_out <= rom_array(33568);
		when "1000001100100001" => data_out <= rom_array(33569);
		when "1000001100100010" => data_out <= rom_array(33570);
		when "1000001100100011" => data_out <= rom_array(33571);
		when "1000001100100100" => data_out <= rom_array(33572);
		when "1000001100100101" => data_out <= rom_array(33573);
		when "1000001100100110" => data_out <= rom_array(33574);
		when "1000001100100111" => data_out <= rom_array(33575);
		when "1000001100101000" => data_out <= rom_array(33576);
		when "1000001100101001" => data_out <= rom_array(33577);
		when "1000001100101010" => data_out <= rom_array(33578);
		when "1000001100101011" => data_out <= rom_array(33579);
		when "1000001100101100" => data_out <= rom_array(33580);
		when "1000001100101101" => data_out <= rom_array(33581);
		when "1000001100101110" => data_out <= rom_array(33582);
		when "1000001100101111" => data_out <= rom_array(33583);
		when "1000001100110000" => data_out <= rom_array(33584);
		when "1000001100110001" => data_out <= rom_array(33585);
		when "1000001100110010" => data_out <= rom_array(33586);
		when "1000001100110011" => data_out <= rom_array(33587);
		when "1000001100110100" => data_out <= rom_array(33588);
		when "1000001100110101" => data_out <= rom_array(33589);
		when "1000001100110110" => data_out <= rom_array(33590);
		when "1000001100110111" => data_out <= rom_array(33591);
		when "1000001100111000" => data_out <= rom_array(33592);
		when "1000001100111001" => data_out <= rom_array(33593);
		when "1000001100111010" => data_out <= rom_array(33594);
		when "1000001100111011" => data_out <= rom_array(33595);
		when "1000001100111100" => data_out <= rom_array(33596);
		when "1000001100111101" => data_out <= rom_array(33597);
		when "1000001100111110" => data_out <= rom_array(33598);
		when "1000001100111111" => data_out <= rom_array(33599);
		when "1000001101000000" => data_out <= rom_array(33600);
		when "1000001101000001" => data_out <= rom_array(33601);
		when "1000001101000010" => data_out <= rom_array(33602);
		when "1000001101000011" => data_out <= rom_array(33603);
		when "1000001101000100" => data_out <= rom_array(33604);
		when "1000001101000101" => data_out <= rom_array(33605);
		when "1000001101000110" => data_out <= rom_array(33606);
		when "1000001101000111" => data_out <= rom_array(33607);
		when "1000001101001000" => data_out <= rom_array(33608);
		when "1000001101001001" => data_out <= rom_array(33609);
		when "1000001101001010" => data_out <= rom_array(33610);
		when "1000001101001011" => data_out <= rom_array(33611);
		when "1000001101001100" => data_out <= rom_array(33612);
		when "1000001101001101" => data_out <= rom_array(33613);
		when "1000001101001110" => data_out <= rom_array(33614);
		when "1000001101001111" => data_out <= rom_array(33615);
		when "1000001101010000" => data_out <= rom_array(33616);
		when "1000001101010001" => data_out <= rom_array(33617);
		when "1000001101010010" => data_out <= rom_array(33618);
		when "1000001101010011" => data_out <= rom_array(33619);
		when "1000001101010100" => data_out <= rom_array(33620);
		when "1000001101010101" => data_out <= rom_array(33621);
		when "1000001101010110" => data_out <= rom_array(33622);
		when "1000001101010111" => data_out <= rom_array(33623);
		when "1000001101011000" => data_out <= rom_array(33624);
		when "1000001101011001" => data_out <= rom_array(33625);
		when "1000001101011010" => data_out <= rom_array(33626);
		when "1000001101011011" => data_out <= rom_array(33627);
		when "1000001101011100" => data_out <= rom_array(33628);
		when "1000001101011101" => data_out <= rom_array(33629);
		when "1000001101011110" => data_out <= rom_array(33630);
		when "1000001101011111" => data_out <= rom_array(33631);
		when "1000001101100000" => data_out <= rom_array(33632);
		when "1000001101100001" => data_out <= rom_array(33633);
		when "1000001101100010" => data_out <= rom_array(33634);
		when "1000001101100011" => data_out <= rom_array(33635);
		when "1000001101100100" => data_out <= rom_array(33636);
		when "1000001101100101" => data_out <= rom_array(33637);
		when "1000001101100110" => data_out <= rom_array(33638);
		when "1000001101100111" => data_out <= rom_array(33639);
		when "1000001101101000" => data_out <= rom_array(33640);
		when "1000001101101001" => data_out <= rom_array(33641);
		when "1000001101101010" => data_out <= rom_array(33642);
		when "1000001101101011" => data_out <= rom_array(33643);
		when "1000001101101100" => data_out <= rom_array(33644);
		when "1000001101101101" => data_out <= rom_array(33645);
		when "1000001101101110" => data_out <= rom_array(33646);
		when "1000001101101111" => data_out <= rom_array(33647);
		when "1000001101110000" => data_out <= rom_array(33648);
		when "1000001101110001" => data_out <= rom_array(33649);
		when "1000001101110010" => data_out <= rom_array(33650);
		when "1000001101110011" => data_out <= rom_array(33651);
		when "1000001101110100" => data_out <= rom_array(33652);
		when "1000001101110101" => data_out <= rom_array(33653);
		when "1000001101110110" => data_out <= rom_array(33654);
		when "1000001101110111" => data_out <= rom_array(33655);
		when "1000001101111000" => data_out <= rom_array(33656);
		when "1000001101111001" => data_out <= rom_array(33657);
		when "1000001101111010" => data_out <= rom_array(33658);
		when "1000001101111011" => data_out <= rom_array(33659);
		when "1000001101111100" => data_out <= rom_array(33660);
		when "1000001101111101" => data_out <= rom_array(33661);
		when "1000001101111110" => data_out <= rom_array(33662);
		when "1000001101111111" => data_out <= rom_array(33663);
		when "1000001110000000" => data_out <= rom_array(33664);
		when "1000001110000001" => data_out <= rom_array(33665);
		when "1000001110000010" => data_out <= rom_array(33666);
		when "1000001110000011" => data_out <= rom_array(33667);
		when "1000001110000100" => data_out <= rom_array(33668);
		when "1000001110000101" => data_out <= rom_array(33669);
		when "1000001110000110" => data_out <= rom_array(33670);
		when "1000001110000111" => data_out <= rom_array(33671);
		when "1000001110001000" => data_out <= rom_array(33672);
		when "1000001110001001" => data_out <= rom_array(33673);
		when "1000001110001010" => data_out <= rom_array(33674);
		when "1000001110001011" => data_out <= rom_array(33675);
		when "1000001110001100" => data_out <= rom_array(33676);
		when "1000001110001101" => data_out <= rom_array(33677);
		when "1000001110001110" => data_out <= rom_array(33678);
		when "1000001110001111" => data_out <= rom_array(33679);
		when "1000001110010000" => data_out <= rom_array(33680);
		when "1000001110010001" => data_out <= rom_array(33681);
		when "1000001110010010" => data_out <= rom_array(33682);
		when "1000001110010011" => data_out <= rom_array(33683);
		when "1000001110010100" => data_out <= rom_array(33684);
		when "1000001110010101" => data_out <= rom_array(33685);
		when "1000001110010110" => data_out <= rom_array(33686);
		when "1000001110010111" => data_out <= rom_array(33687);
		when "1000001110011000" => data_out <= rom_array(33688);
		when "1000001110011001" => data_out <= rom_array(33689);
		when "1000001110011010" => data_out <= rom_array(33690);
		when "1000001110011011" => data_out <= rom_array(33691);
		when "1000001110011100" => data_out <= rom_array(33692);
		when "1000001110011101" => data_out <= rom_array(33693);
		when "1000001110011110" => data_out <= rom_array(33694);
		when "1000001110011111" => data_out <= rom_array(33695);
		when "1000001110100000" => data_out <= rom_array(33696);
		when "1000001110100001" => data_out <= rom_array(33697);
		when "1000001110100010" => data_out <= rom_array(33698);
		when "1000001110100011" => data_out <= rom_array(33699);
		when "1000001110100100" => data_out <= rom_array(33700);
		when "1000001110100101" => data_out <= rom_array(33701);
		when "1000001110100110" => data_out <= rom_array(33702);
		when "1000001110100111" => data_out <= rom_array(33703);
		when "1000001110101000" => data_out <= rom_array(33704);
		when "1000001110101001" => data_out <= rom_array(33705);
		when "1000001110101010" => data_out <= rom_array(33706);
		when "1000001110101011" => data_out <= rom_array(33707);
		when "1000001110101100" => data_out <= rom_array(33708);
		when "1000001110101101" => data_out <= rom_array(33709);
		when "1000001110101110" => data_out <= rom_array(33710);
		when "1000001110101111" => data_out <= rom_array(33711);
		when "1000001110110000" => data_out <= rom_array(33712);
		when "1000001110110001" => data_out <= rom_array(33713);
		when "1000001110110010" => data_out <= rom_array(33714);
		when "1000001110110011" => data_out <= rom_array(33715);
		when "1000001110110100" => data_out <= rom_array(33716);
		when "1000001110110101" => data_out <= rom_array(33717);
		when "1000001110110110" => data_out <= rom_array(33718);
		when "1000001110110111" => data_out <= rom_array(33719);
		when "1000001110111000" => data_out <= rom_array(33720);
		when "1000001110111001" => data_out <= rom_array(33721);
		when "1000001110111010" => data_out <= rom_array(33722);
		when "1000001110111011" => data_out <= rom_array(33723);
		when "1000001110111100" => data_out <= rom_array(33724);
		when "1000001110111101" => data_out <= rom_array(33725);
		when "1000001110111110" => data_out <= rom_array(33726);
		when "1000001110111111" => data_out <= rom_array(33727);
		when "1000001111000000" => data_out <= rom_array(33728);
		when "1000001111000001" => data_out <= rom_array(33729);
		when "1000001111000010" => data_out <= rom_array(33730);
		when "1000001111000011" => data_out <= rom_array(33731);
		when "1000001111000100" => data_out <= rom_array(33732);
		when "1000001111000101" => data_out <= rom_array(33733);
		when "1000001111000110" => data_out <= rom_array(33734);
		when "1000001111000111" => data_out <= rom_array(33735);
		when "1000001111001000" => data_out <= rom_array(33736);
		when "1000001111001001" => data_out <= rom_array(33737);
		when "1000001111001010" => data_out <= rom_array(33738);
		when "1000001111001011" => data_out <= rom_array(33739);
		when "1000001111001100" => data_out <= rom_array(33740);
		when "1000001111001101" => data_out <= rom_array(33741);
		when "1000001111001110" => data_out <= rom_array(33742);
		when "1000001111001111" => data_out <= rom_array(33743);
		when "1000001111010000" => data_out <= rom_array(33744);
		when "1000001111010001" => data_out <= rom_array(33745);
		when "1000001111010010" => data_out <= rom_array(33746);
		when "1000001111010011" => data_out <= rom_array(33747);
		when "1000001111010100" => data_out <= rom_array(33748);
		when "1000001111010101" => data_out <= rom_array(33749);
		when "1000001111010110" => data_out <= rom_array(33750);
		when "1000001111010111" => data_out <= rom_array(33751);
		when "1000001111011000" => data_out <= rom_array(33752);
		when "1000001111011001" => data_out <= rom_array(33753);
		when "1000001111011010" => data_out <= rom_array(33754);
		when "1000001111011011" => data_out <= rom_array(33755);
		when "1000001111011100" => data_out <= rom_array(33756);
		when "1000001111011101" => data_out <= rom_array(33757);
		when "1000001111011110" => data_out <= rom_array(33758);
		when "1000001111011111" => data_out <= rom_array(33759);
		when "1000001111100000" => data_out <= rom_array(33760);
		when "1000001111100001" => data_out <= rom_array(33761);
		when "1000001111100010" => data_out <= rom_array(33762);
		when "1000001111100011" => data_out <= rom_array(33763);
		when "1000001111100100" => data_out <= rom_array(33764);
		when "1000001111100101" => data_out <= rom_array(33765);
		when "1000001111100110" => data_out <= rom_array(33766);
		when "1000001111100111" => data_out <= rom_array(33767);
		when "1000001111101000" => data_out <= rom_array(33768);
		when "1000001111101001" => data_out <= rom_array(33769);
		when "1000001111101010" => data_out <= rom_array(33770);
		when "1000001111101011" => data_out <= rom_array(33771);
		when "1000001111101100" => data_out <= rom_array(33772);
		when "1000001111101101" => data_out <= rom_array(33773);
		when "1000001111101110" => data_out <= rom_array(33774);
		when "1000001111101111" => data_out <= rom_array(33775);
		when "1000001111110000" => data_out <= rom_array(33776);
		when "1000001111110001" => data_out <= rom_array(33777);
		when "1000001111110010" => data_out <= rom_array(33778);
		when "1000001111110011" => data_out <= rom_array(33779);
		when "1000001111110100" => data_out <= rom_array(33780);
		when "1000001111110101" => data_out <= rom_array(33781);
		when "1000001111110110" => data_out <= rom_array(33782);
		when "1000001111110111" => data_out <= rom_array(33783);
		when "1000001111111000" => data_out <= rom_array(33784);
		when "1000001111111001" => data_out <= rom_array(33785);
		when "1000001111111010" => data_out <= rom_array(33786);
		when "1000001111111011" => data_out <= rom_array(33787);
		when "1000001111111100" => data_out <= rom_array(33788);
		when "1000001111111101" => data_out <= rom_array(33789);
		when "1000001111111110" => data_out <= rom_array(33790);
		when "1000001111111111" => data_out <= rom_array(33791);
		when "1000010000000000" => data_out <= rom_array(33792);
		when "1000010000000001" => data_out <= rom_array(33793);
		when "1000010000000010" => data_out <= rom_array(33794);
		when "1000010000000011" => data_out <= rom_array(33795);
		when "1000010000000100" => data_out <= rom_array(33796);
		when "1000010000000101" => data_out <= rom_array(33797);
		when "1000010000000110" => data_out <= rom_array(33798);
		when "1000010000000111" => data_out <= rom_array(33799);
		when "1000010000001000" => data_out <= rom_array(33800);
		when "1000010000001001" => data_out <= rom_array(33801);
		when "1000010000001010" => data_out <= rom_array(33802);
		when "1000010000001011" => data_out <= rom_array(33803);
		when "1000010000001100" => data_out <= rom_array(33804);
		when "1000010000001101" => data_out <= rom_array(33805);
		when "1000010000001110" => data_out <= rom_array(33806);
		when "1000010000001111" => data_out <= rom_array(33807);
		when "1000010000010000" => data_out <= rom_array(33808);
		when "1000010000010001" => data_out <= rom_array(33809);
		when "1000010000010010" => data_out <= rom_array(33810);
		when "1000010000010011" => data_out <= rom_array(33811);
		when "1000010000010100" => data_out <= rom_array(33812);
		when "1000010000010101" => data_out <= rom_array(33813);
		when "1000010000010110" => data_out <= rom_array(33814);
		when "1000010000010111" => data_out <= rom_array(33815);
		when "1000010000011000" => data_out <= rom_array(33816);
		when "1000010000011001" => data_out <= rom_array(33817);
		when "1000010000011010" => data_out <= rom_array(33818);
		when "1000010000011011" => data_out <= rom_array(33819);
		when "1000010000011100" => data_out <= rom_array(33820);
		when "1000010000011101" => data_out <= rom_array(33821);
		when "1000010000011110" => data_out <= rom_array(33822);
		when "1000010000011111" => data_out <= rom_array(33823);
		when "1000010000100000" => data_out <= rom_array(33824);
		when "1000010000100001" => data_out <= rom_array(33825);
		when "1000010000100010" => data_out <= rom_array(33826);
		when "1000010000100011" => data_out <= rom_array(33827);
		when "1000010000100100" => data_out <= rom_array(33828);
		when "1000010000100101" => data_out <= rom_array(33829);
		when "1000010000100110" => data_out <= rom_array(33830);
		when "1000010000100111" => data_out <= rom_array(33831);
		when "1000010000101000" => data_out <= rom_array(33832);
		when "1000010000101001" => data_out <= rom_array(33833);
		when "1000010000101010" => data_out <= rom_array(33834);
		when "1000010000101011" => data_out <= rom_array(33835);
		when "1000010000101100" => data_out <= rom_array(33836);
		when "1000010000101101" => data_out <= rom_array(33837);
		when "1000010000101110" => data_out <= rom_array(33838);
		when "1000010000101111" => data_out <= rom_array(33839);
		when "1000010000110000" => data_out <= rom_array(33840);
		when "1000010000110001" => data_out <= rom_array(33841);
		when "1000010000110010" => data_out <= rom_array(33842);
		when "1000010000110011" => data_out <= rom_array(33843);
		when "1000010000110100" => data_out <= rom_array(33844);
		when "1000010000110101" => data_out <= rom_array(33845);
		when "1000010000110110" => data_out <= rom_array(33846);
		when "1000010000110111" => data_out <= rom_array(33847);
		when "1000010000111000" => data_out <= rom_array(33848);
		when "1000010000111001" => data_out <= rom_array(33849);
		when "1000010000111010" => data_out <= rom_array(33850);
		when "1000010000111011" => data_out <= rom_array(33851);
		when "1000010000111100" => data_out <= rom_array(33852);
		when "1000010000111101" => data_out <= rom_array(33853);
		when "1000010000111110" => data_out <= rom_array(33854);
		when "1000010000111111" => data_out <= rom_array(33855);
		when "1000010001000000" => data_out <= rom_array(33856);
		when "1000010001000001" => data_out <= rom_array(33857);
		when "1000010001000010" => data_out <= rom_array(33858);
		when "1000010001000011" => data_out <= rom_array(33859);
		when "1000010001000100" => data_out <= rom_array(33860);
		when "1000010001000101" => data_out <= rom_array(33861);
		when "1000010001000110" => data_out <= rom_array(33862);
		when "1000010001000111" => data_out <= rom_array(33863);
		when "1000010001001000" => data_out <= rom_array(33864);
		when "1000010001001001" => data_out <= rom_array(33865);
		when "1000010001001010" => data_out <= rom_array(33866);
		when "1000010001001011" => data_out <= rom_array(33867);
		when "1000010001001100" => data_out <= rom_array(33868);
		when "1000010001001101" => data_out <= rom_array(33869);
		when "1000010001001110" => data_out <= rom_array(33870);
		when "1000010001001111" => data_out <= rom_array(33871);
		when "1000010001010000" => data_out <= rom_array(33872);
		when "1000010001010001" => data_out <= rom_array(33873);
		when "1000010001010010" => data_out <= rom_array(33874);
		when "1000010001010011" => data_out <= rom_array(33875);
		when "1000010001010100" => data_out <= rom_array(33876);
		when "1000010001010101" => data_out <= rom_array(33877);
		when "1000010001010110" => data_out <= rom_array(33878);
		when "1000010001010111" => data_out <= rom_array(33879);
		when "1000010001011000" => data_out <= rom_array(33880);
		when "1000010001011001" => data_out <= rom_array(33881);
		when "1000010001011010" => data_out <= rom_array(33882);
		when "1000010001011011" => data_out <= rom_array(33883);
		when "1000010001011100" => data_out <= rom_array(33884);
		when "1000010001011101" => data_out <= rom_array(33885);
		when "1000010001011110" => data_out <= rom_array(33886);
		when "1000010001011111" => data_out <= rom_array(33887);
		when "1000010001100000" => data_out <= rom_array(33888);
		when "1000010001100001" => data_out <= rom_array(33889);
		when "1000010001100010" => data_out <= rom_array(33890);
		when "1000010001100011" => data_out <= rom_array(33891);
		when "1000010001100100" => data_out <= rom_array(33892);
		when "1000010001100101" => data_out <= rom_array(33893);
		when "1000010001100110" => data_out <= rom_array(33894);
		when "1000010001100111" => data_out <= rom_array(33895);
		when "1000010001101000" => data_out <= rom_array(33896);
		when "1000010001101001" => data_out <= rom_array(33897);
		when "1000010001101010" => data_out <= rom_array(33898);
		when "1000010001101011" => data_out <= rom_array(33899);
		when "1000010001101100" => data_out <= rom_array(33900);
		when "1000010001101101" => data_out <= rom_array(33901);
		when "1000010001101110" => data_out <= rom_array(33902);
		when "1000010001101111" => data_out <= rom_array(33903);
		when "1000010001110000" => data_out <= rom_array(33904);
		when "1000010001110001" => data_out <= rom_array(33905);
		when "1000010001110010" => data_out <= rom_array(33906);
		when "1000010001110011" => data_out <= rom_array(33907);
		when "1000010001110100" => data_out <= rom_array(33908);
		when "1000010001110101" => data_out <= rom_array(33909);
		when "1000010001110110" => data_out <= rom_array(33910);
		when "1000010001110111" => data_out <= rom_array(33911);
		when "1000010001111000" => data_out <= rom_array(33912);
		when "1000010001111001" => data_out <= rom_array(33913);
		when "1000010001111010" => data_out <= rom_array(33914);
		when "1000010001111011" => data_out <= rom_array(33915);
		when "1000010001111100" => data_out <= rom_array(33916);
		when "1000010001111101" => data_out <= rom_array(33917);
		when "1000010001111110" => data_out <= rom_array(33918);
		when "1000010001111111" => data_out <= rom_array(33919);
		when "1000010010000000" => data_out <= rom_array(33920);
		when "1000010010000001" => data_out <= rom_array(33921);
		when "1000010010000010" => data_out <= rom_array(33922);
		when "1000010010000011" => data_out <= rom_array(33923);
		when "1000010010000100" => data_out <= rom_array(33924);
		when "1000010010000101" => data_out <= rom_array(33925);
		when "1000010010000110" => data_out <= rom_array(33926);
		when "1000010010000111" => data_out <= rom_array(33927);
		when "1000010010001000" => data_out <= rom_array(33928);
		when "1000010010001001" => data_out <= rom_array(33929);
		when "1000010010001010" => data_out <= rom_array(33930);
		when "1000010010001011" => data_out <= rom_array(33931);
		when "1000010010001100" => data_out <= rom_array(33932);
		when "1000010010001101" => data_out <= rom_array(33933);
		when "1000010010001110" => data_out <= rom_array(33934);
		when "1000010010001111" => data_out <= rom_array(33935);
		when "1000010010010000" => data_out <= rom_array(33936);
		when "1000010010010001" => data_out <= rom_array(33937);
		when "1000010010010010" => data_out <= rom_array(33938);
		when "1000010010010011" => data_out <= rom_array(33939);
		when "1000010010010100" => data_out <= rom_array(33940);
		when "1000010010010101" => data_out <= rom_array(33941);
		when "1000010010010110" => data_out <= rom_array(33942);
		when "1000010010010111" => data_out <= rom_array(33943);
		when "1000010010011000" => data_out <= rom_array(33944);
		when "1000010010011001" => data_out <= rom_array(33945);
		when "1000010010011010" => data_out <= rom_array(33946);
		when "1000010010011011" => data_out <= rom_array(33947);
		when "1000010010011100" => data_out <= rom_array(33948);
		when "1000010010011101" => data_out <= rom_array(33949);
		when "1000010010011110" => data_out <= rom_array(33950);
		when "1000010010011111" => data_out <= rom_array(33951);
		when "1000010010100000" => data_out <= rom_array(33952);
		when "1000010010100001" => data_out <= rom_array(33953);
		when "1000010010100010" => data_out <= rom_array(33954);
		when "1000010010100011" => data_out <= rom_array(33955);
		when "1000010010100100" => data_out <= rom_array(33956);
		when "1000010010100101" => data_out <= rom_array(33957);
		when "1000010010100110" => data_out <= rom_array(33958);
		when "1000010010100111" => data_out <= rom_array(33959);
		when "1000010010101000" => data_out <= rom_array(33960);
		when "1000010010101001" => data_out <= rom_array(33961);
		when "1000010010101010" => data_out <= rom_array(33962);
		when "1000010010101011" => data_out <= rom_array(33963);
		when "1000010010101100" => data_out <= rom_array(33964);
		when "1000010010101101" => data_out <= rom_array(33965);
		when "1000010010101110" => data_out <= rom_array(33966);
		when "1000010010101111" => data_out <= rom_array(33967);
		when "1000010010110000" => data_out <= rom_array(33968);
		when "1000010010110001" => data_out <= rom_array(33969);
		when "1000010010110010" => data_out <= rom_array(33970);
		when "1000010010110011" => data_out <= rom_array(33971);
		when "1000010010110100" => data_out <= rom_array(33972);
		when "1000010010110101" => data_out <= rom_array(33973);
		when "1000010010110110" => data_out <= rom_array(33974);
		when "1000010010110111" => data_out <= rom_array(33975);
		when "1000010010111000" => data_out <= rom_array(33976);
		when "1000010010111001" => data_out <= rom_array(33977);
		when "1000010010111010" => data_out <= rom_array(33978);
		when "1000010010111011" => data_out <= rom_array(33979);
		when "1000010010111100" => data_out <= rom_array(33980);
		when "1000010010111101" => data_out <= rom_array(33981);
		when "1000010010111110" => data_out <= rom_array(33982);
		when "1000010010111111" => data_out <= rom_array(33983);
		when "1000010011000000" => data_out <= rom_array(33984);
		when "1000010011000001" => data_out <= rom_array(33985);
		when "1000010011000010" => data_out <= rom_array(33986);
		when "1000010011000011" => data_out <= rom_array(33987);
		when "1000010011000100" => data_out <= rom_array(33988);
		when "1000010011000101" => data_out <= rom_array(33989);
		when "1000010011000110" => data_out <= rom_array(33990);
		when "1000010011000111" => data_out <= rom_array(33991);
		when "1000010011001000" => data_out <= rom_array(33992);
		when "1000010011001001" => data_out <= rom_array(33993);
		when "1000010011001010" => data_out <= rom_array(33994);
		when "1000010011001011" => data_out <= rom_array(33995);
		when "1000010011001100" => data_out <= rom_array(33996);
		when "1000010011001101" => data_out <= rom_array(33997);
		when "1000010011001110" => data_out <= rom_array(33998);
		when "1000010011001111" => data_out <= rom_array(33999);
		when "1000010011010000" => data_out <= rom_array(34000);
		when "1000010011010001" => data_out <= rom_array(34001);
		when "1000010011010010" => data_out <= rom_array(34002);
		when "1000010011010011" => data_out <= rom_array(34003);
		when "1000010011010100" => data_out <= rom_array(34004);
		when "1000010011010101" => data_out <= rom_array(34005);
		when "1000010011010110" => data_out <= rom_array(34006);
		when "1000010011010111" => data_out <= rom_array(34007);
		when "1000010011011000" => data_out <= rom_array(34008);
		when "1000010011011001" => data_out <= rom_array(34009);
		when "1000010011011010" => data_out <= rom_array(34010);
		when "1000010011011011" => data_out <= rom_array(34011);
		when "1000010011011100" => data_out <= rom_array(34012);
		when "1000010011011101" => data_out <= rom_array(34013);
		when "1000010011011110" => data_out <= rom_array(34014);
		when "1000010011011111" => data_out <= rom_array(34015);
		when "1000010011100000" => data_out <= rom_array(34016);
		when "1000010011100001" => data_out <= rom_array(34017);
		when "1000010011100010" => data_out <= rom_array(34018);
		when "1000010011100011" => data_out <= rom_array(34019);
		when "1000010011100100" => data_out <= rom_array(34020);
		when "1000010011100101" => data_out <= rom_array(34021);
		when "1000010011100110" => data_out <= rom_array(34022);
		when "1000010011100111" => data_out <= rom_array(34023);
		when "1000010011101000" => data_out <= rom_array(34024);
		when "1000010011101001" => data_out <= rom_array(34025);
		when "1000010011101010" => data_out <= rom_array(34026);
		when "1000010011101011" => data_out <= rom_array(34027);
		when "1000010011101100" => data_out <= rom_array(34028);
		when "1000010011101101" => data_out <= rom_array(34029);
		when "1000010011101110" => data_out <= rom_array(34030);
		when "1000010011101111" => data_out <= rom_array(34031);
		when "1000010011110000" => data_out <= rom_array(34032);
		when "1000010011110001" => data_out <= rom_array(34033);
		when "1000010011110010" => data_out <= rom_array(34034);
		when "1000010011110011" => data_out <= rom_array(34035);
		when "1000010011110100" => data_out <= rom_array(34036);
		when "1000010011110101" => data_out <= rom_array(34037);
		when "1000010011110110" => data_out <= rom_array(34038);
		when "1000010011110111" => data_out <= rom_array(34039);
		when "1000010011111000" => data_out <= rom_array(34040);
		when "1000010011111001" => data_out <= rom_array(34041);
		when "1000010011111010" => data_out <= rom_array(34042);
		when "1000010011111011" => data_out <= rom_array(34043);
		when "1000010011111100" => data_out <= rom_array(34044);
		when "1000010011111101" => data_out <= rom_array(34045);
		when "1000010011111110" => data_out <= rom_array(34046);
		when "1000010011111111" => data_out <= rom_array(34047);
		when "1000010100000000" => data_out <= rom_array(34048);
		when "1000010100000001" => data_out <= rom_array(34049);
		when "1000010100000010" => data_out <= rom_array(34050);
		when "1000010100000011" => data_out <= rom_array(34051);
		when "1000010100000100" => data_out <= rom_array(34052);
		when "1000010100000101" => data_out <= rom_array(34053);
		when "1000010100000110" => data_out <= rom_array(34054);
		when "1000010100000111" => data_out <= rom_array(34055);
		when "1000010100001000" => data_out <= rom_array(34056);
		when "1000010100001001" => data_out <= rom_array(34057);
		when "1000010100001010" => data_out <= rom_array(34058);
		when "1000010100001011" => data_out <= rom_array(34059);
		when "1000010100001100" => data_out <= rom_array(34060);
		when "1000010100001101" => data_out <= rom_array(34061);
		when "1000010100001110" => data_out <= rom_array(34062);
		when "1000010100001111" => data_out <= rom_array(34063);
		when "1000010100010000" => data_out <= rom_array(34064);
		when "1000010100010001" => data_out <= rom_array(34065);
		when "1000010100010010" => data_out <= rom_array(34066);
		when "1000010100010011" => data_out <= rom_array(34067);
		when "1000010100010100" => data_out <= rom_array(34068);
		when "1000010100010101" => data_out <= rom_array(34069);
		when "1000010100010110" => data_out <= rom_array(34070);
		when "1000010100010111" => data_out <= rom_array(34071);
		when "1000010100011000" => data_out <= rom_array(34072);
		when "1000010100011001" => data_out <= rom_array(34073);
		when "1000010100011010" => data_out <= rom_array(34074);
		when "1000010100011011" => data_out <= rom_array(34075);
		when "1000010100011100" => data_out <= rom_array(34076);
		when "1000010100011101" => data_out <= rom_array(34077);
		when "1000010100011110" => data_out <= rom_array(34078);
		when "1000010100011111" => data_out <= rom_array(34079);
		when "1000010100100000" => data_out <= rom_array(34080);
		when "1000010100100001" => data_out <= rom_array(34081);
		when "1000010100100010" => data_out <= rom_array(34082);
		when "1000010100100011" => data_out <= rom_array(34083);
		when "1000010100100100" => data_out <= rom_array(34084);
		when "1000010100100101" => data_out <= rom_array(34085);
		when "1000010100100110" => data_out <= rom_array(34086);
		when "1000010100100111" => data_out <= rom_array(34087);
		when "1000010100101000" => data_out <= rom_array(34088);
		when "1000010100101001" => data_out <= rom_array(34089);
		when "1000010100101010" => data_out <= rom_array(34090);
		when "1000010100101011" => data_out <= rom_array(34091);
		when "1000010100101100" => data_out <= rom_array(34092);
		when "1000010100101101" => data_out <= rom_array(34093);
		when "1000010100101110" => data_out <= rom_array(34094);
		when "1000010100101111" => data_out <= rom_array(34095);
		when "1000010100110000" => data_out <= rom_array(34096);
		when "1000010100110001" => data_out <= rom_array(34097);
		when "1000010100110010" => data_out <= rom_array(34098);
		when "1000010100110011" => data_out <= rom_array(34099);
		when "1000010100110100" => data_out <= rom_array(34100);
		when "1000010100110101" => data_out <= rom_array(34101);
		when "1000010100110110" => data_out <= rom_array(34102);
		when "1000010100110111" => data_out <= rom_array(34103);
		when "1000010100111000" => data_out <= rom_array(34104);
		when "1000010100111001" => data_out <= rom_array(34105);
		when "1000010100111010" => data_out <= rom_array(34106);
		when "1000010100111011" => data_out <= rom_array(34107);
		when "1000010100111100" => data_out <= rom_array(34108);
		when "1000010100111101" => data_out <= rom_array(34109);
		when "1000010100111110" => data_out <= rom_array(34110);
		when "1000010100111111" => data_out <= rom_array(34111);
		when "1000010101000000" => data_out <= rom_array(34112);
		when "1000010101000001" => data_out <= rom_array(34113);
		when "1000010101000010" => data_out <= rom_array(34114);
		when "1000010101000011" => data_out <= rom_array(34115);
		when "1000010101000100" => data_out <= rom_array(34116);
		when "1000010101000101" => data_out <= rom_array(34117);
		when "1000010101000110" => data_out <= rom_array(34118);
		when "1000010101000111" => data_out <= rom_array(34119);
		when "1000010101001000" => data_out <= rom_array(34120);
		when "1000010101001001" => data_out <= rom_array(34121);
		when "1000010101001010" => data_out <= rom_array(34122);
		when "1000010101001011" => data_out <= rom_array(34123);
		when "1000010101001100" => data_out <= rom_array(34124);
		when "1000010101001101" => data_out <= rom_array(34125);
		when "1000010101001110" => data_out <= rom_array(34126);
		when "1000010101001111" => data_out <= rom_array(34127);
		when "1000010101010000" => data_out <= rom_array(34128);
		when "1000010101010001" => data_out <= rom_array(34129);
		when "1000010101010010" => data_out <= rom_array(34130);
		when "1000010101010011" => data_out <= rom_array(34131);
		when "1000010101010100" => data_out <= rom_array(34132);
		when "1000010101010101" => data_out <= rom_array(34133);
		when "1000010101010110" => data_out <= rom_array(34134);
		when "1000010101010111" => data_out <= rom_array(34135);
		when "1000010101011000" => data_out <= rom_array(34136);
		when "1000010101011001" => data_out <= rom_array(34137);
		when "1000010101011010" => data_out <= rom_array(34138);
		when "1000010101011011" => data_out <= rom_array(34139);
		when "1000010101011100" => data_out <= rom_array(34140);
		when "1000010101011101" => data_out <= rom_array(34141);
		when "1000010101011110" => data_out <= rom_array(34142);
		when "1000010101011111" => data_out <= rom_array(34143);
		when "1000010101100000" => data_out <= rom_array(34144);
		when "1000010101100001" => data_out <= rom_array(34145);
		when "1000010101100010" => data_out <= rom_array(34146);
		when "1000010101100011" => data_out <= rom_array(34147);
		when "1000010101100100" => data_out <= rom_array(34148);
		when "1000010101100101" => data_out <= rom_array(34149);
		when "1000010101100110" => data_out <= rom_array(34150);
		when "1000010101100111" => data_out <= rom_array(34151);
		when "1000010101101000" => data_out <= rom_array(34152);
		when "1000010101101001" => data_out <= rom_array(34153);
		when "1000010101101010" => data_out <= rom_array(34154);
		when "1000010101101011" => data_out <= rom_array(34155);
		when "1000010101101100" => data_out <= rom_array(34156);
		when "1000010101101101" => data_out <= rom_array(34157);
		when "1000010101101110" => data_out <= rom_array(34158);
		when "1000010101101111" => data_out <= rom_array(34159);
		when "1000010101110000" => data_out <= rom_array(34160);
		when "1000010101110001" => data_out <= rom_array(34161);
		when "1000010101110010" => data_out <= rom_array(34162);
		when "1000010101110011" => data_out <= rom_array(34163);
		when "1000010101110100" => data_out <= rom_array(34164);
		when "1000010101110101" => data_out <= rom_array(34165);
		when "1000010101110110" => data_out <= rom_array(34166);
		when "1000010101110111" => data_out <= rom_array(34167);
		when "1000010101111000" => data_out <= rom_array(34168);
		when "1000010101111001" => data_out <= rom_array(34169);
		when "1000010101111010" => data_out <= rom_array(34170);
		when "1000010101111011" => data_out <= rom_array(34171);
		when "1000010101111100" => data_out <= rom_array(34172);
		when "1000010101111101" => data_out <= rom_array(34173);
		when "1000010101111110" => data_out <= rom_array(34174);
		when "1000010101111111" => data_out <= rom_array(34175);
		when "1000010110000000" => data_out <= rom_array(34176);
		when "1000010110000001" => data_out <= rom_array(34177);
		when "1000010110000010" => data_out <= rom_array(34178);
		when "1000010110000011" => data_out <= rom_array(34179);
		when "1000010110000100" => data_out <= rom_array(34180);
		when "1000010110000101" => data_out <= rom_array(34181);
		when "1000010110000110" => data_out <= rom_array(34182);
		when "1000010110000111" => data_out <= rom_array(34183);
		when "1000010110001000" => data_out <= rom_array(34184);
		when "1000010110001001" => data_out <= rom_array(34185);
		when "1000010110001010" => data_out <= rom_array(34186);
		when "1000010110001011" => data_out <= rom_array(34187);
		when "1000010110001100" => data_out <= rom_array(34188);
		when "1000010110001101" => data_out <= rom_array(34189);
		when "1000010110001110" => data_out <= rom_array(34190);
		when "1000010110001111" => data_out <= rom_array(34191);
		when "1000010110010000" => data_out <= rom_array(34192);
		when "1000010110010001" => data_out <= rom_array(34193);
		when "1000010110010010" => data_out <= rom_array(34194);
		when "1000010110010011" => data_out <= rom_array(34195);
		when "1000010110010100" => data_out <= rom_array(34196);
		when "1000010110010101" => data_out <= rom_array(34197);
		when "1000010110010110" => data_out <= rom_array(34198);
		when "1000010110010111" => data_out <= rom_array(34199);
		when "1000010110011000" => data_out <= rom_array(34200);
		when "1000010110011001" => data_out <= rom_array(34201);
		when "1000010110011010" => data_out <= rom_array(34202);
		when "1000010110011011" => data_out <= rom_array(34203);
		when "1000010110011100" => data_out <= rom_array(34204);
		when "1000010110011101" => data_out <= rom_array(34205);
		when "1000010110011110" => data_out <= rom_array(34206);
		when "1000010110011111" => data_out <= rom_array(34207);
		when "1000010110100000" => data_out <= rom_array(34208);
		when "1000010110100001" => data_out <= rom_array(34209);
		when "1000010110100010" => data_out <= rom_array(34210);
		when "1000010110100011" => data_out <= rom_array(34211);
		when "1000010110100100" => data_out <= rom_array(34212);
		when "1000010110100101" => data_out <= rom_array(34213);
		when "1000010110100110" => data_out <= rom_array(34214);
		when "1000010110100111" => data_out <= rom_array(34215);
		when "1000010110101000" => data_out <= rom_array(34216);
		when "1000010110101001" => data_out <= rom_array(34217);
		when "1000010110101010" => data_out <= rom_array(34218);
		when "1000010110101011" => data_out <= rom_array(34219);
		when "1000010110101100" => data_out <= rom_array(34220);
		when "1000010110101101" => data_out <= rom_array(34221);
		when "1000010110101110" => data_out <= rom_array(34222);
		when "1000010110101111" => data_out <= rom_array(34223);
		when "1000010110110000" => data_out <= rom_array(34224);
		when "1000010110110001" => data_out <= rom_array(34225);
		when "1000010110110010" => data_out <= rom_array(34226);
		when "1000010110110011" => data_out <= rom_array(34227);
		when "1000010110110100" => data_out <= rom_array(34228);
		when "1000010110110101" => data_out <= rom_array(34229);
		when "1000010110110110" => data_out <= rom_array(34230);
		when "1000010110110111" => data_out <= rom_array(34231);
		when "1000010110111000" => data_out <= rom_array(34232);
		when "1000010110111001" => data_out <= rom_array(34233);
		when "1000010110111010" => data_out <= rom_array(34234);
		when "1000010110111011" => data_out <= rom_array(34235);
		when "1000010110111100" => data_out <= rom_array(34236);
		when "1000010110111101" => data_out <= rom_array(34237);
		when "1000010110111110" => data_out <= rom_array(34238);
		when "1000010110111111" => data_out <= rom_array(34239);
		when "1000010111000000" => data_out <= rom_array(34240);
		when "1000010111000001" => data_out <= rom_array(34241);
		when "1000010111000010" => data_out <= rom_array(34242);
		when "1000010111000011" => data_out <= rom_array(34243);
		when "1000010111000100" => data_out <= rom_array(34244);
		when "1000010111000101" => data_out <= rom_array(34245);
		when "1000010111000110" => data_out <= rom_array(34246);
		when "1000010111000111" => data_out <= rom_array(34247);
		when "1000010111001000" => data_out <= rom_array(34248);
		when "1000010111001001" => data_out <= rom_array(34249);
		when "1000010111001010" => data_out <= rom_array(34250);
		when "1000010111001011" => data_out <= rom_array(34251);
		when "1000010111001100" => data_out <= rom_array(34252);
		when "1000010111001101" => data_out <= rom_array(34253);
		when "1000010111001110" => data_out <= rom_array(34254);
		when "1000010111001111" => data_out <= rom_array(34255);
		when "1000010111010000" => data_out <= rom_array(34256);
		when "1000010111010001" => data_out <= rom_array(34257);
		when "1000010111010010" => data_out <= rom_array(34258);
		when "1000010111010011" => data_out <= rom_array(34259);
		when "1000010111010100" => data_out <= rom_array(34260);
		when "1000010111010101" => data_out <= rom_array(34261);
		when "1000010111010110" => data_out <= rom_array(34262);
		when "1000010111010111" => data_out <= rom_array(34263);
		when "1000010111011000" => data_out <= rom_array(34264);
		when "1000010111011001" => data_out <= rom_array(34265);
		when "1000010111011010" => data_out <= rom_array(34266);
		when "1000010111011011" => data_out <= rom_array(34267);
		when "1000010111011100" => data_out <= rom_array(34268);
		when "1000010111011101" => data_out <= rom_array(34269);
		when "1000010111011110" => data_out <= rom_array(34270);
		when "1000010111011111" => data_out <= rom_array(34271);
		when "1000010111100000" => data_out <= rom_array(34272);
		when "1000010111100001" => data_out <= rom_array(34273);
		when "1000010111100010" => data_out <= rom_array(34274);
		when "1000010111100011" => data_out <= rom_array(34275);
		when "1000010111100100" => data_out <= rom_array(34276);
		when "1000010111100101" => data_out <= rom_array(34277);
		when "1000010111100110" => data_out <= rom_array(34278);
		when "1000010111100111" => data_out <= rom_array(34279);
		when "1000010111101000" => data_out <= rom_array(34280);
		when "1000010111101001" => data_out <= rom_array(34281);
		when "1000010111101010" => data_out <= rom_array(34282);
		when "1000010111101011" => data_out <= rom_array(34283);
		when "1000010111101100" => data_out <= rom_array(34284);
		when "1000010111101101" => data_out <= rom_array(34285);
		when "1000010111101110" => data_out <= rom_array(34286);
		when "1000010111101111" => data_out <= rom_array(34287);
		when "1000010111110000" => data_out <= rom_array(34288);
		when "1000010111110001" => data_out <= rom_array(34289);
		when "1000010111110010" => data_out <= rom_array(34290);
		when "1000010111110011" => data_out <= rom_array(34291);
		when "1000010111110100" => data_out <= rom_array(34292);
		when "1000010111110101" => data_out <= rom_array(34293);
		when "1000010111110110" => data_out <= rom_array(34294);
		when "1000010111110111" => data_out <= rom_array(34295);
		when "1000010111111000" => data_out <= rom_array(34296);
		when "1000010111111001" => data_out <= rom_array(34297);
		when "1000010111111010" => data_out <= rom_array(34298);
		when "1000010111111011" => data_out <= rom_array(34299);
		when "1000010111111100" => data_out <= rom_array(34300);
		when "1000010111111101" => data_out <= rom_array(34301);
		when "1000010111111110" => data_out <= rom_array(34302);
		when "1000010111111111" => data_out <= rom_array(34303);
		when "1000011000000000" => data_out <= rom_array(34304);
		when "1000011000000001" => data_out <= rom_array(34305);
		when "1000011000000010" => data_out <= rom_array(34306);
		when "1000011000000011" => data_out <= rom_array(34307);
		when "1000011000000100" => data_out <= rom_array(34308);
		when "1000011000000101" => data_out <= rom_array(34309);
		when "1000011000000110" => data_out <= rom_array(34310);
		when "1000011000000111" => data_out <= rom_array(34311);
		when "1000011000001000" => data_out <= rom_array(34312);
		when "1000011000001001" => data_out <= rom_array(34313);
		when "1000011000001010" => data_out <= rom_array(34314);
		when "1000011000001011" => data_out <= rom_array(34315);
		when "1000011000001100" => data_out <= rom_array(34316);
		when "1000011000001101" => data_out <= rom_array(34317);
		when "1000011000001110" => data_out <= rom_array(34318);
		when "1000011000001111" => data_out <= rom_array(34319);
		when "1000011000010000" => data_out <= rom_array(34320);
		when "1000011000010001" => data_out <= rom_array(34321);
		when "1000011000010010" => data_out <= rom_array(34322);
		when "1000011000010011" => data_out <= rom_array(34323);
		when "1000011000010100" => data_out <= rom_array(34324);
		when "1000011000010101" => data_out <= rom_array(34325);
		when "1000011000010110" => data_out <= rom_array(34326);
		when "1000011000010111" => data_out <= rom_array(34327);
		when "1000011000011000" => data_out <= rom_array(34328);
		when "1000011000011001" => data_out <= rom_array(34329);
		when "1000011000011010" => data_out <= rom_array(34330);
		when "1000011000011011" => data_out <= rom_array(34331);
		when "1000011000011100" => data_out <= rom_array(34332);
		when "1000011000011101" => data_out <= rom_array(34333);
		when "1000011000011110" => data_out <= rom_array(34334);
		when "1000011000011111" => data_out <= rom_array(34335);
		when "1000011000100000" => data_out <= rom_array(34336);
		when "1000011000100001" => data_out <= rom_array(34337);
		when "1000011000100010" => data_out <= rom_array(34338);
		when "1000011000100011" => data_out <= rom_array(34339);
		when "1000011000100100" => data_out <= rom_array(34340);
		when "1000011000100101" => data_out <= rom_array(34341);
		when "1000011000100110" => data_out <= rom_array(34342);
		when "1000011000100111" => data_out <= rom_array(34343);
		when "1000011000101000" => data_out <= rom_array(34344);
		when "1000011000101001" => data_out <= rom_array(34345);
		when "1000011000101010" => data_out <= rom_array(34346);
		when "1000011000101011" => data_out <= rom_array(34347);
		when "1000011000101100" => data_out <= rom_array(34348);
		when "1000011000101101" => data_out <= rom_array(34349);
		when "1000011000101110" => data_out <= rom_array(34350);
		when "1000011000101111" => data_out <= rom_array(34351);
		when "1000011000110000" => data_out <= rom_array(34352);
		when "1000011000110001" => data_out <= rom_array(34353);
		when "1000011000110010" => data_out <= rom_array(34354);
		when "1000011000110011" => data_out <= rom_array(34355);
		when "1000011000110100" => data_out <= rom_array(34356);
		when "1000011000110101" => data_out <= rom_array(34357);
		when "1000011000110110" => data_out <= rom_array(34358);
		when "1000011000110111" => data_out <= rom_array(34359);
		when "1000011000111000" => data_out <= rom_array(34360);
		when "1000011000111001" => data_out <= rom_array(34361);
		when "1000011000111010" => data_out <= rom_array(34362);
		when "1000011000111011" => data_out <= rom_array(34363);
		when "1000011000111100" => data_out <= rom_array(34364);
		when "1000011000111101" => data_out <= rom_array(34365);
		when "1000011000111110" => data_out <= rom_array(34366);
		when "1000011000111111" => data_out <= rom_array(34367);
		when "1000011001000000" => data_out <= rom_array(34368);
		when "1000011001000001" => data_out <= rom_array(34369);
		when "1000011001000010" => data_out <= rom_array(34370);
		when "1000011001000011" => data_out <= rom_array(34371);
		when "1000011001000100" => data_out <= rom_array(34372);
		when "1000011001000101" => data_out <= rom_array(34373);
		when "1000011001000110" => data_out <= rom_array(34374);
		when "1000011001000111" => data_out <= rom_array(34375);
		when "1000011001001000" => data_out <= rom_array(34376);
		when "1000011001001001" => data_out <= rom_array(34377);
		when "1000011001001010" => data_out <= rom_array(34378);
		when "1000011001001011" => data_out <= rom_array(34379);
		when "1000011001001100" => data_out <= rom_array(34380);
		when "1000011001001101" => data_out <= rom_array(34381);
		when "1000011001001110" => data_out <= rom_array(34382);
		when "1000011001001111" => data_out <= rom_array(34383);
		when "1000011001010000" => data_out <= rom_array(34384);
		when "1000011001010001" => data_out <= rom_array(34385);
		when "1000011001010010" => data_out <= rom_array(34386);
		when "1000011001010011" => data_out <= rom_array(34387);
		when "1000011001010100" => data_out <= rom_array(34388);
		when "1000011001010101" => data_out <= rom_array(34389);
		when "1000011001010110" => data_out <= rom_array(34390);
		when "1000011001010111" => data_out <= rom_array(34391);
		when "1000011001011000" => data_out <= rom_array(34392);
		when "1000011001011001" => data_out <= rom_array(34393);
		when "1000011001011010" => data_out <= rom_array(34394);
		when "1000011001011011" => data_out <= rom_array(34395);
		when "1000011001011100" => data_out <= rom_array(34396);
		when "1000011001011101" => data_out <= rom_array(34397);
		when "1000011001011110" => data_out <= rom_array(34398);
		when "1000011001011111" => data_out <= rom_array(34399);
		when "1000011001100000" => data_out <= rom_array(34400);
		when "1000011001100001" => data_out <= rom_array(34401);
		when "1000011001100010" => data_out <= rom_array(34402);
		when "1000011001100011" => data_out <= rom_array(34403);
		when "1000011001100100" => data_out <= rom_array(34404);
		when "1000011001100101" => data_out <= rom_array(34405);
		when "1000011001100110" => data_out <= rom_array(34406);
		when "1000011001100111" => data_out <= rom_array(34407);
		when "1000011001101000" => data_out <= rom_array(34408);
		when "1000011001101001" => data_out <= rom_array(34409);
		when "1000011001101010" => data_out <= rom_array(34410);
		when "1000011001101011" => data_out <= rom_array(34411);
		when "1000011001101100" => data_out <= rom_array(34412);
		when "1000011001101101" => data_out <= rom_array(34413);
		when "1000011001101110" => data_out <= rom_array(34414);
		when "1000011001101111" => data_out <= rom_array(34415);
		when "1000011001110000" => data_out <= rom_array(34416);
		when "1000011001110001" => data_out <= rom_array(34417);
		when "1000011001110010" => data_out <= rom_array(34418);
		when "1000011001110011" => data_out <= rom_array(34419);
		when "1000011001110100" => data_out <= rom_array(34420);
		when "1000011001110101" => data_out <= rom_array(34421);
		when "1000011001110110" => data_out <= rom_array(34422);
		when "1000011001110111" => data_out <= rom_array(34423);
		when "1000011001111000" => data_out <= rom_array(34424);
		when "1000011001111001" => data_out <= rom_array(34425);
		when "1000011001111010" => data_out <= rom_array(34426);
		when "1000011001111011" => data_out <= rom_array(34427);
		when "1000011001111100" => data_out <= rom_array(34428);
		when "1000011001111101" => data_out <= rom_array(34429);
		when "1000011001111110" => data_out <= rom_array(34430);
		when "1000011001111111" => data_out <= rom_array(34431);
		when "1000011010000000" => data_out <= rom_array(34432);
		when "1000011010000001" => data_out <= rom_array(34433);
		when "1000011010000010" => data_out <= rom_array(34434);
		when "1000011010000011" => data_out <= rom_array(34435);
		when "1000011010000100" => data_out <= rom_array(34436);
		when "1000011010000101" => data_out <= rom_array(34437);
		when "1000011010000110" => data_out <= rom_array(34438);
		when "1000011010000111" => data_out <= rom_array(34439);
		when "1000011010001000" => data_out <= rom_array(34440);
		when "1000011010001001" => data_out <= rom_array(34441);
		when "1000011010001010" => data_out <= rom_array(34442);
		when "1000011010001011" => data_out <= rom_array(34443);
		when "1000011010001100" => data_out <= rom_array(34444);
		when "1000011010001101" => data_out <= rom_array(34445);
		when "1000011010001110" => data_out <= rom_array(34446);
		when "1000011010001111" => data_out <= rom_array(34447);
		when "1000011010010000" => data_out <= rom_array(34448);
		when "1000011010010001" => data_out <= rom_array(34449);
		when "1000011010010010" => data_out <= rom_array(34450);
		when "1000011010010011" => data_out <= rom_array(34451);
		when "1000011010010100" => data_out <= rom_array(34452);
		when "1000011010010101" => data_out <= rom_array(34453);
		when "1000011010010110" => data_out <= rom_array(34454);
		when "1000011010010111" => data_out <= rom_array(34455);
		when "1000011010011000" => data_out <= rom_array(34456);
		when "1000011010011001" => data_out <= rom_array(34457);
		when "1000011010011010" => data_out <= rom_array(34458);
		when "1000011010011011" => data_out <= rom_array(34459);
		when "1000011010011100" => data_out <= rom_array(34460);
		when "1000011010011101" => data_out <= rom_array(34461);
		when "1000011010011110" => data_out <= rom_array(34462);
		when "1000011010011111" => data_out <= rom_array(34463);
		when "1000011010100000" => data_out <= rom_array(34464);
		when "1000011010100001" => data_out <= rom_array(34465);
		when "1000011010100010" => data_out <= rom_array(34466);
		when "1000011010100011" => data_out <= rom_array(34467);
		when "1000011010100100" => data_out <= rom_array(34468);
		when "1000011010100101" => data_out <= rom_array(34469);
		when "1000011010100110" => data_out <= rom_array(34470);
		when "1000011010100111" => data_out <= rom_array(34471);
		when "1000011010101000" => data_out <= rom_array(34472);
		when "1000011010101001" => data_out <= rom_array(34473);
		when "1000011010101010" => data_out <= rom_array(34474);
		when "1000011010101011" => data_out <= rom_array(34475);
		when "1000011010101100" => data_out <= rom_array(34476);
		when "1000011010101101" => data_out <= rom_array(34477);
		when "1000011010101110" => data_out <= rom_array(34478);
		when "1000011010101111" => data_out <= rom_array(34479);
		when "1000011010110000" => data_out <= rom_array(34480);
		when "1000011010110001" => data_out <= rom_array(34481);
		when "1000011010110010" => data_out <= rom_array(34482);
		when "1000011010110011" => data_out <= rom_array(34483);
		when "1000011010110100" => data_out <= rom_array(34484);
		when "1000011010110101" => data_out <= rom_array(34485);
		when "1000011010110110" => data_out <= rom_array(34486);
		when "1000011010110111" => data_out <= rom_array(34487);
		when "1000011010111000" => data_out <= rom_array(34488);
		when "1000011010111001" => data_out <= rom_array(34489);
		when "1000011010111010" => data_out <= rom_array(34490);
		when "1000011010111011" => data_out <= rom_array(34491);
		when "1000011010111100" => data_out <= rom_array(34492);
		when "1000011010111101" => data_out <= rom_array(34493);
		when "1000011010111110" => data_out <= rom_array(34494);
		when "1000011010111111" => data_out <= rom_array(34495);
		when "1000011011000000" => data_out <= rom_array(34496);
		when "1000011011000001" => data_out <= rom_array(34497);
		when "1000011011000010" => data_out <= rom_array(34498);
		when "1000011011000011" => data_out <= rom_array(34499);
		when "1000011011000100" => data_out <= rom_array(34500);
		when "1000011011000101" => data_out <= rom_array(34501);
		when "1000011011000110" => data_out <= rom_array(34502);
		when "1000011011000111" => data_out <= rom_array(34503);
		when "1000011011001000" => data_out <= rom_array(34504);
		when "1000011011001001" => data_out <= rom_array(34505);
		when "1000011011001010" => data_out <= rom_array(34506);
		when "1000011011001011" => data_out <= rom_array(34507);
		when "1000011011001100" => data_out <= rom_array(34508);
		when "1000011011001101" => data_out <= rom_array(34509);
		when "1000011011001110" => data_out <= rom_array(34510);
		when "1000011011001111" => data_out <= rom_array(34511);
		when "1000011011010000" => data_out <= rom_array(34512);
		when "1000011011010001" => data_out <= rom_array(34513);
		when "1000011011010010" => data_out <= rom_array(34514);
		when "1000011011010011" => data_out <= rom_array(34515);
		when "1000011011010100" => data_out <= rom_array(34516);
		when "1000011011010101" => data_out <= rom_array(34517);
		when "1000011011010110" => data_out <= rom_array(34518);
		when "1000011011010111" => data_out <= rom_array(34519);
		when "1000011011011000" => data_out <= rom_array(34520);
		when "1000011011011001" => data_out <= rom_array(34521);
		when "1000011011011010" => data_out <= rom_array(34522);
		when "1000011011011011" => data_out <= rom_array(34523);
		when "1000011011011100" => data_out <= rom_array(34524);
		when "1000011011011101" => data_out <= rom_array(34525);
		when "1000011011011110" => data_out <= rom_array(34526);
		when "1000011011011111" => data_out <= rom_array(34527);
		when "1000011011100000" => data_out <= rom_array(34528);
		when "1000011011100001" => data_out <= rom_array(34529);
		when "1000011011100010" => data_out <= rom_array(34530);
		when "1000011011100011" => data_out <= rom_array(34531);
		when "1000011011100100" => data_out <= rom_array(34532);
		when "1000011011100101" => data_out <= rom_array(34533);
		when "1000011011100110" => data_out <= rom_array(34534);
		when "1000011011100111" => data_out <= rom_array(34535);
		when "1000011011101000" => data_out <= rom_array(34536);
		when "1000011011101001" => data_out <= rom_array(34537);
		when "1000011011101010" => data_out <= rom_array(34538);
		when "1000011011101011" => data_out <= rom_array(34539);
		when "1000011011101100" => data_out <= rom_array(34540);
		when "1000011011101101" => data_out <= rom_array(34541);
		when "1000011011101110" => data_out <= rom_array(34542);
		when "1000011011101111" => data_out <= rom_array(34543);
		when "1000011011110000" => data_out <= rom_array(34544);
		when "1000011011110001" => data_out <= rom_array(34545);
		when "1000011011110010" => data_out <= rom_array(34546);
		when "1000011011110011" => data_out <= rom_array(34547);
		when "1000011011110100" => data_out <= rom_array(34548);
		when "1000011011110101" => data_out <= rom_array(34549);
		when "1000011011110110" => data_out <= rom_array(34550);
		when "1000011011110111" => data_out <= rom_array(34551);
		when "1000011011111000" => data_out <= rom_array(34552);
		when "1000011011111001" => data_out <= rom_array(34553);
		when "1000011011111010" => data_out <= rom_array(34554);
		when "1000011011111011" => data_out <= rom_array(34555);
		when "1000011011111100" => data_out <= rom_array(34556);
		when "1000011011111101" => data_out <= rom_array(34557);
		when "1000011011111110" => data_out <= rom_array(34558);
		when "1000011011111111" => data_out <= rom_array(34559);
		when "1000011100000000" => data_out <= rom_array(34560);
		when "1000011100000001" => data_out <= rom_array(34561);
		when "1000011100000010" => data_out <= rom_array(34562);
		when "1000011100000011" => data_out <= rom_array(34563);
		when "1000011100000100" => data_out <= rom_array(34564);
		when "1000011100000101" => data_out <= rom_array(34565);
		when "1000011100000110" => data_out <= rom_array(34566);
		when "1000011100000111" => data_out <= rom_array(34567);
		when "1000011100001000" => data_out <= rom_array(34568);
		when "1000011100001001" => data_out <= rom_array(34569);
		when "1000011100001010" => data_out <= rom_array(34570);
		when "1000011100001011" => data_out <= rom_array(34571);
		when "1000011100001100" => data_out <= rom_array(34572);
		when "1000011100001101" => data_out <= rom_array(34573);
		when "1000011100001110" => data_out <= rom_array(34574);
		when "1000011100001111" => data_out <= rom_array(34575);
		when "1000011100010000" => data_out <= rom_array(34576);
		when "1000011100010001" => data_out <= rom_array(34577);
		when "1000011100010010" => data_out <= rom_array(34578);
		when "1000011100010011" => data_out <= rom_array(34579);
		when "1000011100010100" => data_out <= rom_array(34580);
		when "1000011100010101" => data_out <= rom_array(34581);
		when "1000011100010110" => data_out <= rom_array(34582);
		when "1000011100010111" => data_out <= rom_array(34583);
		when "1000011100011000" => data_out <= rom_array(34584);
		when "1000011100011001" => data_out <= rom_array(34585);
		when "1000011100011010" => data_out <= rom_array(34586);
		when "1000011100011011" => data_out <= rom_array(34587);
		when "1000011100011100" => data_out <= rom_array(34588);
		when "1000011100011101" => data_out <= rom_array(34589);
		when "1000011100011110" => data_out <= rom_array(34590);
		when "1000011100011111" => data_out <= rom_array(34591);
		when "1000011100100000" => data_out <= rom_array(34592);
		when "1000011100100001" => data_out <= rom_array(34593);
		when "1000011100100010" => data_out <= rom_array(34594);
		when "1000011100100011" => data_out <= rom_array(34595);
		when "1000011100100100" => data_out <= rom_array(34596);
		when "1000011100100101" => data_out <= rom_array(34597);
		when "1000011100100110" => data_out <= rom_array(34598);
		when "1000011100100111" => data_out <= rom_array(34599);
		when "1000011100101000" => data_out <= rom_array(34600);
		when "1000011100101001" => data_out <= rom_array(34601);
		when "1000011100101010" => data_out <= rom_array(34602);
		when "1000011100101011" => data_out <= rom_array(34603);
		when "1000011100101100" => data_out <= rom_array(34604);
		when "1000011100101101" => data_out <= rom_array(34605);
		when "1000011100101110" => data_out <= rom_array(34606);
		when "1000011100101111" => data_out <= rom_array(34607);
		when "1000011100110000" => data_out <= rom_array(34608);
		when "1000011100110001" => data_out <= rom_array(34609);
		when "1000011100110010" => data_out <= rom_array(34610);
		when "1000011100110011" => data_out <= rom_array(34611);
		when "1000011100110100" => data_out <= rom_array(34612);
		when "1000011100110101" => data_out <= rom_array(34613);
		when "1000011100110110" => data_out <= rom_array(34614);
		when "1000011100110111" => data_out <= rom_array(34615);
		when "1000011100111000" => data_out <= rom_array(34616);
		when "1000011100111001" => data_out <= rom_array(34617);
		when "1000011100111010" => data_out <= rom_array(34618);
		when "1000011100111011" => data_out <= rom_array(34619);
		when "1000011100111100" => data_out <= rom_array(34620);
		when "1000011100111101" => data_out <= rom_array(34621);
		when "1000011100111110" => data_out <= rom_array(34622);
		when "1000011100111111" => data_out <= rom_array(34623);
		when "1000011101000000" => data_out <= rom_array(34624);
		when "1000011101000001" => data_out <= rom_array(34625);
		when "1000011101000010" => data_out <= rom_array(34626);
		when "1000011101000011" => data_out <= rom_array(34627);
		when "1000011101000100" => data_out <= rom_array(34628);
		when "1000011101000101" => data_out <= rom_array(34629);
		when "1000011101000110" => data_out <= rom_array(34630);
		when "1000011101000111" => data_out <= rom_array(34631);
		when "1000011101001000" => data_out <= rom_array(34632);
		when "1000011101001001" => data_out <= rom_array(34633);
		when "1000011101001010" => data_out <= rom_array(34634);
		when "1000011101001011" => data_out <= rom_array(34635);
		when "1000011101001100" => data_out <= rom_array(34636);
		when "1000011101001101" => data_out <= rom_array(34637);
		when "1000011101001110" => data_out <= rom_array(34638);
		when "1000011101001111" => data_out <= rom_array(34639);
		when "1000011101010000" => data_out <= rom_array(34640);
		when "1000011101010001" => data_out <= rom_array(34641);
		when "1000011101010010" => data_out <= rom_array(34642);
		when "1000011101010011" => data_out <= rom_array(34643);
		when "1000011101010100" => data_out <= rom_array(34644);
		when "1000011101010101" => data_out <= rom_array(34645);
		when "1000011101010110" => data_out <= rom_array(34646);
		when "1000011101010111" => data_out <= rom_array(34647);
		when "1000011101011000" => data_out <= rom_array(34648);
		when "1000011101011001" => data_out <= rom_array(34649);
		when "1000011101011010" => data_out <= rom_array(34650);
		when "1000011101011011" => data_out <= rom_array(34651);
		when "1000011101011100" => data_out <= rom_array(34652);
		when "1000011101011101" => data_out <= rom_array(34653);
		when "1000011101011110" => data_out <= rom_array(34654);
		when "1000011101011111" => data_out <= rom_array(34655);
		when "1000011101100000" => data_out <= rom_array(34656);
		when "1000011101100001" => data_out <= rom_array(34657);
		when "1000011101100010" => data_out <= rom_array(34658);
		when "1000011101100011" => data_out <= rom_array(34659);
		when "1000011101100100" => data_out <= rom_array(34660);
		when "1000011101100101" => data_out <= rom_array(34661);
		when "1000011101100110" => data_out <= rom_array(34662);
		when "1000011101100111" => data_out <= rom_array(34663);
		when "1000011101101000" => data_out <= rom_array(34664);
		when "1000011101101001" => data_out <= rom_array(34665);
		when "1000011101101010" => data_out <= rom_array(34666);
		when "1000011101101011" => data_out <= rom_array(34667);
		when "1000011101101100" => data_out <= rom_array(34668);
		when "1000011101101101" => data_out <= rom_array(34669);
		when "1000011101101110" => data_out <= rom_array(34670);
		when "1000011101101111" => data_out <= rom_array(34671);
		when "1000011101110000" => data_out <= rom_array(34672);
		when "1000011101110001" => data_out <= rom_array(34673);
		when "1000011101110010" => data_out <= rom_array(34674);
		when "1000011101110011" => data_out <= rom_array(34675);
		when "1000011101110100" => data_out <= rom_array(34676);
		when "1000011101110101" => data_out <= rom_array(34677);
		when "1000011101110110" => data_out <= rom_array(34678);
		when "1000011101110111" => data_out <= rom_array(34679);
		when "1000011101111000" => data_out <= rom_array(34680);
		when "1000011101111001" => data_out <= rom_array(34681);
		when "1000011101111010" => data_out <= rom_array(34682);
		when "1000011101111011" => data_out <= rom_array(34683);
		when "1000011101111100" => data_out <= rom_array(34684);
		when "1000011101111101" => data_out <= rom_array(34685);
		when "1000011101111110" => data_out <= rom_array(34686);
		when "1000011101111111" => data_out <= rom_array(34687);
		when "1000011110000000" => data_out <= rom_array(34688);
		when "1000011110000001" => data_out <= rom_array(34689);
		when "1000011110000010" => data_out <= rom_array(34690);
		when "1000011110000011" => data_out <= rom_array(34691);
		when "1000011110000100" => data_out <= rom_array(34692);
		when "1000011110000101" => data_out <= rom_array(34693);
		when "1000011110000110" => data_out <= rom_array(34694);
		when "1000011110000111" => data_out <= rom_array(34695);
		when "1000011110001000" => data_out <= rom_array(34696);
		when "1000011110001001" => data_out <= rom_array(34697);
		when "1000011110001010" => data_out <= rom_array(34698);
		when "1000011110001011" => data_out <= rom_array(34699);
		when "1000011110001100" => data_out <= rom_array(34700);
		when "1000011110001101" => data_out <= rom_array(34701);
		when "1000011110001110" => data_out <= rom_array(34702);
		when "1000011110001111" => data_out <= rom_array(34703);
		when "1000011110010000" => data_out <= rom_array(34704);
		when "1000011110010001" => data_out <= rom_array(34705);
		when "1000011110010010" => data_out <= rom_array(34706);
		when "1000011110010011" => data_out <= rom_array(34707);
		when "1000011110010100" => data_out <= rom_array(34708);
		when "1000011110010101" => data_out <= rom_array(34709);
		when "1000011110010110" => data_out <= rom_array(34710);
		when "1000011110010111" => data_out <= rom_array(34711);
		when "1000011110011000" => data_out <= rom_array(34712);
		when "1000011110011001" => data_out <= rom_array(34713);
		when "1000011110011010" => data_out <= rom_array(34714);
		when "1000011110011011" => data_out <= rom_array(34715);
		when "1000011110011100" => data_out <= rom_array(34716);
		when "1000011110011101" => data_out <= rom_array(34717);
		when "1000011110011110" => data_out <= rom_array(34718);
		when "1000011110011111" => data_out <= rom_array(34719);
		when "1000011110100000" => data_out <= rom_array(34720);
		when "1000011110100001" => data_out <= rom_array(34721);
		when "1000011110100010" => data_out <= rom_array(34722);
		when "1000011110100011" => data_out <= rom_array(34723);
		when "1000011110100100" => data_out <= rom_array(34724);
		when "1000011110100101" => data_out <= rom_array(34725);
		when "1000011110100110" => data_out <= rom_array(34726);
		when "1000011110100111" => data_out <= rom_array(34727);
		when "1000011110101000" => data_out <= rom_array(34728);
		when "1000011110101001" => data_out <= rom_array(34729);
		when "1000011110101010" => data_out <= rom_array(34730);
		when "1000011110101011" => data_out <= rom_array(34731);
		when "1000011110101100" => data_out <= rom_array(34732);
		when "1000011110101101" => data_out <= rom_array(34733);
		when "1000011110101110" => data_out <= rom_array(34734);
		when "1000011110101111" => data_out <= rom_array(34735);
		when "1000011110110000" => data_out <= rom_array(34736);
		when "1000011110110001" => data_out <= rom_array(34737);
		when "1000011110110010" => data_out <= rom_array(34738);
		when "1000011110110011" => data_out <= rom_array(34739);
		when "1000011110110100" => data_out <= rom_array(34740);
		when "1000011110110101" => data_out <= rom_array(34741);
		when "1000011110110110" => data_out <= rom_array(34742);
		when "1000011110110111" => data_out <= rom_array(34743);
		when "1000011110111000" => data_out <= rom_array(34744);
		when "1000011110111001" => data_out <= rom_array(34745);
		when "1000011110111010" => data_out <= rom_array(34746);
		when "1000011110111011" => data_out <= rom_array(34747);
		when "1000011110111100" => data_out <= rom_array(34748);
		when "1000011110111101" => data_out <= rom_array(34749);
		when "1000011110111110" => data_out <= rom_array(34750);
		when "1000011110111111" => data_out <= rom_array(34751);
		when "1000011111000000" => data_out <= rom_array(34752);
		when "1000011111000001" => data_out <= rom_array(34753);
		when "1000011111000010" => data_out <= rom_array(34754);
		when "1000011111000011" => data_out <= rom_array(34755);
		when "1000011111000100" => data_out <= rom_array(34756);
		when "1000011111000101" => data_out <= rom_array(34757);
		when "1000011111000110" => data_out <= rom_array(34758);
		when "1000011111000111" => data_out <= rom_array(34759);
		when "1000011111001000" => data_out <= rom_array(34760);
		when "1000011111001001" => data_out <= rom_array(34761);
		when "1000011111001010" => data_out <= rom_array(34762);
		when "1000011111001011" => data_out <= rom_array(34763);
		when "1000011111001100" => data_out <= rom_array(34764);
		when "1000011111001101" => data_out <= rom_array(34765);
		when "1000011111001110" => data_out <= rom_array(34766);
		when "1000011111001111" => data_out <= rom_array(34767);
		when "1000011111010000" => data_out <= rom_array(34768);
		when "1000011111010001" => data_out <= rom_array(34769);
		when "1000011111010010" => data_out <= rom_array(34770);
		when "1000011111010011" => data_out <= rom_array(34771);
		when "1000011111010100" => data_out <= rom_array(34772);
		when "1000011111010101" => data_out <= rom_array(34773);
		when "1000011111010110" => data_out <= rom_array(34774);
		when "1000011111010111" => data_out <= rom_array(34775);
		when "1000011111011000" => data_out <= rom_array(34776);
		when "1000011111011001" => data_out <= rom_array(34777);
		when "1000011111011010" => data_out <= rom_array(34778);
		when "1000011111011011" => data_out <= rom_array(34779);
		when "1000011111011100" => data_out <= rom_array(34780);
		when "1000011111011101" => data_out <= rom_array(34781);
		when "1000011111011110" => data_out <= rom_array(34782);
		when "1000011111011111" => data_out <= rom_array(34783);
		when "1000011111100000" => data_out <= rom_array(34784);
		when "1000011111100001" => data_out <= rom_array(34785);
		when "1000011111100010" => data_out <= rom_array(34786);
		when "1000011111100011" => data_out <= rom_array(34787);
		when "1000011111100100" => data_out <= rom_array(34788);
		when "1000011111100101" => data_out <= rom_array(34789);
		when "1000011111100110" => data_out <= rom_array(34790);
		when "1000011111100111" => data_out <= rom_array(34791);
		when "1000011111101000" => data_out <= rom_array(34792);
		when "1000011111101001" => data_out <= rom_array(34793);
		when "1000011111101010" => data_out <= rom_array(34794);
		when "1000011111101011" => data_out <= rom_array(34795);
		when "1000011111101100" => data_out <= rom_array(34796);
		when "1000011111101101" => data_out <= rom_array(34797);
		when "1000011111101110" => data_out <= rom_array(34798);
		when "1000011111101111" => data_out <= rom_array(34799);
		when "1000011111110000" => data_out <= rom_array(34800);
		when "1000011111110001" => data_out <= rom_array(34801);
		when "1000011111110010" => data_out <= rom_array(34802);
		when "1000011111110011" => data_out <= rom_array(34803);
		when "1000011111110100" => data_out <= rom_array(34804);
		when "1000011111110101" => data_out <= rom_array(34805);
		when "1000011111110110" => data_out <= rom_array(34806);
		when "1000011111110111" => data_out <= rom_array(34807);
		when "1000011111111000" => data_out <= rom_array(34808);
		when "1000011111111001" => data_out <= rom_array(34809);
		when "1000011111111010" => data_out <= rom_array(34810);
		when "1000011111111011" => data_out <= rom_array(34811);
		when "1000011111111100" => data_out <= rom_array(34812);
		when "1000011111111101" => data_out <= rom_array(34813);
		when "1000011111111110" => data_out <= rom_array(34814);
		when "1000011111111111" => data_out <= rom_array(34815);
		when "1000100000000000" => data_out <= rom_array(34816);
		when "1000100000000001" => data_out <= rom_array(34817);
		when "1000100000000010" => data_out <= rom_array(34818);
		when "1000100000000011" => data_out <= rom_array(34819);
		when "1000100000000100" => data_out <= rom_array(34820);
		when "1000100000000101" => data_out <= rom_array(34821);
		when "1000100000000110" => data_out <= rom_array(34822);
		when "1000100000000111" => data_out <= rom_array(34823);
		when "1000100000001000" => data_out <= rom_array(34824);
		when "1000100000001001" => data_out <= rom_array(34825);
		when "1000100000001010" => data_out <= rom_array(34826);
		when "1000100000001011" => data_out <= rom_array(34827);
		when "1000100000001100" => data_out <= rom_array(34828);
		when "1000100000001101" => data_out <= rom_array(34829);
		when "1000100000001110" => data_out <= rom_array(34830);
		when "1000100000001111" => data_out <= rom_array(34831);
		when "1000100000010000" => data_out <= rom_array(34832);
		when "1000100000010001" => data_out <= rom_array(34833);
		when "1000100000010010" => data_out <= rom_array(34834);
		when "1000100000010011" => data_out <= rom_array(34835);
		when "1000100000010100" => data_out <= rom_array(34836);
		when "1000100000010101" => data_out <= rom_array(34837);
		when "1000100000010110" => data_out <= rom_array(34838);
		when "1000100000010111" => data_out <= rom_array(34839);
		when "1000100000011000" => data_out <= rom_array(34840);
		when "1000100000011001" => data_out <= rom_array(34841);
		when "1000100000011010" => data_out <= rom_array(34842);
		when "1000100000011011" => data_out <= rom_array(34843);
		when "1000100000011100" => data_out <= rom_array(34844);
		when "1000100000011101" => data_out <= rom_array(34845);
		when "1000100000011110" => data_out <= rom_array(34846);
		when "1000100000011111" => data_out <= rom_array(34847);
		when "1000100000100000" => data_out <= rom_array(34848);
		when "1000100000100001" => data_out <= rom_array(34849);
		when "1000100000100010" => data_out <= rom_array(34850);
		when "1000100000100011" => data_out <= rom_array(34851);
		when "1000100000100100" => data_out <= rom_array(34852);
		when "1000100000100101" => data_out <= rom_array(34853);
		when "1000100000100110" => data_out <= rom_array(34854);
		when "1000100000100111" => data_out <= rom_array(34855);
		when "1000100000101000" => data_out <= rom_array(34856);
		when "1000100000101001" => data_out <= rom_array(34857);
		when "1000100000101010" => data_out <= rom_array(34858);
		when "1000100000101011" => data_out <= rom_array(34859);
		when "1000100000101100" => data_out <= rom_array(34860);
		when "1000100000101101" => data_out <= rom_array(34861);
		when "1000100000101110" => data_out <= rom_array(34862);
		when "1000100000101111" => data_out <= rom_array(34863);
		when "1000100000110000" => data_out <= rom_array(34864);
		when "1000100000110001" => data_out <= rom_array(34865);
		when "1000100000110010" => data_out <= rom_array(34866);
		when "1000100000110011" => data_out <= rom_array(34867);
		when "1000100000110100" => data_out <= rom_array(34868);
		when "1000100000110101" => data_out <= rom_array(34869);
		when "1000100000110110" => data_out <= rom_array(34870);
		when "1000100000110111" => data_out <= rom_array(34871);
		when "1000100000111000" => data_out <= rom_array(34872);
		when "1000100000111001" => data_out <= rom_array(34873);
		when "1000100000111010" => data_out <= rom_array(34874);
		when "1000100000111011" => data_out <= rom_array(34875);
		when "1000100000111100" => data_out <= rom_array(34876);
		when "1000100000111101" => data_out <= rom_array(34877);
		when "1000100000111110" => data_out <= rom_array(34878);
		when "1000100000111111" => data_out <= rom_array(34879);
		when "1000100001000000" => data_out <= rom_array(34880);
		when "1000100001000001" => data_out <= rom_array(34881);
		when "1000100001000010" => data_out <= rom_array(34882);
		when "1000100001000011" => data_out <= rom_array(34883);
		when "1000100001000100" => data_out <= rom_array(34884);
		when "1000100001000101" => data_out <= rom_array(34885);
		when "1000100001000110" => data_out <= rom_array(34886);
		when "1000100001000111" => data_out <= rom_array(34887);
		when "1000100001001000" => data_out <= rom_array(34888);
		when "1000100001001001" => data_out <= rom_array(34889);
		when "1000100001001010" => data_out <= rom_array(34890);
		when "1000100001001011" => data_out <= rom_array(34891);
		when "1000100001001100" => data_out <= rom_array(34892);
		when "1000100001001101" => data_out <= rom_array(34893);
		when "1000100001001110" => data_out <= rom_array(34894);
		when "1000100001001111" => data_out <= rom_array(34895);
		when "1000100001010000" => data_out <= rom_array(34896);
		when "1000100001010001" => data_out <= rom_array(34897);
		when "1000100001010010" => data_out <= rom_array(34898);
		when "1000100001010011" => data_out <= rom_array(34899);
		when "1000100001010100" => data_out <= rom_array(34900);
		when "1000100001010101" => data_out <= rom_array(34901);
		when "1000100001010110" => data_out <= rom_array(34902);
		when "1000100001010111" => data_out <= rom_array(34903);
		when "1000100001011000" => data_out <= rom_array(34904);
		when "1000100001011001" => data_out <= rom_array(34905);
		when "1000100001011010" => data_out <= rom_array(34906);
		when "1000100001011011" => data_out <= rom_array(34907);
		when "1000100001011100" => data_out <= rom_array(34908);
		when "1000100001011101" => data_out <= rom_array(34909);
		when "1000100001011110" => data_out <= rom_array(34910);
		when "1000100001011111" => data_out <= rom_array(34911);
		when "1000100001100000" => data_out <= rom_array(34912);
		when "1000100001100001" => data_out <= rom_array(34913);
		when "1000100001100010" => data_out <= rom_array(34914);
		when "1000100001100011" => data_out <= rom_array(34915);
		when "1000100001100100" => data_out <= rom_array(34916);
		when "1000100001100101" => data_out <= rom_array(34917);
		when "1000100001100110" => data_out <= rom_array(34918);
		when "1000100001100111" => data_out <= rom_array(34919);
		when "1000100001101000" => data_out <= rom_array(34920);
		when "1000100001101001" => data_out <= rom_array(34921);
		when "1000100001101010" => data_out <= rom_array(34922);
		when "1000100001101011" => data_out <= rom_array(34923);
		when "1000100001101100" => data_out <= rom_array(34924);
		when "1000100001101101" => data_out <= rom_array(34925);
		when "1000100001101110" => data_out <= rom_array(34926);
		when "1000100001101111" => data_out <= rom_array(34927);
		when "1000100001110000" => data_out <= rom_array(34928);
		when "1000100001110001" => data_out <= rom_array(34929);
		when "1000100001110010" => data_out <= rom_array(34930);
		when "1000100001110011" => data_out <= rom_array(34931);
		when "1000100001110100" => data_out <= rom_array(34932);
		when "1000100001110101" => data_out <= rom_array(34933);
		when "1000100001110110" => data_out <= rom_array(34934);
		when "1000100001110111" => data_out <= rom_array(34935);
		when "1000100001111000" => data_out <= rom_array(34936);
		when "1000100001111001" => data_out <= rom_array(34937);
		when "1000100001111010" => data_out <= rom_array(34938);
		when "1000100001111011" => data_out <= rom_array(34939);
		when "1000100001111100" => data_out <= rom_array(34940);
		when "1000100001111101" => data_out <= rom_array(34941);
		when "1000100001111110" => data_out <= rom_array(34942);
		when "1000100001111111" => data_out <= rom_array(34943);
		when "1000100010000000" => data_out <= rom_array(34944);
		when "1000100010000001" => data_out <= rom_array(34945);
		when "1000100010000010" => data_out <= rom_array(34946);
		when "1000100010000011" => data_out <= rom_array(34947);
		when "1000100010000100" => data_out <= rom_array(34948);
		when "1000100010000101" => data_out <= rom_array(34949);
		when "1000100010000110" => data_out <= rom_array(34950);
		when "1000100010000111" => data_out <= rom_array(34951);
		when "1000100010001000" => data_out <= rom_array(34952);
		when "1000100010001001" => data_out <= rom_array(34953);
		when "1000100010001010" => data_out <= rom_array(34954);
		when "1000100010001011" => data_out <= rom_array(34955);
		when "1000100010001100" => data_out <= rom_array(34956);
		when "1000100010001101" => data_out <= rom_array(34957);
		when "1000100010001110" => data_out <= rom_array(34958);
		when "1000100010001111" => data_out <= rom_array(34959);
		when "1000100010010000" => data_out <= rom_array(34960);
		when "1000100010010001" => data_out <= rom_array(34961);
		when "1000100010010010" => data_out <= rom_array(34962);
		when "1000100010010011" => data_out <= rom_array(34963);
		when "1000100010010100" => data_out <= rom_array(34964);
		when "1000100010010101" => data_out <= rom_array(34965);
		when "1000100010010110" => data_out <= rom_array(34966);
		when "1000100010010111" => data_out <= rom_array(34967);
		when "1000100010011000" => data_out <= rom_array(34968);
		when "1000100010011001" => data_out <= rom_array(34969);
		when "1000100010011010" => data_out <= rom_array(34970);
		when "1000100010011011" => data_out <= rom_array(34971);
		when "1000100010011100" => data_out <= rom_array(34972);
		when "1000100010011101" => data_out <= rom_array(34973);
		when "1000100010011110" => data_out <= rom_array(34974);
		when "1000100010011111" => data_out <= rom_array(34975);
		when "1000100010100000" => data_out <= rom_array(34976);
		when "1000100010100001" => data_out <= rom_array(34977);
		when "1000100010100010" => data_out <= rom_array(34978);
		when "1000100010100011" => data_out <= rom_array(34979);
		when "1000100010100100" => data_out <= rom_array(34980);
		when "1000100010100101" => data_out <= rom_array(34981);
		when "1000100010100110" => data_out <= rom_array(34982);
		when "1000100010100111" => data_out <= rom_array(34983);
		when "1000100010101000" => data_out <= rom_array(34984);
		when "1000100010101001" => data_out <= rom_array(34985);
		when "1000100010101010" => data_out <= rom_array(34986);
		when "1000100010101011" => data_out <= rom_array(34987);
		when "1000100010101100" => data_out <= rom_array(34988);
		when "1000100010101101" => data_out <= rom_array(34989);
		when "1000100010101110" => data_out <= rom_array(34990);
		when "1000100010101111" => data_out <= rom_array(34991);
		when "1000100010110000" => data_out <= rom_array(34992);
		when "1000100010110001" => data_out <= rom_array(34993);
		when "1000100010110010" => data_out <= rom_array(34994);
		when "1000100010110011" => data_out <= rom_array(34995);
		when "1000100010110100" => data_out <= rom_array(34996);
		when "1000100010110101" => data_out <= rom_array(34997);
		when "1000100010110110" => data_out <= rom_array(34998);
		when "1000100010110111" => data_out <= rom_array(34999);
		when "1000100010111000" => data_out <= rom_array(35000);
		when "1000100010111001" => data_out <= rom_array(35001);
		when "1000100010111010" => data_out <= rom_array(35002);
		when "1000100010111011" => data_out <= rom_array(35003);
		when "1000100010111100" => data_out <= rom_array(35004);
		when "1000100010111101" => data_out <= rom_array(35005);
		when "1000100010111110" => data_out <= rom_array(35006);
		when "1000100010111111" => data_out <= rom_array(35007);
		when "1000100011000000" => data_out <= rom_array(35008);
		when "1000100011000001" => data_out <= rom_array(35009);
		when "1000100011000010" => data_out <= rom_array(35010);
		when "1000100011000011" => data_out <= rom_array(35011);
		when "1000100011000100" => data_out <= rom_array(35012);
		when "1000100011000101" => data_out <= rom_array(35013);
		when "1000100011000110" => data_out <= rom_array(35014);
		when "1000100011000111" => data_out <= rom_array(35015);
		when "1000100011001000" => data_out <= rom_array(35016);
		when "1000100011001001" => data_out <= rom_array(35017);
		when "1000100011001010" => data_out <= rom_array(35018);
		when "1000100011001011" => data_out <= rom_array(35019);
		when "1000100011001100" => data_out <= rom_array(35020);
		when "1000100011001101" => data_out <= rom_array(35021);
		when "1000100011001110" => data_out <= rom_array(35022);
		when "1000100011001111" => data_out <= rom_array(35023);
		when "1000100011010000" => data_out <= rom_array(35024);
		when "1000100011010001" => data_out <= rom_array(35025);
		when "1000100011010010" => data_out <= rom_array(35026);
		when "1000100011010011" => data_out <= rom_array(35027);
		when "1000100011010100" => data_out <= rom_array(35028);
		when "1000100011010101" => data_out <= rom_array(35029);
		when "1000100011010110" => data_out <= rom_array(35030);
		when "1000100011010111" => data_out <= rom_array(35031);
		when "1000100011011000" => data_out <= rom_array(35032);
		when "1000100011011001" => data_out <= rom_array(35033);
		when "1000100011011010" => data_out <= rom_array(35034);
		when "1000100011011011" => data_out <= rom_array(35035);
		when "1000100011011100" => data_out <= rom_array(35036);
		when "1000100011011101" => data_out <= rom_array(35037);
		when "1000100011011110" => data_out <= rom_array(35038);
		when "1000100011011111" => data_out <= rom_array(35039);
		when "1000100011100000" => data_out <= rom_array(35040);
		when "1000100011100001" => data_out <= rom_array(35041);
		when "1000100011100010" => data_out <= rom_array(35042);
		when "1000100011100011" => data_out <= rom_array(35043);
		when "1000100011100100" => data_out <= rom_array(35044);
		when "1000100011100101" => data_out <= rom_array(35045);
		when "1000100011100110" => data_out <= rom_array(35046);
		when "1000100011100111" => data_out <= rom_array(35047);
		when "1000100011101000" => data_out <= rom_array(35048);
		when "1000100011101001" => data_out <= rom_array(35049);
		when "1000100011101010" => data_out <= rom_array(35050);
		when "1000100011101011" => data_out <= rom_array(35051);
		when "1000100011101100" => data_out <= rom_array(35052);
		when "1000100011101101" => data_out <= rom_array(35053);
		when "1000100011101110" => data_out <= rom_array(35054);
		when "1000100011101111" => data_out <= rom_array(35055);
		when "1000100011110000" => data_out <= rom_array(35056);
		when "1000100011110001" => data_out <= rom_array(35057);
		when "1000100011110010" => data_out <= rom_array(35058);
		when "1000100011110011" => data_out <= rom_array(35059);
		when "1000100011110100" => data_out <= rom_array(35060);
		when "1000100011110101" => data_out <= rom_array(35061);
		when "1000100011110110" => data_out <= rom_array(35062);
		when "1000100011110111" => data_out <= rom_array(35063);
		when "1000100011111000" => data_out <= rom_array(35064);
		when "1000100011111001" => data_out <= rom_array(35065);
		when "1000100011111010" => data_out <= rom_array(35066);
		when "1000100011111011" => data_out <= rom_array(35067);
		when "1000100011111100" => data_out <= rom_array(35068);
		when "1000100011111101" => data_out <= rom_array(35069);
		when "1000100011111110" => data_out <= rom_array(35070);
		when "1000100011111111" => data_out <= rom_array(35071);
		when "1000100100000000" => data_out <= rom_array(35072);
		when "1000100100000001" => data_out <= rom_array(35073);
		when "1000100100000010" => data_out <= rom_array(35074);
		when "1000100100000011" => data_out <= rom_array(35075);
		when "1000100100000100" => data_out <= rom_array(35076);
		when "1000100100000101" => data_out <= rom_array(35077);
		when "1000100100000110" => data_out <= rom_array(35078);
		when "1000100100000111" => data_out <= rom_array(35079);
		when "1000100100001000" => data_out <= rom_array(35080);
		when "1000100100001001" => data_out <= rom_array(35081);
		when "1000100100001010" => data_out <= rom_array(35082);
		when "1000100100001011" => data_out <= rom_array(35083);
		when "1000100100001100" => data_out <= rom_array(35084);
		when "1000100100001101" => data_out <= rom_array(35085);
		when "1000100100001110" => data_out <= rom_array(35086);
		when "1000100100001111" => data_out <= rom_array(35087);
		when "1000100100010000" => data_out <= rom_array(35088);
		when "1000100100010001" => data_out <= rom_array(35089);
		when "1000100100010010" => data_out <= rom_array(35090);
		when "1000100100010011" => data_out <= rom_array(35091);
		when "1000100100010100" => data_out <= rom_array(35092);
		when "1000100100010101" => data_out <= rom_array(35093);
		when "1000100100010110" => data_out <= rom_array(35094);
		when "1000100100010111" => data_out <= rom_array(35095);
		when "1000100100011000" => data_out <= rom_array(35096);
		when "1000100100011001" => data_out <= rom_array(35097);
		when "1000100100011010" => data_out <= rom_array(35098);
		when "1000100100011011" => data_out <= rom_array(35099);
		when "1000100100011100" => data_out <= rom_array(35100);
		when "1000100100011101" => data_out <= rom_array(35101);
		when "1000100100011110" => data_out <= rom_array(35102);
		when "1000100100011111" => data_out <= rom_array(35103);
		when "1000100100100000" => data_out <= rom_array(35104);
		when "1000100100100001" => data_out <= rom_array(35105);
		when "1000100100100010" => data_out <= rom_array(35106);
		when "1000100100100011" => data_out <= rom_array(35107);
		when "1000100100100100" => data_out <= rom_array(35108);
		when "1000100100100101" => data_out <= rom_array(35109);
		when "1000100100100110" => data_out <= rom_array(35110);
		when "1000100100100111" => data_out <= rom_array(35111);
		when "1000100100101000" => data_out <= rom_array(35112);
		when "1000100100101001" => data_out <= rom_array(35113);
		when "1000100100101010" => data_out <= rom_array(35114);
		when "1000100100101011" => data_out <= rom_array(35115);
		when "1000100100101100" => data_out <= rom_array(35116);
		when "1000100100101101" => data_out <= rom_array(35117);
		when "1000100100101110" => data_out <= rom_array(35118);
		when "1000100100101111" => data_out <= rom_array(35119);
		when "1000100100110000" => data_out <= rom_array(35120);
		when "1000100100110001" => data_out <= rom_array(35121);
		when "1000100100110010" => data_out <= rom_array(35122);
		when "1000100100110011" => data_out <= rom_array(35123);
		when "1000100100110100" => data_out <= rom_array(35124);
		when "1000100100110101" => data_out <= rom_array(35125);
		when "1000100100110110" => data_out <= rom_array(35126);
		when "1000100100110111" => data_out <= rom_array(35127);
		when "1000100100111000" => data_out <= rom_array(35128);
		when "1000100100111001" => data_out <= rom_array(35129);
		when "1000100100111010" => data_out <= rom_array(35130);
		when "1000100100111011" => data_out <= rom_array(35131);
		when "1000100100111100" => data_out <= rom_array(35132);
		when "1000100100111101" => data_out <= rom_array(35133);
		when "1000100100111110" => data_out <= rom_array(35134);
		when "1000100100111111" => data_out <= rom_array(35135);
		when "1000100101000000" => data_out <= rom_array(35136);
		when "1000100101000001" => data_out <= rom_array(35137);
		when "1000100101000010" => data_out <= rom_array(35138);
		when "1000100101000011" => data_out <= rom_array(35139);
		when "1000100101000100" => data_out <= rom_array(35140);
		when "1000100101000101" => data_out <= rom_array(35141);
		when "1000100101000110" => data_out <= rom_array(35142);
		when "1000100101000111" => data_out <= rom_array(35143);
		when "1000100101001000" => data_out <= rom_array(35144);
		when "1000100101001001" => data_out <= rom_array(35145);
		when "1000100101001010" => data_out <= rom_array(35146);
		when "1000100101001011" => data_out <= rom_array(35147);
		when "1000100101001100" => data_out <= rom_array(35148);
		when "1000100101001101" => data_out <= rom_array(35149);
		when "1000100101001110" => data_out <= rom_array(35150);
		when "1000100101001111" => data_out <= rom_array(35151);
		when "1000100101010000" => data_out <= rom_array(35152);
		when "1000100101010001" => data_out <= rom_array(35153);
		when "1000100101010010" => data_out <= rom_array(35154);
		when "1000100101010011" => data_out <= rom_array(35155);
		when "1000100101010100" => data_out <= rom_array(35156);
		when "1000100101010101" => data_out <= rom_array(35157);
		when "1000100101010110" => data_out <= rom_array(35158);
		when "1000100101010111" => data_out <= rom_array(35159);
		when "1000100101011000" => data_out <= rom_array(35160);
		when "1000100101011001" => data_out <= rom_array(35161);
		when "1000100101011010" => data_out <= rom_array(35162);
		when "1000100101011011" => data_out <= rom_array(35163);
		when "1000100101011100" => data_out <= rom_array(35164);
		when "1000100101011101" => data_out <= rom_array(35165);
		when "1000100101011110" => data_out <= rom_array(35166);
		when "1000100101011111" => data_out <= rom_array(35167);
		when "1000100101100000" => data_out <= rom_array(35168);
		when "1000100101100001" => data_out <= rom_array(35169);
		when "1000100101100010" => data_out <= rom_array(35170);
		when "1000100101100011" => data_out <= rom_array(35171);
		when "1000100101100100" => data_out <= rom_array(35172);
		when "1000100101100101" => data_out <= rom_array(35173);
		when "1000100101100110" => data_out <= rom_array(35174);
		when "1000100101100111" => data_out <= rom_array(35175);
		when "1000100101101000" => data_out <= rom_array(35176);
		when "1000100101101001" => data_out <= rom_array(35177);
		when "1000100101101010" => data_out <= rom_array(35178);
		when "1000100101101011" => data_out <= rom_array(35179);
		when "1000100101101100" => data_out <= rom_array(35180);
		when "1000100101101101" => data_out <= rom_array(35181);
		when "1000100101101110" => data_out <= rom_array(35182);
		when "1000100101101111" => data_out <= rom_array(35183);
		when "1000100101110000" => data_out <= rom_array(35184);
		when "1000100101110001" => data_out <= rom_array(35185);
		when "1000100101110010" => data_out <= rom_array(35186);
		when "1000100101110011" => data_out <= rom_array(35187);
		when "1000100101110100" => data_out <= rom_array(35188);
		when "1000100101110101" => data_out <= rom_array(35189);
		when "1000100101110110" => data_out <= rom_array(35190);
		when "1000100101110111" => data_out <= rom_array(35191);
		when "1000100101111000" => data_out <= rom_array(35192);
		when "1000100101111001" => data_out <= rom_array(35193);
		when "1000100101111010" => data_out <= rom_array(35194);
		when "1000100101111011" => data_out <= rom_array(35195);
		when "1000100101111100" => data_out <= rom_array(35196);
		when "1000100101111101" => data_out <= rom_array(35197);
		when "1000100101111110" => data_out <= rom_array(35198);
		when "1000100101111111" => data_out <= rom_array(35199);
		when "1000100110000000" => data_out <= rom_array(35200);
		when "1000100110000001" => data_out <= rom_array(35201);
		when "1000100110000010" => data_out <= rom_array(35202);
		when "1000100110000011" => data_out <= rom_array(35203);
		when "1000100110000100" => data_out <= rom_array(35204);
		when "1000100110000101" => data_out <= rom_array(35205);
		when "1000100110000110" => data_out <= rom_array(35206);
		when "1000100110000111" => data_out <= rom_array(35207);
		when "1000100110001000" => data_out <= rom_array(35208);
		when "1000100110001001" => data_out <= rom_array(35209);
		when "1000100110001010" => data_out <= rom_array(35210);
		when "1000100110001011" => data_out <= rom_array(35211);
		when "1000100110001100" => data_out <= rom_array(35212);
		when "1000100110001101" => data_out <= rom_array(35213);
		when "1000100110001110" => data_out <= rom_array(35214);
		when "1000100110001111" => data_out <= rom_array(35215);
		when "1000100110010000" => data_out <= rom_array(35216);
		when "1000100110010001" => data_out <= rom_array(35217);
		when "1000100110010010" => data_out <= rom_array(35218);
		when "1000100110010011" => data_out <= rom_array(35219);
		when "1000100110010100" => data_out <= rom_array(35220);
		when "1000100110010101" => data_out <= rom_array(35221);
		when "1000100110010110" => data_out <= rom_array(35222);
		when "1000100110010111" => data_out <= rom_array(35223);
		when "1000100110011000" => data_out <= rom_array(35224);
		when "1000100110011001" => data_out <= rom_array(35225);
		when "1000100110011010" => data_out <= rom_array(35226);
		when "1000100110011011" => data_out <= rom_array(35227);
		when "1000100110011100" => data_out <= rom_array(35228);
		when "1000100110011101" => data_out <= rom_array(35229);
		when "1000100110011110" => data_out <= rom_array(35230);
		when "1000100110011111" => data_out <= rom_array(35231);
		when "1000100110100000" => data_out <= rom_array(35232);
		when "1000100110100001" => data_out <= rom_array(35233);
		when "1000100110100010" => data_out <= rom_array(35234);
		when "1000100110100011" => data_out <= rom_array(35235);
		when "1000100110100100" => data_out <= rom_array(35236);
		when "1000100110100101" => data_out <= rom_array(35237);
		when "1000100110100110" => data_out <= rom_array(35238);
		when "1000100110100111" => data_out <= rom_array(35239);
		when "1000100110101000" => data_out <= rom_array(35240);
		when "1000100110101001" => data_out <= rom_array(35241);
		when "1000100110101010" => data_out <= rom_array(35242);
		when "1000100110101011" => data_out <= rom_array(35243);
		when "1000100110101100" => data_out <= rom_array(35244);
		when "1000100110101101" => data_out <= rom_array(35245);
		when "1000100110101110" => data_out <= rom_array(35246);
		when "1000100110101111" => data_out <= rom_array(35247);
		when "1000100110110000" => data_out <= rom_array(35248);
		when "1000100110110001" => data_out <= rom_array(35249);
		when "1000100110110010" => data_out <= rom_array(35250);
		when "1000100110110011" => data_out <= rom_array(35251);
		when "1000100110110100" => data_out <= rom_array(35252);
		when "1000100110110101" => data_out <= rom_array(35253);
		when "1000100110110110" => data_out <= rom_array(35254);
		when "1000100110110111" => data_out <= rom_array(35255);
		when "1000100110111000" => data_out <= rom_array(35256);
		when "1000100110111001" => data_out <= rom_array(35257);
		when "1000100110111010" => data_out <= rom_array(35258);
		when "1000100110111011" => data_out <= rom_array(35259);
		when "1000100110111100" => data_out <= rom_array(35260);
		when "1000100110111101" => data_out <= rom_array(35261);
		when "1000100110111110" => data_out <= rom_array(35262);
		when "1000100110111111" => data_out <= rom_array(35263);
		when "1000100111000000" => data_out <= rom_array(35264);
		when "1000100111000001" => data_out <= rom_array(35265);
		when "1000100111000010" => data_out <= rom_array(35266);
		when "1000100111000011" => data_out <= rom_array(35267);
		when "1000100111000100" => data_out <= rom_array(35268);
		when "1000100111000101" => data_out <= rom_array(35269);
		when "1000100111000110" => data_out <= rom_array(35270);
		when "1000100111000111" => data_out <= rom_array(35271);
		when "1000100111001000" => data_out <= rom_array(35272);
		when "1000100111001001" => data_out <= rom_array(35273);
		when "1000100111001010" => data_out <= rom_array(35274);
		when "1000100111001011" => data_out <= rom_array(35275);
		when "1000100111001100" => data_out <= rom_array(35276);
		when "1000100111001101" => data_out <= rom_array(35277);
		when "1000100111001110" => data_out <= rom_array(35278);
		when "1000100111001111" => data_out <= rom_array(35279);
		when "1000100111010000" => data_out <= rom_array(35280);
		when "1000100111010001" => data_out <= rom_array(35281);
		when "1000100111010010" => data_out <= rom_array(35282);
		when "1000100111010011" => data_out <= rom_array(35283);
		when "1000100111010100" => data_out <= rom_array(35284);
		when "1000100111010101" => data_out <= rom_array(35285);
		when "1000100111010110" => data_out <= rom_array(35286);
		when "1000100111010111" => data_out <= rom_array(35287);
		when "1000100111011000" => data_out <= rom_array(35288);
		when "1000100111011001" => data_out <= rom_array(35289);
		when "1000100111011010" => data_out <= rom_array(35290);
		when "1000100111011011" => data_out <= rom_array(35291);
		when "1000100111011100" => data_out <= rom_array(35292);
		when "1000100111011101" => data_out <= rom_array(35293);
		when "1000100111011110" => data_out <= rom_array(35294);
		when "1000100111011111" => data_out <= rom_array(35295);
		when "1000100111100000" => data_out <= rom_array(35296);
		when "1000100111100001" => data_out <= rom_array(35297);
		when "1000100111100010" => data_out <= rom_array(35298);
		when "1000100111100011" => data_out <= rom_array(35299);
		when "1000100111100100" => data_out <= rom_array(35300);
		when "1000100111100101" => data_out <= rom_array(35301);
		when "1000100111100110" => data_out <= rom_array(35302);
		when "1000100111100111" => data_out <= rom_array(35303);
		when "1000100111101000" => data_out <= rom_array(35304);
		when "1000100111101001" => data_out <= rom_array(35305);
		when "1000100111101010" => data_out <= rom_array(35306);
		when "1000100111101011" => data_out <= rom_array(35307);
		when "1000100111101100" => data_out <= rom_array(35308);
		when "1000100111101101" => data_out <= rom_array(35309);
		when "1000100111101110" => data_out <= rom_array(35310);
		when "1000100111101111" => data_out <= rom_array(35311);
		when "1000100111110000" => data_out <= rom_array(35312);
		when "1000100111110001" => data_out <= rom_array(35313);
		when "1000100111110010" => data_out <= rom_array(35314);
		when "1000100111110011" => data_out <= rom_array(35315);
		when "1000100111110100" => data_out <= rom_array(35316);
		when "1000100111110101" => data_out <= rom_array(35317);
		when "1000100111110110" => data_out <= rom_array(35318);
		when "1000100111110111" => data_out <= rom_array(35319);
		when "1000100111111000" => data_out <= rom_array(35320);
		when "1000100111111001" => data_out <= rom_array(35321);
		when "1000100111111010" => data_out <= rom_array(35322);
		when "1000100111111011" => data_out <= rom_array(35323);
		when "1000100111111100" => data_out <= rom_array(35324);
		when "1000100111111101" => data_out <= rom_array(35325);
		when "1000100111111110" => data_out <= rom_array(35326);
		when "1000100111111111" => data_out <= rom_array(35327);
		when "1000101000000000" => data_out <= rom_array(35328);
		when "1000101000000001" => data_out <= rom_array(35329);
		when "1000101000000010" => data_out <= rom_array(35330);
		when "1000101000000011" => data_out <= rom_array(35331);
		when "1000101000000100" => data_out <= rom_array(35332);
		when "1000101000000101" => data_out <= rom_array(35333);
		when "1000101000000110" => data_out <= rom_array(35334);
		when "1000101000000111" => data_out <= rom_array(35335);
		when "1000101000001000" => data_out <= rom_array(35336);
		when "1000101000001001" => data_out <= rom_array(35337);
		when "1000101000001010" => data_out <= rom_array(35338);
		when "1000101000001011" => data_out <= rom_array(35339);
		when "1000101000001100" => data_out <= rom_array(35340);
		when "1000101000001101" => data_out <= rom_array(35341);
		when "1000101000001110" => data_out <= rom_array(35342);
		when "1000101000001111" => data_out <= rom_array(35343);
		when "1000101000010000" => data_out <= rom_array(35344);
		when "1000101000010001" => data_out <= rom_array(35345);
		when "1000101000010010" => data_out <= rom_array(35346);
		when "1000101000010011" => data_out <= rom_array(35347);
		when "1000101000010100" => data_out <= rom_array(35348);
		when "1000101000010101" => data_out <= rom_array(35349);
		when "1000101000010110" => data_out <= rom_array(35350);
		when "1000101000010111" => data_out <= rom_array(35351);
		when "1000101000011000" => data_out <= rom_array(35352);
		when "1000101000011001" => data_out <= rom_array(35353);
		when "1000101000011010" => data_out <= rom_array(35354);
		when "1000101000011011" => data_out <= rom_array(35355);
		when "1000101000011100" => data_out <= rom_array(35356);
		when "1000101000011101" => data_out <= rom_array(35357);
		when "1000101000011110" => data_out <= rom_array(35358);
		when "1000101000011111" => data_out <= rom_array(35359);
		when "1000101000100000" => data_out <= rom_array(35360);
		when "1000101000100001" => data_out <= rom_array(35361);
		when "1000101000100010" => data_out <= rom_array(35362);
		when "1000101000100011" => data_out <= rom_array(35363);
		when "1000101000100100" => data_out <= rom_array(35364);
		when "1000101000100101" => data_out <= rom_array(35365);
		when "1000101000100110" => data_out <= rom_array(35366);
		when "1000101000100111" => data_out <= rom_array(35367);
		when "1000101000101000" => data_out <= rom_array(35368);
		when "1000101000101001" => data_out <= rom_array(35369);
		when "1000101000101010" => data_out <= rom_array(35370);
		when "1000101000101011" => data_out <= rom_array(35371);
		when "1000101000101100" => data_out <= rom_array(35372);
		when "1000101000101101" => data_out <= rom_array(35373);
		when "1000101000101110" => data_out <= rom_array(35374);
		when "1000101000101111" => data_out <= rom_array(35375);
		when "1000101000110000" => data_out <= rom_array(35376);
		when "1000101000110001" => data_out <= rom_array(35377);
		when "1000101000110010" => data_out <= rom_array(35378);
		when "1000101000110011" => data_out <= rom_array(35379);
		when "1000101000110100" => data_out <= rom_array(35380);
		when "1000101000110101" => data_out <= rom_array(35381);
		when "1000101000110110" => data_out <= rom_array(35382);
		when "1000101000110111" => data_out <= rom_array(35383);
		when "1000101000111000" => data_out <= rom_array(35384);
		when "1000101000111001" => data_out <= rom_array(35385);
		when "1000101000111010" => data_out <= rom_array(35386);
		when "1000101000111011" => data_out <= rom_array(35387);
		when "1000101000111100" => data_out <= rom_array(35388);
		when "1000101000111101" => data_out <= rom_array(35389);
		when "1000101000111110" => data_out <= rom_array(35390);
		when "1000101000111111" => data_out <= rom_array(35391);
		when "1000101001000000" => data_out <= rom_array(35392);
		when "1000101001000001" => data_out <= rom_array(35393);
		when "1000101001000010" => data_out <= rom_array(35394);
		when "1000101001000011" => data_out <= rom_array(35395);
		when "1000101001000100" => data_out <= rom_array(35396);
		when "1000101001000101" => data_out <= rom_array(35397);
		when "1000101001000110" => data_out <= rom_array(35398);
		when "1000101001000111" => data_out <= rom_array(35399);
		when "1000101001001000" => data_out <= rom_array(35400);
		when "1000101001001001" => data_out <= rom_array(35401);
		when "1000101001001010" => data_out <= rom_array(35402);
		when "1000101001001011" => data_out <= rom_array(35403);
		when "1000101001001100" => data_out <= rom_array(35404);
		when "1000101001001101" => data_out <= rom_array(35405);
		when "1000101001001110" => data_out <= rom_array(35406);
		when "1000101001001111" => data_out <= rom_array(35407);
		when "1000101001010000" => data_out <= rom_array(35408);
		when "1000101001010001" => data_out <= rom_array(35409);
		when "1000101001010010" => data_out <= rom_array(35410);
		when "1000101001010011" => data_out <= rom_array(35411);
		when "1000101001010100" => data_out <= rom_array(35412);
		when "1000101001010101" => data_out <= rom_array(35413);
		when "1000101001010110" => data_out <= rom_array(35414);
		when "1000101001010111" => data_out <= rom_array(35415);
		when "1000101001011000" => data_out <= rom_array(35416);
		when "1000101001011001" => data_out <= rom_array(35417);
		when "1000101001011010" => data_out <= rom_array(35418);
		when "1000101001011011" => data_out <= rom_array(35419);
		when "1000101001011100" => data_out <= rom_array(35420);
		when "1000101001011101" => data_out <= rom_array(35421);
		when "1000101001011110" => data_out <= rom_array(35422);
		when "1000101001011111" => data_out <= rom_array(35423);
		when "1000101001100000" => data_out <= rom_array(35424);
		when "1000101001100001" => data_out <= rom_array(35425);
		when "1000101001100010" => data_out <= rom_array(35426);
		when "1000101001100011" => data_out <= rom_array(35427);
		when "1000101001100100" => data_out <= rom_array(35428);
		when "1000101001100101" => data_out <= rom_array(35429);
		when "1000101001100110" => data_out <= rom_array(35430);
		when "1000101001100111" => data_out <= rom_array(35431);
		when "1000101001101000" => data_out <= rom_array(35432);
		when "1000101001101001" => data_out <= rom_array(35433);
		when "1000101001101010" => data_out <= rom_array(35434);
		when "1000101001101011" => data_out <= rom_array(35435);
		when "1000101001101100" => data_out <= rom_array(35436);
		when "1000101001101101" => data_out <= rom_array(35437);
		when "1000101001101110" => data_out <= rom_array(35438);
		when "1000101001101111" => data_out <= rom_array(35439);
		when "1000101001110000" => data_out <= rom_array(35440);
		when "1000101001110001" => data_out <= rom_array(35441);
		when "1000101001110010" => data_out <= rom_array(35442);
		when "1000101001110011" => data_out <= rom_array(35443);
		when "1000101001110100" => data_out <= rom_array(35444);
		when "1000101001110101" => data_out <= rom_array(35445);
		when "1000101001110110" => data_out <= rom_array(35446);
		when "1000101001110111" => data_out <= rom_array(35447);
		when "1000101001111000" => data_out <= rom_array(35448);
		when "1000101001111001" => data_out <= rom_array(35449);
		when "1000101001111010" => data_out <= rom_array(35450);
		when "1000101001111011" => data_out <= rom_array(35451);
		when "1000101001111100" => data_out <= rom_array(35452);
		when "1000101001111101" => data_out <= rom_array(35453);
		when "1000101001111110" => data_out <= rom_array(35454);
		when "1000101001111111" => data_out <= rom_array(35455);
		when "1000101010000000" => data_out <= rom_array(35456);
		when "1000101010000001" => data_out <= rom_array(35457);
		when "1000101010000010" => data_out <= rom_array(35458);
		when "1000101010000011" => data_out <= rom_array(35459);
		when "1000101010000100" => data_out <= rom_array(35460);
		when "1000101010000101" => data_out <= rom_array(35461);
		when "1000101010000110" => data_out <= rom_array(35462);
		when "1000101010000111" => data_out <= rom_array(35463);
		when "1000101010001000" => data_out <= rom_array(35464);
		when "1000101010001001" => data_out <= rom_array(35465);
		when "1000101010001010" => data_out <= rom_array(35466);
		when "1000101010001011" => data_out <= rom_array(35467);
		when "1000101010001100" => data_out <= rom_array(35468);
		when "1000101010001101" => data_out <= rom_array(35469);
		when "1000101010001110" => data_out <= rom_array(35470);
		when "1000101010001111" => data_out <= rom_array(35471);
		when "1000101010010000" => data_out <= rom_array(35472);
		when "1000101010010001" => data_out <= rom_array(35473);
		when "1000101010010010" => data_out <= rom_array(35474);
		when "1000101010010011" => data_out <= rom_array(35475);
		when "1000101010010100" => data_out <= rom_array(35476);
		when "1000101010010101" => data_out <= rom_array(35477);
		when "1000101010010110" => data_out <= rom_array(35478);
		when "1000101010010111" => data_out <= rom_array(35479);
		when "1000101010011000" => data_out <= rom_array(35480);
		when "1000101010011001" => data_out <= rom_array(35481);
		when "1000101010011010" => data_out <= rom_array(35482);
		when "1000101010011011" => data_out <= rom_array(35483);
		when "1000101010011100" => data_out <= rom_array(35484);
		when "1000101010011101" => data_out <= rom_array(35485);
		when "1000101010011110" => data_out <= rom_array(35486);
		when "1000101010011111" => data_out <= rom_array(35487);
		when "1000101010100000" => data_out <= rom_array(35488);
		when "1000101010100001" => data_out <= rom_array(35489);
		when "1000101010100010" => data_out <= rom_array(35490);
		when "1000101010100011" => data_out <= rom_array(35491);
		when "1000101010100100" => data_out <= rom_array(35492);
		when "1000101010100101" => data_out <= rom_array(35493);
		when "1000101010100110" => data_out <= rom_array(35494);
		when "1000101010100111" => data_out <= rom_array(35495);
		when "1000101010101000" => data_out <= rom_array(35496);
		when "1000101010101001" => data_out <= rom_array(35497);
		when "1000101010101010" => data_out <= rom_array(35498);
		when "1000101010101011" => data_out <= rom_array(35499);
		when "1000101010101100" => data_out <= rom_array(35500);
		when "1000101010101101" => data_out <= rom_array(35501);
		when "1000101010101110" => data_out <= rom_array(35502);
		when "1000101010101111" => data_out <= rom_array(35503);
		when "1000101010110000" => data_out <= rom_array(35504);
		when "1000101010110001" => data_out <= rom_array(35505);
		when "1000101010110010" => data_out <= rom_array(35506);
		when "1000101010110011" => data_out <= rom_array(35507);
		when "1000101010110100" => data_out <= rom_array(35508);
		when "1000101010110101" => data_out <= rom_array(35509);
		when "1000101010110110" => data_out <= rom_array(35510);
		when "1000101010110111" => data_out <= rom_array(35511);
		when "1000101010111000" => data_out <= rom_array(35512);
		when "1000101010111001" => data_out <= rom_array(35513);
		when "1000101010111010" => data_out <= rom_array(35514);
		when "1000101010111011" => data_out <= rom_array(35515);
		when "1000101010111100" => data_out <= rom_array(35516);
		when "1000101010111101" => data_out <= rom_array(35517);
		when "1000101010111110" => data_out <= rom_array(35518);
		when "1000101010111111" => data_out <= rom_array(35519);
		when "1000101011000000" => data_out <= rom_array(35520);
		when "1000101011000001" => data_out <= rom_array(35521);
		when "1000101011000010" => data_out <= rom_array(35522);
		when "1000101011000011" => data_out <= rom_array(35523);
		when "1000101011000100" => data_out <= rom_array(35524);
		when "1000101011000101" => data_out <= rom_array(35525);
		when "1000101011000110" => data_out <= rom_array(35526);
		when "1000101011000111" => data_out <= rom_array(35527);
		when "1000101011001000" => data_out <= rom_array(35528);
		when "1000101011001001" => data_out <= rom_array(35529);
		when "1000101011001010" => data_out <= rom_array(35530);
		when "1000101011001011" => data_out <= rom_array(35531);
		when "1000101011001100" => data_out <= rom_array(35532);
		when "1000101011001101" => data_out <= rom_array(35533);
		when "1000101011001110" => data_out <= rom_array(35534);
		when "1000101011001111" => data_out <= rom_array(35535);
		when "1000101011010000" => data_out <= rom_array(35536);
		when "1000101011010001" => data_out <= rom_array(35537);
		when "1000101011010010" => data_out <= rom_array(35538);
		when "1000101011010011" => data_out <= rom_array(35539);
		when "1000101011010100" => data_out <= rom_array(35540);
		when "1000101011010101" => data_out <= rom_array(35541);
		when "1000101011010110" => data_out <= rom_array(35542);
		when "1000101011010111" => data_out <= rom_array(35543);
		when "1000101011011000" => data_out <= rom_array(35544);
		when "1000101011011001" => data_out <= rom_array(35545);
		when "1000101011011010" => data_out <= rom_array(35546);
		when "1000101011011011" => data_out <= rom_array(35547);
		when "1000101011011100" => data_out <= rom_array(35548);
		when "1000101011011101" => data_out <= rom_array(35549);
		when "1000101011011110" => data_out <= rom_array(35550);
		when "1000101011011111" => data_out <= rom_array(35551);
		when "1000101011100000" => data_out <= rom_array(35552);
		when "1000101011100001" => data_out <= rom_array(35553);
		when "1000101011100010" => data_out <= rom_array(35554);
		when "1000101011100011" => data_out <= rom_array(35555);
		when "1000101011100100" => data_out <= rom_array(35556);
		when "1000101011100101" => data_out <= rom_array(35557);
		when "1000101011100110" => data_out <= rom_array(35558);
		when "1000101011100111" => data_out <= rom_array(35559);
		when "1000101011101000" => data_out <= rom_array(35560);
		when "1000101011101001" => data_out <= rom_array(35561);
		when "1000101011101010" => data_out <= rom_array(35562);
		when "1000101011101011" => data_out <= rom_array(35563);
		when "1000101011101100" => data_out <= rom_array(35564);
		when "1000101011101101" => data_out <= rom_array(35565);
		when "1000101011101110" => data_out <= rom_array(35566);
		when "1000101011101111" => data_out <= rom_array(35567);
		when "1000101011110000" => data_out <= rom_array(35568);
		when "1000101011110001" => data_out <= rom_array(35569);
		when "1000101011110010" => data_out <= rom_array(35570);
		when "1000101011110011" => data_out <= rom_array(35571);
		when "1000101011110100" => data_out <= rom_array(35572);
		when "1000101011110101" => data_out <= rom_array(35573);
		when "1000101011110110" => data_out <= rom_array(35574);
		when "1000101011110111" => data_out <= rom_array(35575);
		when "1000101011111000" => data_out <= rom_array(35576);
		when "1000101011111001" => data_out <= rom_array(35577);
		when "1000101011111010" => data_out <= rom_array(35578);
		when "1000101011111011" => data_out <= rom_array(35579);
		when "1000101011111100" => data_out <= rom_array(35580);
		when "1000101011111101" => data_out <= rom_array(35581);
		when "1000101011111110" => data_out <= rom_array(35582);
		when "1000101011111111" => data_out <= rom_array(35583);
		when "1000101100000000" => data_out <= rom_array(35584);
		when "1000101100000001" => data_out <= rom_array(35585);
		when "1000101100000010" => data_out <= rom_array(35586);
		when "1000101100000011" => data_out <= rom_array(35587);
		when "1000101100000100" => data_out <= rom_array(35588);
		when "1000101100000101" => data_out <= rom_array(35589);
		when "1000101100000110" => data_out <= rom_array(35590);
		when "1000101100000111" => data_out <= rom_array(35591);
		when "1000101100001000" => data_out <= rom_array(35592);
		when "1000101100001001" => data_out <= rom_array(35593);
		when "1000101100001010" => data_out <= rom_array(35594);
		when "1000101100001011" => data_out <= rom_array(35595);
		when "1000101100001100" => data_out <= rom_array(35596);
		when "1000101100001101" => data_out <= rom_array(35597);
		when "1000101100001110" => data_out <= rom_array(35598);
		when "1000101100001111" => data_out <= rom_array(35599);
		when "1000101100010000" => data_out <= rom_array(35600);
		when "1000101100010001" => data_out <= rom_array(35601);
		when "1000101100010010" => data_out <= rom_array(35602);
		when "1000101100010011" => data_out <= rom_array(35603);
		when "1000101100010100" => data_out <= rom_array(35604);
		when "1000101100010101" => data_out <= rom_array(35605);
		when "1000101100010110" => data_out <= rom_array(35606);
		when "1000101100010111" => data_out <= rom_array(35607);
		when "1000101100011000" => data_out <= rom_array(35608);
		when "1000101100011001" => data_out <= rom_array(35609);
		when "1000101100011010" => data_out <= rom_array(35610);
		when "1000101100011011" => data_out <= rom_array(35611);
		when "1000101100011100" => data_out <= rom_array(35612);
		when "1000101100011101" => data_out <= rom_array(35613);
		when "1000101100011110" => data_out <= rom_array(35614);
		when "1000101100011111" => data_out <= rom_array(35615);
		when "1000101100100000" => data_out <= rom_array(35616);
		when "1000101100100001" => data_out <= rom_array(35617);
		when "1000101100100010" => data_out <= rom_array(35618);
		when "1000101100100011" => data_out <= rom_array(35619);
		when "1000101100100100" => data_out <= rom_array(35620);
		when "1000101100100101" => data_out <= rom_array(35621);
		when "1000101100100110" => data_out <= rom_array(35622);
		when "1000101100100111" => data_out <= rom_array(35623);
		when "1000101100101000" => data_out <= rom_array(35624);
		when "1000101100101001" => data_out <= rom_array(35625);
		when "1000101100101010" => data_out <= rom_array(35626);
		when "1000101100101011" => data_out <= rom_array(35627);
		when "1000101100101100" => data_out <= rom_array(35628);
		when "1000101100101101" => data_out <= rom_array(35629);
		when "1000101100101110" => data_out <= rom_array(35630);
		when "1000101100101111" => data_out <= rom_array(35631);
		when "1000101100110000" => data_out <= rom_array(35632);
		when "1000101100110001" => data_out <= rom_array(35633);
		when "1000101100110010" => data_out <= rom_array(35634);
		when "1000101100110011" => data_out <= rom_array(35635);
		when "1000101100110100" => data_out <= rom_array(35636);
		when "1000101100110101" => data_out <= rom_array(35637);
		when "1000101100110110" => data_out <= rom_array(35638);
		when "1000101100110111" => data_out <= rom_array(35639);
		when "1000101100111000" => data_out <= rom_array(35640);
		when "1000101100111001" => data_out <= rom_array(35641);
		when "1000101100111010" => data_out <= rom_array(35642);
		when "1000101100111011" => data_out <= rom_array(35643);
		when "1000101100111100" => data_out <= rom_array(35644);
		when "1000101100111101" => data_out <= rom_array(35645);
		when "1000101100111110" => data_out <= rom_array(35646);
		when "1000101100111111" => data_out <= rom_array(35647);
		when "1000101101000000" => data_out <= rom_array(35648);
		when "1000101101000001" => data_out <= rom_array(35649);
		when "1000101101000010" => data_out <= rom_array(35650);
		when "1000101101000011" => data_out <= rom_array(35651);
		when "1000101101000100" => data_out <= rom_array(35652);
		when "1000101101000101" => data_out <= rom_array(35653);
		when "1000101101000110" => data_out <= rom_array(35654);
		when "1000101101000111" => data_out <= rom_array(35655);
		when "1000101101001000" => data_out <= rom_array(35656);
		when "1000101101001001" => data_out <= rom_array(35657);
		when "1000101101001010" => data_out <= rom_array(35658);
		when "1000101101001011" => data_out <= rom_array(35659);
		when "1000101101001100" => data_out <= rom_array(35660);
		when "1000101101001101" => data_out <= rom_array(35661);
		when "1000101101001110" => data_out <= rom_array(35662);
		when "1000101101001111" => data_out <= rom_array(35663);
		when "1000101101010000" => data_out <= rom_array(35664);
		when "1000101101010001" => data_out <= rom_array(35665);
		when "1000101101010010" => data_out <= rom_array(35666);
		when "1000101101010011" => data_out <= rom_array(35667);
		when "1000101101010100" => data_out <= rom_array(35668);
		when "1000101101010101" => data_out <= rom_array(35669);
		when "1000101101010110" => data_out <= rom_array(35670);
		when "1000101101010111" => data_out <= rom_array(35671);
		when "1000101101011000" => data_out <= rom_array(35672);
		when "1000101101011001" => data_out <= rom_array(35673);
		when "1000101101011010" => data_out <= rom_array(35674);
		when "1000101101011011" => data_out <= rom_array(35675);
		when "1000101101011100" => data_out <= rom_array(35676);
		when "1000101101011101" => data_out <= rom_array(35677);
		when "1000101101011110" => data_out <= rom_array(35678);
		when "1000101101011111" => data_out <= rom_array(35679);
		when "1000101101100000" => data_out <= rom_array(35680);
		when "1000101101100001" => data_out <= rom_array(35681);
		when "1000101101100010" => data_out <= rom_array(35682);
		when "1000101101100011" => data_out <= rom_array(35683);
		when "1000101101100100" => data_out <= rom_array(35684);
		when "1000101101100101" => data_out <= rom_array(35685);
		when "1000101101100110" => data_out <= rom_array(35686);
		when "1000101101100111" => data_out <= rom_array(35687);
		when "1000101101101000" => data_out <= rom_array(35688);
		when "1000101101101001" => data_out <= rom_array(35689);
		when "1000101101101010" => data_out <= rom_array(35690);
		when "1000101101101011" => data_out <= rom_array(35691);
		when "1000101101101100" => data_out <= rom_array(35692);
		when "1000101101101101" => data_out <= rom_array(35693);
		when "1000101101101110" => data_out <= rom_array(35694);
		when "1000101101101111" => data_out <= rom_array(35695);
		when "1000101101110000" => data_out <= rom_array(35696);
		when "1000101101110001" => data_out <= rom_array(35697);
		when "1000101101110010" => data_out <= rom_array(35698);
		when "1000101101110011" => data_out <= rom_array(35699);
		when "1000101101110100" => data_out <= rom_array(35700);
		when "1000101101110101" => data_out <= rom_array(35701);
		when "1000101101110110" => data_out <= rom_array(35702);
		when "1000101101110111" => data_out <= rom_array(35703);
		when "1000101101111000" => data_out <= rom_array(35704);
		when "1000101101111001" => data_out <= rom_array(35705);
		when "1000101101111010" => data_out <= rom_array(35706);
		when "1000101101111011" => data_out <= rom_array(35707);
		when "1000101101111100" => data_out <= rom_array(35708);
		when "1000101101111101" => data_out <= rom_array(35709);
		when "1000101101111110" => data_out <= rom_array(35710);
		when "1000101101111111" => data_out <= rom_array(35711);
		when "1000101110000000" => data_out <= rom_array(35712);
		when "1000101110000001" => data_out <= rom_array(35713);
		when "1000101110000010" => data_out <= rom_array(35714);
		when "1000101110000011" => data_out <= rom_array(35715);
		when "1000101110000100" => data_out <= rom_array(35716);
		when "1000101110000101" => data_out <= rom_array(35717);
		when "1000101110000110" => data_out <= rom_array(35718);
		when "1000101110000111" => data_out <= rom_array(35719);
		when "1000101110001000" => data_out <= rom_array(35720);
		when "1000101110001001" => data_out <= rom_array(35721);
		when "1000101110001010" => data_out <= rom_array(35722);
		when "1000101110001011" => data_out <= rom_array(35723);
		when "1000101110001100" => data_out <= rom_array(35724);
		when "1000101110001101" => data_out <= rom_array(35725);
		when "1000101110001110" => data_out <= rom_array(35726);
		when "1000101110001111" => data_out <= rom_array(35727);
		when "1000101110010000" => data_out <= rom_array(35728);
		when "1000101110010001" => data_out <= rom_array(35729);
		when "1000101110010010" => data_out <= rom_array(35730);
		when "1000101110010011" => data_out <= rom_array(35731);
		when "1000101110010100" => data_out <= rom_array(35732);
		when "1000101110010101" => data_out <= rom_array(35733);
		when "1000101110010110" => data_out <= rom_array(35734);
		when "1000101110010111" => data_out <= rom_array(35735);
		when "1000101110011000" => data_out <= rom_array(35736);
		when "1000101110011001" => data_out <= rom_array(35737);
		when "1000101110011010" => data_out <= rom_array(35738);
		when "1000101110011011" => data_out <= rom_array(35739);
		when "1000101110011100" => data_out <= rom_array(35740);
		when "1000101110011101" => data_out <= rom_array(35741);
		when "1000101110011110" => data_out <= rom_array(35742);
		when "1000101110011111" => data_out <= rom_array(35743);
		when "1000101110100000" => data_out <= rom_array(35744);
		when "1000101110100001" => data_out <= rom_array(35745);
		when "1000101110100010" => data_out <= rom_array(35746);
		when "1000101110100011" => data_out <= rom_array(35747);
		when "1000101110100100" => data_out <= rom_array(35748);
		when "1000101110100101" => data_out <= rom_array(35749);
		when "1000101110100110" => data_out <= rom_array(35750);
		when "1000101110100111" => data_out <= rom_array(35751);
		when "1000101110101000" => data_out <= rom_array(35752);
		when "1000101110101001" => data_out <= rom_array(35753);
		when "1000101110101010" => data_out <= rom_array(35754);
		when "1000101110101011" => data_out <= rom_array(35755);
		when "1000101110101100" => data_out <= rom_array(35756);
		when "1000101110101101" => data_out <= rom_array(35757);
		when "1000101110101110" => data_out <= rom_array(35758);
		when "1000101110101111" => data_out <= rom_array(35759);
		when "1000101110110000" => data_out <= rom_array(35760);
		when "1000101110110001" => data_out <= rom_array(35761);
		when "1000101110110010" => data_out <= rom_array(35762);
		when "1000101110110011" => data_out <= rom_array(35763);
		when "1000101110110100" => data_out <= rom_array(35764);
		when "1000101110110101" => data_out <= rom_array(35765);
		when "1000101110110110" => data_out <= rom_array(35766);
		when "1000101110110111" => data_out <= rom_array(35767);
		when "1000101110111000" => data_out <= rom_array(35768);
		when "1000101110111001" => data_out <= rom_array(35769);
		when "1000101110111010" => data_out <= rom_array(35770);
		when "1000101110111011" => data_out <= rom_array(35771);
		when "1000101110111100" => data_out <= rom_array(35772);
		when "1000101110111101" => data_out <= rom_array(35773);
		when "1000101110111110" => data_out <= rom_array(35774);
		when "1000101110111111" => data_out <= rom_array(35775);
		when "1000101111000000" => data_out <= rom_array(35776);
		when "1000101111000001" => data_out <= rom_array(35777);
		when "1000101111000010" => data_out <= rom_array(35778);
		when "1000101111000011" => data_out <= rom_array(35779);
		when "1000101111000100" => data_out <= rom_array(35780);
		when "1000101111000101" => data_out <= rom_array(35781);
		when "1000101111000110" => data_out <= rom_array(35782);
		when "1000101111000111" => data_out <= rom_array(35783);
		when "1000101111001000" => data_out <= rom_array(35784);
		when "1000101111001001" => data_out <= rom_array(35785);
		when "1000101111001010" => data_out <= rom_array(35786);
		when "1000101111001011" => data_out <= rom_array(35787);
		when "1000101111001100" => data_out <= rom_array(35788);
		when "1000101111001101" => data_out <= rom_array(35789);
		when "1000101111001110" => data_out <= rom_array(35790);
		when "1000101111001111" => data_out <= rom_array(35791);
		when "1000101111010000" => data_out <= rom_array(35792);
		when "1000101111010001" => data_out <= rom_array(35793);
		when "1000101111010010" => data_out <= rom_array(35794);
		when "1000101111010011" => data_out <= rom_array(35795);
		when "1000101111010100" => data_out <= rom_array(35796);
		when "1000101111010101" => data_out <= rom_array(35797);
		when "1000101111010110" => data_out <= rom_array(35798);
		when "1000101111010111" => data_out <= rom_array(35799);
		when "1000101111011000" => data_out <= rom_array(35800);
		when "1000101111011001" => data_out <= rom_array(35801);
		when "1000101111011010" => data_out <= rom_array(35802);
		when "1000101111011011" => data_out <= rom_array(35803);
		when "1000101111011100" => data_out <= rom_array(35804);
		when "1000101111011101" => data_out <= rom_array(35805);
		when "1000101111011110" => data_out <= rom_array(35806);
		when "1000101111011111" => data_out <= rom_array(35807);
		when "1000101111100000" => data_out <= rom_array(35808);
		when "1000101111100001" => data_out <= rom_array(35809);
		when "1000101111100010" => data_out <= rom_array(35810);
		when "1000101111100011" => data_out <= rom_array(35811);
		when "1000101111100100" => data_out <= rom_array(35812);
		when "1000101111100101" => data_out <= rom_array(35813);
		when "1000101111100110" => data_out <= rom_array(35814);
		when "1000101111100111" => data_out <= rom_array(35815);
		when "1000101111101000" => data_out <= rom_array(35816);
		when "1000101111101001" => data_out <= rom_array(35817);
		when "1000101111101010" => data_out <= rom_array(35818);
		when "1000101111101011" => data_out <= rom_array(35819);
		when "1000101111101100" => data_out <= rom_array(35820);
		when "1000101111101101" => data_out <= rom_array(35821);
		when "1000101111101110" => data_out <= rom_array(35822);
		when "1000101111101111" => data_out <= rom_array(35823);
		when "1000101111110000" => data_out <= rom_array(35824);
		when "1000101111110001" => data_out <= rom_array(35825);
		when "1000101111110010" => data_out <= rom_array(35826);
		when "1000101111110011" => data_out <= rom_array(35827);
		when "1000101111110100" => data_out <= rom_array(35828);
		when "1000101111110101" => data_out <= rom_array(35829);
		when "1000101111110110" => data_out <= rom_array(35830);
		when "1000101111110111" => data_out <= rom_array(35831);
		when "1000101111111000" => data_out <= rom_array(35832);
		when "1000101111111001" => data_out <= rom_array(35833);
		when "1000101111111010" => data_out <= rom_array(35834);
		when "1000101111111011" => data_out <= rom_array(35835);
		when "1000101111111100" => data_out <= rom_array(35836);
		when "1000101111111101" => data_out <= rom_array(35837);
		when "1000101111111110" => data_out <= rom_array(35838);
		when "1000101111111111" => data_out <= rom_array(35839);
		when "1000110000000000" => data_out <= rom_array(35840);
		when "1000110000000001" => data_out <= rom_array(35841);
		when "1000110000000010" => data_out <= rom_array(35842);
		when "1000110000000011" => data_out <= rom_array(35843);
		when "1000110000000100" => data_out <= rom_array(35844);
		when "1000110000000101" => data_out <= rom_array(35845);
		when "1000110000000110" => data_out <= rom_array(35846);
		when "1000110000000111" => data_out <= rom_array(35847);
		when "1000110000001000" => data_out <= rom_array(35848);
		when "1000110000001001" => data_out <= rom_array(35849);
		when "1000110000001010" => data_out <= rom_array(35850);
		when "1000110000001011" => data_out <= rom_array(35851);
		when "1000110000001100" => data_out <= rom_array(35852);
		when "1000110000001101" => data_out <= rom_array(35853);
		when "1000110000001110" => data_out <= rom_array(35854);
		when "1000110000001111" => data_out <= rom_array(35855);
		when "1000110000010000" => data_out <= rom_array(35856);
		when "1000110000010001" => data_out <= rom_array(35857);
		when "1000110000010010" => data_out <= rom_array(35858);
		when "1000110000010011" => data_out <= rom_array(35859);
		when "1000110000010100" => data_out <= rom_array(35860);
		when "1000110000010101" => data_out <= rom_array(35861);
		when "1000110000010110" => data_out <= rom_array(35862);
		when "1000110000010111" => data_out <= rom_array(35863);
		when "1000110000011000" => data_out <= rom_array(35864);
		when "1000110000011001" => data_out <= rom_array(35865);
		when "1000110000011010" => data_out <= rom_array(35866);
		when "1000110000011011" => data_out <= rom_array(35867);
		when "1000110000011100" => data_out <= rom_array(35868);
		when "1000110000011101" => data_out <= rom_array(35869);
		when "1000110000011110" => data_out <= rom_array(35870);
		when "1000110000011111" => data_out <= rom_array(35871);
		when "1000110000100000" => data_out <= rom_array(35872);
		when "1000110000100001" => data_out <= rom_array(35873);
		when "1000110000100010" => data_out <= rom_array(35874);
		when "1000110000100011" => data_out <= rom_array(35875);
		when "1000110000100100" => data_out <= rom_array(35876);
		when "1000110000100101" => data_out <= rom_array(35877);
		when "1000110000100110" => data_out <= rom_array(35878);
		when "1000110000100111" => data_out <= rom_array(35879);
		when "1000110000101000" => data_out <= rom_array(35880);
		when "1000110000101001" => data_out <= rom_array(35881);
		when "1000110000101010" => data_out <= rom_array(35882);
		when "1000110000101011" => data_out <= rom_array(35883);
		when "1000110000101100" => data_out <= rom_array(35884);
		when "1000110000101101" => data_out <= rom_array(35885);
		when "1000110000101110" => data_out <= rom_array(35886);
		when "1000110000101111" => data_out <= rom_array(35887);
		when "1000110000110000" => data_out <= rom_array(35888);
		when "1000110000110001" => data_out <= rom_array(35889);
		when "1000110000110010" => data_out <= rom_array(35890);
		when "1000110000110011" => data_out <= rom_array(35891);
		when "1000110000110100" => data_out <= rom_array(35892);
		when "1000110000110101" => data_out <= rom_array(35893);
		when "1000110000110110" => data_out <= rom_array(35894);
		when "1000110000110111" => data_out <= rom_array(35895);
		when "1000110000111000" => data_out <= rom_array(35896);
		when "1000110000111001" => data_out <= rom_array(35897);
		when "1000110000111010" => data_out <= rom_array(35898);
		when "1000110000111011" => data_out <= rom_array(35899);
		when "1000110000111100" => data_out <= rom_array(35900);
		when "1000110000111101" => data_out <= rom_array(35901);
		when "1000110000111110" => data_out <= rom_array(35902);
		when "1000110000111111" => data_out <= rom_array(35903);
		when "1000110001000000" => data_out <= rom_array(35904);
		when "1000110001000001" => data_out <= rom_array(35905);
		when "1000110001000010" => data_out <= rom_array(35906);
		when "1000110001000011" => data_out <= rom_array(35907);
		when "1000110001000100" => data_out <= rom_array(35908);
		when "1000110001000101" => data_out <= rom_array(35909);
		when "1000110001000110" => data_out <= rom_array(35910);
		when "1000110001000111" => data_out <= rom_array(35911);
		when "1000110001001000" => data_out <= rom_array(35912);
		when "1000110001001001" => data_out <= rom_array(35913);
		when "1000110001001010" => data_out <= rom_array(35914);
		when "1000110001001011" => data_out <= rom_array(35915);
		when "1000110001001100" => data_out <= rom_array(35916);
		when "1000110001001101" => data_out <= rom_array(35917);
		when "1000110001001110" => data_out <= rom_array(35918);
		when "1000110001001111" => data_out <= rom_array(35919);
		when "1000110001010000" => data_out <= rom_array(35920);
		when "1000110001010001" => data_out <= rom_array(35921);
		when "1000110001010010" => data_out <= rom_array(35922);
		when "1000110001010011" => data_out <= rom_array(35923);
		when "1000110001010100" => data_out <= rom_array(35924);
		when "1000110001010101" => data_out <= rom_array(35925);
		when "1000110001010110" => data_out <= rom_array(35926);
		when "1000110001010111" => data_out <= rom_array(35927);
		when "1000110001011000" => data_out <= rom_array(35928);
		when "1000110001011001" => data_out <= rom_array(35929);
		when "1000110001011010" => data_out <= rom_array(35930);
		when "1000110001011011" => data_out <= rom_array(35931);
		when "1000110001011100" => data_out <= rom_array(35932);
		when "1000110001011101" => data_out <= rom_array(35933);
		when "1000110001011110" => data_out <= rom_array(35934);
		when "1000110001011111" => data_out <= rom_array(35935);
		when "1000110001100000" => data_out <= rom_array(35936);
		when "1000110001100001" => data_out <= rom_array(35937);
		when "1000110001100010" => data_out <= rom_array(35938);
		when "1000110001100011" => data_out <= rom_array(35939);
		when "1000110001100100" => data_out <= rom_array(35940);
		when "1000110001100101" => data_out <= rom_array(35941);
		when "1000110001100110" => data_out <= rom_array(35942);
		when "1000110001100111" => data_out <= rom_array(35943);
		when "1000110001101000" => data_out <= rom_array(35944);
		when "1000110001101001" => data_out <= rom_array(35945);
		when "1000110001101010" => data_out <= rom_array(35946);
		when "1000110001101011" => data_out <= rom_array(35947);
		when "1000110001101100" => data_out <= rom_array(35948);
		when "1000110001101101" => data_out <= rom_array(35949);
		when "1000110001101110" => data_out <= rom_array(35950);
		when "1000110001101111" => data_out <= rom_array(35951);
		when "1000110001110000" => data_out <= rom_array(35952);
		when "1000110001110001" => data_out <= rom_array(35953);
		when "1000110001110010" => data_out <= rom_array(35954);
		when "1000110001110011" => data_out <= rom_array(35955);
		when "1000110001110100" => data_out <= rom_array(35956);
		when "1000110001110101" => data_out <= rom_array(35957);
		when "1000110001110110" => data_out <= rom_array(35958);
		when "1000110001110111" => data_out <= rom_array(35959);
		when "1000110001111000" => data_out <= rom_array(35960);
		when "1000110001111001" => data_out <= rom_array(35961);
		when "1000110001111010" => data_out <= rom_array(35962);
		when "1000110001111011" => data_out <= rom_array(35963);
		when "1000110001111100" => data_out <= rom_array(35964);
		when "1000110001111101" => data_out <= rom_array(35965);
		when "1000110001111110" => data_out <= rom_array(35966);
		when "1000110001111111" => data_out <= rom_array(35967);
		when "1000110010000000" => data_out <= rom_array(35968);
		when "1000110010000001" => data_out <= rom_array(35969);
		when "1000110010000010" => data_out <= rom_array(35970);
		when "1000110010000011" => data_out <= rom_array(35971);
		when "1000110010000100" => data_out <= rom_array(35972);
		when "1000110010000101" => data_out <= rom_array(35973);
		when "1000110010000110" => data_out <= rom_array(35974);
		when "1000110010000111" => data_out <= rom_array(35975);
		when "1000110010001000" => data_out <= rom_array(35976);
		when "1000110010001001" => data_out <= rom_array(35977);
		when "1000110010001010" => data_out <= rom_array(35978);
		when "1000110010001011" => data_out <= rom_array(35979);
		when "1000110010001100" => data_out <= rom_array(35980);
		when "1000110010001101" => data_out <= rom_array(35981);
		when "1000110010001110" => data_out <= rom_array(35982);
		when "1000110010001111" => data_out <= rom_array(35983);
		when "1000110010010000" => data_out <= rom_array(35984);
		when "1000110010010001" => data_out <= rom_array(35985);
		when "1000110010010010" => data_out <= rom_array(35986);
		when "1000110010010011" => data_out <= rom_array(35987);
		when "1000110010010100" => data_out <= rom_array(35988);
		when "1000110010010101" => data_out <= rom_array(35989);
		when "1000110010010110" => data_out <= rom_array(35990);
		when "1000110010010111" => data_out <= rom_array(35991);
		when "1000110010011000" => data_out <= rom_array(35992);
		when "1000110010011001" => data_out <= rom_array(35993);
		when "1000110010011010" => data_out <= rom_array(35994);
		when "1000110010011011" => data_out <= rom_array(35995);
		when "1000110010011100" => data_out <= rom_array(35996);
		when "1000110010011101" => data_out <= rom_array(35997);
		when "1000110010011110" => data_out <= rom_array(35998);
		when "1000110010011111" => data_out <= rom_array(35999);
		when "1000110010100000" => data_out <= rom_array(36000);
		when "1000110010100001" => data_out <= rom_array(36001);
		when "1000110010100010" => data_out <= rom_array(36002);
		when "1000110010100011" => data_out <= rom_array(36003);
		when "1000110010100100" => data_out <= rom_array(36004);
		when "1000110010100101" => data_out <= rom_array(36005);
		when "1000110010100110" => data_out <= rom_array(36006);
		when "1000110010100111" => data_out <= rom_array(36007);
		when "1000110010101000" => data_out <= rom_array(36008);
		when "1000110010101001" => data_out <= rom_array(36009);
		when "1000110010101010" => data_out <= rom_array(36010);
		when "1000110010101011" => data_out <= rom_array(36011);
		when "1000110010101100" => data_out <= rom_array(36012);
		when "1000110010101101" => data_out <= rom_array(36013);
		when "1000110010101110" => data_out <= rom_array(36014);
		when "1000110010101111" => data_out <= rom_array(36015);
		when "1000110010110000" => data_out <= rom_array(36016);
		when "1000110010110001" => data_out <= rom_array(36017);
		when "1000110010110010" => data_out <= rom_array(36018);
		when "1000110010110011" => data_out <= rom_array(36019);
		when "1000110010110100" => data_out <= rom_array(36020);
		when "1000110010110101" => data_out <= rom_array(36021);
		when "1000110010110110" => data_out <= rom_array(36022);
		when "1000110010110111" => data_out <= rom_array(36023);
		when "1000110010111000" => data_out <= rom_array(36024);
		when "1000110010111001" => data_out <= rom_array(36025);
		when "1000110010111010" => data_out <= rom_array(36026);
		when "1000110010111011" => data_out <= rom_array(36027);
		when "1000110010111100" => data_out <= rom_array(36028);
		when "1000110010111101" => data_out <= rom_array(36029);
		when "1000110010111110" => data_out <= rom_array(36030);
		when "1000110010111111" => data_out <= rom_array(36031);
		when "1000110011000000" => data_out <= rom_array(36032);
		when "1000110011000001" => data_out <= rom_array(36033);
		when "1000110011000010" => data_out <= rom_array(36034);
		when "1000110011000011" => data_out <= rom_array(36035);
		when "1000110011000100" => data_out <= rom_array(36036);
		when "1000110011000101" => data_out <= rom_array(36037);
		when "1000110011000110" => data_out <= rom_array(36038);
		when "1000110011000111" => data_out <= rom_array(36039);
		when "1000110011001000" => data_out <= rom_array(36040);
		when "1000110011001001" => data_out <= rom_array(36041);
		when "1000110011001010" => data_out <= rom_array(36042);
		when "1000110011001011" => data_out <= rom_array(36043);
		when "1000110011001100" => data_out <= rom_array(36044);
		when "1000110011001101" => data_out <= rom_array(36045);
		when "1000110011001110" => data_out <= rom_array(36046);
		when "1000110011001111" => data_out <= rom_array(36047);
		when "1000110011010000" => data_out <= rom_array(36048);
		when "1000110011010001" => data_out <= rom_array(36049);
		when "1000110011010010" => data_out <= rom_array(36050);
		when "1000110011010011" => data_out <= rom_array(36051);
		when "1000110011010100" => data_out <= rom_array(36052);
		when "1000110011010101" => data_out <= rom_array(36053);
		when "1000110011010110" => data_out <= rom_array(36054);
		when "1000110011010111" => data_out <= rom_array(36055);
		when "1000110011011000" => data_out <= rom_array(36056);
		when "1000110011011001" => data_out <= rom_array(36057);
		when "1000110011011010" => data_out <= rom_array(36058);
		when "1000110011011011" => data_out <= rom_array(36059);
		when "1000110011011100" => data_out <= rom_array(36060);
		when "1000110011011101" => data_out <= rom_array(36061);
		when "1000110011011110" => data_out <= rom_array(36062);
		when "1000110011011111" => data_out <= rom_array(36063);
		when "1000110011100000" => data_out <= rom_array(36064);
		when "1000110011100001" => data_out <= rom_array(36065);
		when "1000110011100010" => data_out <= rom_array(36066);
		when "1000110011100011" => data_out <= rom_array(36067);
		when "1000110011100100" => data_out <= rom_array(36068);
		when "1000110011100101" => data_out <= rom_array(36069);
		when "1000110011100110" => data_out <= rom_array(36070);
		when "1000110011100111" => data_out <= rom_array(36071);
		when "1000110011101000" => data_out <= rom_array(36072);
		when "1000110011101001" => data_out <= rom_array(36073);
		when "1000110011101010" => data_out <= rom_array(36074);
		when "1000110011101011" => data_out <= rom_array(36075);
		when "1000110011101100" => data_out <= rom_array(36076);
		when "1000110011101101" => data_out <= rom_array(36077);
		when "1000110011101110" => data_out <= rom_array(36078);
		when "1000110011101111" => data_out <= rom_array(36079);
		when "1000110011110000" => data_out <= rom_array(36080);
		when "1000110011110001" => data_out <= rom_array(36081);
		when "1000110011110010" => data_out <= rom_array(36082);
		when "1000110011110011" => data_out <= rom_array(36083);
		when "1000110011110100" => data_out <= rom_array(36084);
		when "1000110011110101" => data_out <= rom_array(36085);
		when "1000110011110110" => data_out <= rom_array(36086);
		when "1000110011110111" => data_out <= rom_array(36087);
		when "1000110011111000" => data_out <= rom_array(36088);
		when "1000110011111001" => data_out <= rom_array(36089);
		when "1000110011111010" => data_out <= rom_array(36090);
		when "1000110011111011" => data_out <= rom_array(36091);
		when "1000110011111100" => data_out <= rom_array(36092);
		when "1000110011111101" => data_out <= rom_array(36093);
		when "1000110011111110" => data_out <= rom_array(36094);
		when "1000110011111111" => data_out <= rom_array(36095);
		when "1000110100000000" => data_out <= rom_array(36096);
		when "1000110100000001" => data_out <= rom_array(36097);
		when "1000110100000010" => data_out <= rom_array(36098);
		when "1000110100000011" => data_out <= rom_array(36099);
		when "1000110100000100" => data_out <= rom_array(36100);
		when "1000110100000101" => data_out <= rom_array(36101);
		when "1000110100000110" => data_out <= rom_array(36102);
		when "1000110100000111" => data_out <= rom_array(36103);
		when "1000110100001000" => data_out <= rom_array(36104);
		when "1000110100001001" => data_out <= rom_array(36105);
		when "1000110100001010" => data_out <= rom_array(36106);
		when "1000110100001011" => data_out <= rom_array(36107);
		when "1000110100001100" => data_out <= rom_array(36108);
		when "1000110100001101" => data_out <= rom_array(36109);
		when "1000110100001110" => data_out <= rom_array(36110);
		when "1000110100001111" => data_out <= rom_array(36111);
		when "1000110100010000" => data_out <= rom_array(36112);
		when "1000110100010001" => data_out <= rom_array(36113);
		when "1000110100010010" => data_out <= rom_array(36114);
		when "1000110100010011" => data_out <= rom_array(36115);
		when "1000110100010100" => data_out <= rom_array(36116);
		when "1000110100010101" => data_out <= rom_array(36117);
		when "1000110100010110" => data_out <= rom_array(36118);
		when "1000110100010111" => data_out <= rom_array(36119);
		when "1000110100011000" => data_out <= rom_array(36120);
		when "1000110100011001" => data_out <= rom_array(36121);
		when "1000110100011010" => data_out <= rom_array(36122);
		when "1000110100011011" => data_out <= rom_array(36123);
		when "1000110100011100" => data_out <= rom_array(36124);
		when "1000110100011101" => data_out <= rom_array(36125);
		when "1000110100011110" => data_out <= rom_array(36126);
		when "1000110100011111" => data_out <= rom_array(36127);
		when "1000110100100000" => data_out <= rom_array(36128);
		when "1000110100100001" => data_out <= rom_array(36129);
		when "1000110100100010" => data_out <= rom_array(36130);
		when "1000110100100011" => data_out <= rom_array(36131);
		when "1000110100100100" => data_out <= rom_array(36132);
		when "1000110100100101" => data_out <= rom_array(36133);
		when "1000110100100110" => data_out <= rom_array(36134);
		when "1000110100100111" => data_out <= rom_array(36135);
		when "1000110100101000" => data_out <= rom_array(36136);
		when "1000110100101001" => data_out <= rom_array(36137);
		when "1000110100101010" => data_out <= rom_array(36138);
		when "1000110100101011" => data_out <= rom_array(36139);
		when "1000110100101100" => data_out <= rom_array(36140);
		when "1000110100101101" => data_out <= rom_array(36141);
		when "1000110100101110" => data_out <= rom_array(36142);
		when "1000110100101111" => data_out <= rom_array(36143);
		when "1000110100110000" => data_out <= rom_array(36144);
		when "1000110100110001" => data_out <= rom_array(36145);
		when "1000110100110010" => data_out <= rom_array(36146);
		when "1000110100110011" => data_out <= rom_array(36147);
		when "1000110100110100" => data_out <= rom_array(36148);
		when "1000110100110101" => data_out <= rom_array(36149);
		when "1000110100110110" => data_out <= rom_array(36150);
		when "1000110100110111" => data_out <= rom_array(36151);
		when "1000110100111000" => data_out <= rom_array(36152);
		when "1000110100111001" => data_out <= rom_array(36153);
		when "1000110100111010" => data_out <= rom_array(36154);
		when "1000110100111011" => data_out <= rom_array(36155);
		when "1000110100111100" => data_out <= rom_array(36156);
		when "1000110100111101" => data_out <= rom_array(36157);
		when "1000110100111110" => data_out <= rom_array(36158);
		when "1000110100111111" => data_out <= rom_array(36159);
		when "1000110101000000" => data_out <= rom_array(36160);
		when "1000110101000001" => data_out <= rom_array(36161);
		when "1000110101000010" => data_out <= rom_array(36162);
		when "1000110101000011" => data_out <= rom_array(36163);
		when "1000110101000100" => data_out <= rom_array(36164);
		when "1000110101000101" => data_out <= rom_array(36165);
		when "1000110101000110" => data_out <= rom_array(36166);
		when "1000110101000111" => data_out <= rom_array(36167);
		when "1000110101001000" => data_out <= rom_array(36168);
		when "1000110101001001" => data_out <= rom_array(36169);
		when "1000110101001010" => data_out <= rom_array(36170);
		when "1000110101001011" => data_out <= rom_array(36171);
		when "1000110101001100" => data_out <= rom_array(36172);
		when "1000110101001101" => data_out <= rom_array(36173);
		when "1000110101001110" => data_out <= rom_array(36174);
		when "1000110101001111" => data_out <= rom_array(36175);
		when "1000110101010000" => data_out <= rom_array(36176);
		when "1000110101010001" => data_out <= rom_array(36177);
		when "1000110101010010" => data_out <= rom_array(36178);
		when "1000110101010011" => data_out <= rom_array(36179);
		when "1000110101010100" => data_out <= rom_array(36180);
		when "1000110101010101" => data_out <= rom_array(36181);
		when "1000110101010110" => data_out <= rom_array(36182);
		when "1000110101010111" => data_out <= rom_array(36183);
		when "1000110101011000" => data_out <= rom_array(36184);
		when "1000110101011001" => data_out <= rom_array(36185);
		when "1000110101011010" => data_out <= rom_array(36186);
		when "1000110101011011" => data_out <= rom_array(36187);
		when "1000110101011100" => data_out <= rom_array(36188);
		when "1000110101011101" => data_out <= rom_array(36189);
		when "1000110101011110" => data_out <= rom_array(36190);
		when "1000110101011111" => data_out <= rom_array(36191);
		when "1000110101100000" => data_out <= rom_array(36192);
		when "1000110101100001" => data_out <= rom_array(36193);
		when "1000110101100010" => data_out <= rom_array(36194);
		when "1000110101100011" => data_out <= rom_array(36195);
		when "1000110101100100" => data_out <= rom_array(36196);
		when "1000110101100101" => data_out <= rom_array(36197);
		when "1000110101100110" => data_out <= rom_array(36198);
		when "1000110101100111" => data_out <= rom_array(36199);
		when "1000110101101000" => data_out <= rom_array(36200);
		when "1000110101101001" => data_out <= rom_array(36201);
		when "1000110101101010" => data_out <= rom_array(36202);
		when "1000110101101011" => data_out <= rom_array(36203);
		when "1000110101101100" => data_out <= rom_array(36204);
		when "1000110101101101" => data_out <= rom_array(36205);
		when "1000110101101110" => data_out <= rom_array(36206);
		when "1000110101101111" => data_out <= rom_array(36207);
		when "1000110101110000" => data_out <= rom_array(36208);
		when "1000110101110001" => data_out <= rom_array(36209);
		when "1000110101110010" => data_out <= rom_array(36210);
		when "1000110101110011" => data_out <= rom_array(36211);
		when "1000110101110100" => data_out <= rom_array(36212);
		when "1000110101110101" => data_out <= rom_array(36213);
		when "1000110101110110" => data_out <= rom_array(36214);
		when "1000110101110111" => data_out <= rom_array(36215);
		when "1000110101111000" => data_out <= rom_array(36216);
		when "1000110101111001" => data_out <= rom_array(36217);
		when "1000110101111010" => data_out <= rom_array(36218);
		when "1000110101111011" => data_out <= rom_array(36219);
		when "1000110101111100" => data_out <= rom_array(36220);
		when "1000110101111101" => data_out <= rom_array(36221);
		when "1000110101111110" => data_out <= rom_array(36222);
		when "1000110101111111" => data_out <= rom_array(36223);
		when "1000110110000000" => data_out <= rom_array(36224);
		when "1000110110000001" => data_out <= rom_array(36225);
		when "1000110110000010" => data_out <= rom_array(36226);
		when "1000110110000011" => data_out <= rom_array(36227);
		when "1000110110000100" => data_out <= rom_array(36228);
		when "1000110110000101" => data_out <= rom_array(36229);
		when "1000110110000110" => data_out <= rom_array(36230);
		when "1000110110000111" => data_out <= rom_array(36231);
		when "1000110110001000" => data_out <= rom_array(36232);
		when "1000110110001001" => data_out <= rom_array(36233);
		when "1000110110001010" => data_out <= rom_array(36234);
		when "1000110110001011" => data_out <= rom_array(36235);
		when "1000110110001100" => data_out <= rom_array(36236);
		when "1000110110001101" => data_out <= rom_array(36237);
		when "1000110110001110" => data_out <= rom_array(36238);
		when "1000110110001111" => data_out <= rom_array(36239);
		when "1000110110010000" => data_out <= rom_array(36240);
		when "1000110110010001" => data_out <= rom_array(36241);
		when "1000110110010010" => data_out <= rom_array(36242);
		when "1000110110010011" => data_out <= rom_array(36243);
		when "1000110110010100" => data_out <= rom_array(36244);
		when "1000110110010101" => data_out <= rom_array(36245);
		when "1000110110010110" => data_out <= rom_array(36246);
		when "1000110110010111" => data_out <= rom_array(36247);
		when "1000110110011000" => data_out <= rom_array(36248);
		when "1000110110011001" => data_out <= rom_array(36249);
		when "1000110110011010" => data_out <= rom_array(36250);
		when "1000110110011011" => data_out <= rom_array(36251);
		when "1000110110011100" => data_out <= rom_array(36252);
		when "1000110110011101" => data_out <= rom_array(36253);
		when "1000110110011110" => data_out <= rom_array(36254);
		when "1000110110011111" => data_out <= rom_array(36255);
		when "1000110110100000" => data_out <= rom_array(36256);
		when "1000110110100001" => data_out <= rom_array(36257);
		when "1000110110100010" => data_out <= rom_array(36258);
		when "1000110110100011" => data_out <= rom_array(36259);
		when "1000110110100100" => data_out <= rom_array(36260);
		when "1000110110100101" => data_out <= rom_array(36261);
		when "1000110110100110" => data_out <= rom_array(36262);
		when "1000110110100111" => data_out <= rom_array(36263);
		when "1000110110101000" => data_out <= rom_array(36264);
		when "1000110110101001" => data_out <= rom_array(36265);
		when "1000110110101010" => data_out <= rom_array(36266);
		when "1000110110101011" => data_out <= rom_array(36267);
		when "1000110110101100" => data_out <= rom_array(36268);
		when "1000110110101101" => data_out <= rom_array(36269);
		when "1000110110101110" => data_out <= rom_array(36270);
		when "1000110110101111" => data_out <= rom_array(36271);
		when "1000110110110000" => data_out <= rom_array(36272);
		when "1000110110110001" => data_out <= rom_array(36273);
		when "1000110110110010" => data_out <= rom_array(36274);
		when "1000110110110011" => data_out <= rom_array(36275);
		when "1000110110110100" => data_out <= rom_array(36276);
		when "1000110110110101" => data_out <= rom_array(36277);
		when "1000110110110110" => data_out <= rom_array(36278);
		when "1000110110110111" => data_out <= rom_array(36279);
		when "1000110110111000" => data_out <= rom_array(36280);
		when "1000110110111001" => data_out <= rom_array(36281);
		when "1000110110111010" => data_out <= rom_array(36282);
		when "1000110110111011" => data_out <= rom_array(36283);
		when "1000110110111100" => data_out <= rom_array(36284);
		when "1000110110111101" => data_out <= rom_array(36285);
		when "1000110110111110" => data_out <= rom_array(36286);
		when "1000110110111111" => data_out <= rom_array(36287);
		when "1000110111000000" => data_out <= rom_array(36288);
		when "1000110111000001" => data_out <= rom_array(36289);
		when "1000110111000010" => data_out <= rom_array(36290);
		when "1000110111000011" => data_out <= rom_array(36291);
		when "1000110111000100" => data_out <= rom_array(36292);
		when "1000110111000101" => data_out <= rom_array(36293);
		when "1000110111000110" => data_out <= rom_array(36294);
		when "1000110111000111" => data_out <= rom_array(36295);
		when "1000110111001000" => data_out <= rom_array(36296);
		when "1000110111001001" => data_out <= rom_array(36297);
		when "1000110111001010" => data_out <= rom_array(36298);
		when "1000110111001011" => data_out <= rom_array(36299);
		when "1000110111001100" => data_out <= rom_array(36300);
		when "1000110111001101" => data_out <= rom_array(36301);
		when "1000110111001110" => data_out <= rom_array(36302);
		when "1000110111001111" => data_out <= rom_array(36303);
		when "1000110111010000" => data_out <= rom_array(36304);
		when "1000110111010001" => data_out <= rom_array(36305);
		when "1000110111010010" => data_out <= rom_array(36306);
		when "1000110111010011" => data_out <= rom_array(36307);
		when "1000110111010100" => data_out <= rom_array(36308);
		when "1000110111010101" => data_out <= rom_array(36309);
		when "1000110111010110" => data_out <= rom_array(36310);
		when "1000110111010111" => data_out <= rom_array(36311);
		when "1000110111011000" => data_out <= rom_array(36312);
		when "1000110111011001" => data_out <= rom_array(36313);
		when "1000110111011010" => data_out <= rom_array(36314);
		when "1000110111011011" => data_out <= rom_array(36315);
		when "1000110111011100" => data_out <= rom_array(36316);
		when "1000110111011101" => data_out <= rom_array(36317);
		when "1000110111011110" => data_out <= rom_array(36318);
		when "1000110111011111" => data_out <= rom_array(36319);
		when "1000110111100000" => data_out <= rom_array(36320);
		when "1000110111100001" => data_out <= rom_array(36321);
		when "1000110111100010" => data_out <= rom_array(36322);
		when "1000110111100011" => data_out <= rom_array(36323);
		when "1000110111100100" => data_out <= rom_array(36324);
		when "1000110111100101" => data_out <= rom_array(36325);
		when "1000110111100110" => data_out <= rom_array(36326);
		when "1000110111100111" => data_out <= rom_array(36327);
		when "1000110111101000" => data_out <= rom_array(36328);
		when "1000110111101001" => data_out <= rom_array(36329);
		when "1000110111101010" => data_out <= rom_array(36330);
		when "1000110111101011" => data_out <= rom_array(36331);
		when "1000110111101100" => data_out <= rom_array(36332);
		when "1000110111101101" => data_out <= rom_array(36333);
		when "1000110111101110" => data_out <= rom_array(36334);
		when "1000110111101111" => data_out <= rom_array(36335);
		when "1000110111110000" => data_out <= rom_array(36336);
		when "1000110111110001" => data_out <= rom_array(36337);
		when "1000110111110010" => data_out <= rom_array(36338);
		when "1000110111110011" => data_out <= rom_array(36339);
		when "1000110111110100" => data_out <= rom_array(36340);
		when "1000110111110101" => data_out <= rom_array(36341);
		when "1000110111110110" => data_out <= rom_array(36342);
		when "1000110111110111" => data_out <= rom_array(36343);
		when "1000110111111000" => data_out <= rom_array(36344);
		when "1000110111111001" => data_out <= rom_array(36345);
		when "1000110111111010" => data_out <= rom_array(36346);
		when "1000110111111011" => data_out <= rom_array(36347);
		when "1000110111111100" => data_out <= rom_array(36348);
		when "1000110111111101" => data_out <= rom_array(36349);
		when "1000110111111110" => data_out <= rom_array(36350);
		when "1000110111111111" => data_out <= rom_array(36351);
		when "1000111000000000" => data_out <= rom_array(36352);
		when "1000111000000001" => data_out <= rom_array(36353);
		when "1000111000000010" => data_out <= rom_array(36354);
		when "1000111000000011" => data_out <= rom_array(36355);
		when "1000111000000100" => data_out <= rom_array(36356);
		when "1000111000000101" => data_out <= rom_array(36357);
		when "1000111000000110" => data_out <= rom_array(36358);
		when "1000111000000111" => data_out <= rom_array(36359);
		when "1000111000001000" => data_out <= rom_array(36360);
		when "1000111000001001" => data_out <= rom_array(36361);
		when "1000111000001010" => data_out <= rom_array(36362);
		when "1000111000001011" => data_out <= rom_array(36363);
		when "1000111000001100" => data_out <= rom_array(36364);
		when "1000111000001101" => data_out <= rom_array(36365);
		when "1000111000001110" => data_out <= rom_array(36366);
		when "1000111000001111" => data_out <= rom_array(36367);
		when "1000111000010000" => data_out <= rom_array(36368);
		when "1000111000010001" => data_out <= rom_array(36369);
		when "1000111000010010" => data_out <= rom_array(36370);
		when "1000111000010011" => data_out <= rom_array(36371);
		when "1000111000010100" => data_out <= rom_array(36372);
		when "1000111000010101" => data_out <= rom_array(36373);
		when "1000111000010110" => data_out <= rom_array(36374);
		when "1000111000010111" => data_out <= rom_array(36375);
		when "1000111000011000" => data_out <= rom_array(36376);
		when "1000111000011001" => data_out <= rom_array(36377);
		when "1000111000011010" => data_out <= rom_array(36378);
		when "1000111000011011" => data_out <= rom_array(36379);
		when "1000111000011100" => data_out <= rom_array(36380);
		when "1000111000011101" => data_out <= rom_array(36381);
		when "1000111000011110" => data_out <= rom_array(36382);
		when "1000111000011111" => data_out <= rom_array(36383);
		when "1000111000100000" => data_out <= rom_array(36384);
		when "1000111000100001" => data_out <= rom_array(36385);
		when "1000111000100010" => data_out <= rom_array(36386);
		when "1000111000100011" => data_out <= rom_array(36387);
		when "1000111000100100" => data_out <= rom_array(36388);
		when "1000111000100101" => data_out <= rom_array(36389);
		when "1000111000100110" => data_out <= rom_array(36390);
		when "1000111000100111" => data_out <= rom_array(36391);
		when "1000111000101000" => data_out <= rom_array(36392);
		when "1000111000101001" => data_out <= rom_array(36393);
		when "1000111000101010" => data_out <= rom_array(36394);
		when "1000111000101011" => data_out <= rom_array(36395);
		when "1000111000101100" => data_out <= rom_array(36396);
		when "1000111000101101" => data_out <= rom_array(36397);
		when "1000111000101110" => data_out <= rom_array(36398);
		when "1000111000101111" => data_out <= rom_array(36399);
		when "1000111000110000" => data_out <= rom_array(36400);
		when "1000111000110001" => data_out <= rom_array(36401);
		when "1000111000110010" => data_out <= rom_array(36402);
		when "1000111000110011" => data_out <= rom_array(36403);
		when "1000111000110100" => data_out <= rom_array(36404);
		when "1000111000110101" => data_out <= rom_array(36405);
		when "1000111000110110" => data_out <= rom_array(36406);
		when "1000111000110111" => data_out <= rom_array(36407);
		when "1000111000111000" => data_out <= rom_array(36408);
		when "1000111000111001" => data_out <= rom_array(36409);
		when "1000111000111010" => data_out <= rom_array(36410);
		when "1000111000111011" => data_out <= rom_array(36411);
		when "1000111000111100" => data_out <= rom_array(36412);
		when "1000111000111101" => data_out <= rom_array(36413);
		when "1000111000111110" => data_out <= rom_array(36414);
		when "1000111000111111" => data_out <= rom_array(36415);
		when "1000111001000000" => data_out <= rom_array(36416);
		when "1000111001000001" => data_out <= rom_array(36417);
		when "1000111001000010" => data_out <= rom_array(36418);
		when "1000111001000011" => data_out <= rom_array(36419);
		when "1000111001000100" => data_out <= rom_array(36420);
		when "1000111001000101" => data_out <= rom_array(36421);
		when "1000111001000110" => data_out <= rom_array(36422);
		when "1000111001000111" => data_out <= rom_array(36423);
		when "1000111001001000" => data_out <= rom_array(36424);
		when "1000111001001001" => data_out <= rom_array(36425);
		when "1000111001001010" => data_out <= rom_array(36426);
		when "1000111001001011" => data_out <= rom_array(36427);
		when "1000111001001100" => data_out <= rom_array(36428);
		when "1000111001001101" => data_out <= rom_array(36429);
		when "1000111001001110" => data_out <= rom_array(36430);
		when "1000111001001111" => data_out <= rom_array(36431);
		when "1000111001010000" => data_out <= rom_array(36432);
		when "1000111001010001" => data_out <= rom_array(36433);
		when "1000111001010010" => data_out <= rom_array(36434);
		when "1000111001010011" => data_out <= rom_array(36435);
		when "1000111001010100" => data_out <= rom_array(36436);
		when "1000111001010101" => data_out <= rom_array(36437);
		when "1000111001010110" => data_out <= rom_array(36438);
		when "1000111001010111" => data_out <= rom_array(36439);
		when "1000111001011000" => data_out <= rom_array(36440);
		when "1000111001011001" => data_out <= rom_array(36441);
		when "1000111001011010" => data_out <= rom_array(36442);
		when "1000111001011011" => data_out <= rom_array(36443);
		when "1000111001011100" => data_out <= rom_array(36444);
		when "1000111001011101" => data_out <= rom_array(36445);
		when "1000111001011110" => data_out <= rom_array(36446);
		when "1000111001011111" => data_out <= rom_array(36447);
		when "1000111001100000" => data_out <= rom_array(36448);
		when "1000111001100001" => data_out <= rom_array(36449);
		when "1000111001100010" => data_out <= rom_array(36450);
		when "1000111001100011" => data_out <= rom_array(36451);
		when "1000111001100100" => data_out <= rom_array(36452);
		when "1000111001100101" => data_out <= rom_array(36453);
		when "1000111001100110" => data_out <= rom_array(36454);
		when "1000111001100111" => data_out <= rom_array(36455);
		when "1000111001101000" => data_out <= rom_array(36456);
		when "1000111001101001" => data_out <= rom_array(36457);
		when "1000111001101010" => data_out <= rom_array(36458);
		when "1000111001101011" => data_out <= rom_array(36459);
		when "1000111001101100" => data_out <= rom_array(36460);
		when "1000111001101101" => data_out <= rom_array(36461);
		when "1000111001101110" => data_out <= rom_array(36462);
		when "1000111001101111" => data_out <= rom_array(36463);
		when "1000111001110000" => data_out <= rom_array(36464);
		when "1000111001110001" => data_out <= rom_array(36465);
		when "1000111001110010" => data_out <= rom_array(36466);
		when "1000111001110011" => data_out <= rom_array(36467);
		when "1000111001110100" => data_out <= rom_array(36468);
		when "1000111001110101" => data_out <= rom_array(36469);
		when "1000111001110110" => data_out <= rom_array(36470);
		when "1000111001110111" => data_out <= rom_array(36471);
		when "1000111001111000" => data_out <= rom_array(36472);
		when "1000111001111001" => data_out <= rom_array(36473);
		when "1000111001111010" => data_out <= rom_array(36474);
		when "1000111001111011" => data_out <= rom_array(36475);
		when "1000111001111100" => data_out <= rom_array(36476);
		when "1000111001111101" => data_out <= rom_array(36477);
		when "1000111001111110" => data_out <= rom_array(36478);
		when "1000111001111111" => data_out <= rom_array(36479);
		when "1000111010000000" => data_out <= rom_array(36480);
		when "1000111010000001" => data_out <= rom_array(36481);
		when "1000111010000010" => data_out <= rom_array(36482);
		when "1000111010000011" => data_out <= rom_array(36483);
		when "1000111010000100" => data_out <= rom_array(36484);
		when "1000111010000101" => data_out <= rom_array(36485);
		when "1000111010000110" => data_out <= rom_array(36486);
		when "1000111010000111" => data_out <= rom_array(36487);
		when "1000111010001000" => data_out <= rom_array(36488);
		when "1000111010001001" => data_out <= rom_array(36489);
		when "1000111010001010" => data_out <= rom_array(36490);
		when "1000111010001011" => data_out <= rom_array(36491);
		when "1000111010001100" => data_out <= rom_array(36492);
		when "1000111010001101" => data_out <= rom_array(36493);
		when "1000111010001110" => data_out <= rom_array(36494);
		when "1000111010001111" => data_out <= rom_array(36495);
		when "1000111010010000" => data_out <= rom_array(36496);
		when "1000111010010001" => data_out <= rom_array(36497);
		when "1000111010010010" => data_out <= rom_array(36498);
		when "1000111010010011" => data_out <= rom_array(36499);
		when "1000111010010100" => data_out <= rom_array(36500);
		when "1000111010010101" => data_out <= rom_array(36501);
		when "1000111010010110" => data_out <= rom_array(36502);
		when "1000111010010111" => data_out <= rom_array(36503);
		when "1000111010011000" => data_out <= rom_array(36504);
		when "1000111010011001" => data_out <= rom_array(36505);
		when "1000111010011010" => data_out <= rom_array(36506);
		when "1000111010011011" => data_out <= rom_array(36507);
		when "1000111010011100" => data_out <= rom_array(36508);
		when "1000111010011101" => data_out <= rom_array(36509);
		when "1000111010011110" => data_out <= rom_array(36510);
		when "1000111010011111" => data_out <= rom_array(36511);
		when "1000111010100000" => data_out <= rom_array(36512);
		when "1000111010100001" => data_out <= rom_array(36513);
		when "1000111010100010" => data_out <= rom_array(36514);
		when "1000111010100011" => data_out <= rom_array(36515);
		when "1000111010100100" => data_out <= rom_array(36516);
		when "1000111010100101" => data_out <= rom_array(36517);
		when "1000111010100110" => data_out <= rom_array(36518);
		when "1000111010100111" => data_out <= rom_array(36519);
		when "1000111010101000" => data_out <= rom_array(36520);
		when "1000111010101001" => data_out <= rom_array(36521);
		when "1000111010101010" => data_out <= rom_array(36522);
		when "1000111010101011" => data_out <= rom_array(36523);
		when "1000111010101100" => data_out <= rom_array(36524);
		when "1000111010101101" => data_out <= rom_array(36525);
		when "1000111010101110" => data_out <= rom_array(36526);
		when "1000111010101111" => data_out <= rom_array(36527);
		when "1000111010110000" => data_out <= rom_array(36528);
		when "1000111010110001" => data_out <= rom_array(36529);
		when "1000111010110010" => data_out <= rom_array(36530);
		when "1000111010110011" => data_out <= rom_array(36531);
		when "1000111010110100" => data_out <= rom_array(36532);
		when "1000111010110101" => data_out <= rom_array(36533);
		when "1000111010110110" => data_out <= rom_array(36534);
		when "1000111010110111" => data_out <= rom_array(36535);
		when "1000111010111000" => data_out <= rom_array(36536);
		when "1000111010111001" => data_out <= rom_array(36537);
		when "1000111010111010" => data_out <= rom_array(36538);
		when "1000111010111011" => data_out <= rom_array(36539);
		when "1000111010111100" => data_out <= rom_array(36540);
		when "1000111010111101" => data_out <= rom_array(36541);
		when "1000111010111110" => data_out <= rom_array(36542);
		when "1000111010111111" => data_out <= rom_array(36543);
		when "1000111011000000" => data_out <= rom_array(36544);
		when "1000111011000001" => data_out <= rom_array(36545);
		when "1000111011000010" => data_out <= rom_array(36546);
		when "1000111011000011" => data_out <= rom_array(36547);
		when "1000111011000100" => data_out <= rom_array(36548);
		when "1000111011000101" => data_out <= rom_array(36549);
		when "1000111011000110" => data_out <= rom_array(36550);
		when "1000111011000111" => data_out <= rom_array(36551);
		when "1000111011001000" => data_out <= rom_array(36552);
		when "1000111011001001" => data_out <= rom_array(36553);
		when "1000111011001010" => data_out <= rom_array(36554);
		when "1000111011001011" => data_out <= rom_array(36555);
		when "1000111011001100" => data_out <= rom_array(36556);
		when "1000111011001101" => data_out <= rom_array(36557);
		when "1000111011001110" => data_out <= rom_array(36558);
		when "1000111011001111" => data_out <= rom_array(36559);
		when "1000111011010000" => data_out <= rom_array(36560);
		when "1000111011010001" => data_out <= rom_array(36561);
		when "1000111011010010" => data_out <= rom_array(36562);
		when "1000111011010011" => data_out <= rom_array(36563);
		when "1000111011010100" => data_out <= rom_array(36564);
		when "1000111011010101" => data_out <= rom_array(36565);
		when "1000111011010110" => data_out <= rom_array(36566);
		when "1000111011010111" => data_out <= rom_array(36567);
		when "1000111011011000" => data_out <= rom_array(36568);
		when "1000111011011001" => data_out <= rom_array(36569);
		when "1000111011011010" => data_out <= rom_array(36570);
		when "1000111011011011" => data_out <= rom_array(36571);
		when "1000111011011100" => data_out <= rom_array(36572);
		when "1000111011011101" => data_out <= rom_array(36573);
		when "1000111011011110" => data_out <= rom_array(36574);
		when "1000111011011111" => data_out <= rom_array(36575);
		when "1000111011100000" => data_out <= rom_array(36576);
		when "1000111011100001" => data_out <= rom_array(36577);
		when "1000111011100010" => data_out <= rom_array(36578);
		when "1000111011100011" => data_out <= rom_array(36579);
		when "1000111011100100" => data_out <= rom_array(36580);
		when "1000111011100101" => data_out <= rom_array(36581);
		when "1000111011100110" => data_out <= rom_array(36582);
		when "1000111011100111" => data_out <= rom_array(36583);
		when "1000111011101000" => data_out <= rom_array(36584);
		when "1000111011101001" => data_out <= rom_array(36585);
		when "1000111011101010" => data_out <= rom_array(36586);
		when "1000111011101011" => data_out <= rom_array(36587);
		when "1000111011101100" => data_out <= rom_array(36588);
		when "1000111011101101" => data_out <= rom_array(36589);
		when "1000111011101110" => data_out <= rom_array(36590);
		when "1000111011101111" => data_out <= rom_array(36591);
		when "1000111011110000" => data_out <= rom_array(36592);
		when "1000111011110001" => data_out <= rom_array(36593);
		when "1000111011110010" => data_out <= rom_array(36594);
		when "1000111011110011" => data_out <= rom_array(36595);
		when "1000111011110100" => data_out <= rom_array(36596);
		when "1000111011110101" => data_out <= rom_array(36597);
		when "1000111011110110" => data_out <= rom_array(36598);
		when "1000111011110111" => data_out <= rom_array(36599);
		when "1000111011111000" => data_out <= rom_array(36600);
		when "1000111011111001" => data_out <= rom_array(36601);
		when "1000111011111010" => data_out <= rom_array(36602);
		when "1000111011111011" => data_out <= rom_array(36603);
		when "1000111011111100" => data_out <= rom_array(36604);
		when "1000111011111101" => data_out <= rom_array(36605);
		when "1000111011111110" => data_out <= rom_array(36606);
		when "1000111011111111" => data_out <= rom_array(36607);
		when "1000111100000000" => data_out <= rom_array(36608);
		when "1000111100000001" => data_out <= rom_array(36609);
		when "1000111100000010" => data_out <= rom_array(36610);
		when "1000111100000011" => data_out <= rom_array(36611);
		when "1000111100000100" => data_out <= rom_array(36612);
		when "1000111100000101" => data_out <= rom_array(36613);
		when "1000111100000110" => data_out <= rom_array(36614);
		when "1000111100000111" => data_out <= rom_array(36615);
		when "1000111100001000" => data_out <= rom_array(36616);
		when "1000111100001001" => data_out <= rom_array(36617);
		when "1000111100001010" => data_out <= rom_array(36618);
		when "1000111100001011" => data_out <= rom_array(36619);
		when "1000111100001100" => data_out <= rom_array(36620);
		when "1000111100001101" => data_out <= rom_array(36621);
		when "1000111100001110" => data_out <= rom_array(36622);
		when "1000111100001111" => data_out <= rom_array(36623);
		when "1000111100010000" => data_out <= rom_array(36624);
		when "1000111100010001" => data_out <= rom_array(36625);
		when "1000111100010010" => data_out <= rom_array(36626);
		when "1000111100010011" => data_out <= rom_array(36627);
		when "1000111100010100" => data_out <= rom_array(36628);
		when "1000111100010101" => data_out <= rom_array(36629);
		when "1000111100010110" => data_out <= rom_array(36630);
		when "1000111100010111" => data_out <= rom_array(36631);
		when "1000111100011000" => data_out <= rom_array(36632);
		when "1000111100011001" => data_out <= rom_array(36633);
		when "1000111100011010" => data_out <= rom_array(36634);
		when "1000111100011011" => data_out <= rom_array(36635);
		when "1000111100011100" => data_out <= rom_array(36636);
		when "1000111100011101" => data_out <= rom_array(36637);
		when "1000111100011110" => data_out <= rom_array(36638);
		when "1000111100011111" => data_out <= rom_array(36639);
		when "1000111100100000" => data_out <= rom_array(36640);
		when "1000111100100001" => data_out <= rom_array(36641);
		when "1000111100100010" => data_out <= rom_array(36642);
		when "1000111100100011" => data_out <= rom_array(36643);
		when "1000111100100100" => data_out <= rom_array(36644);
		when "1000111100100101" => data_out <= rom_array(36645);
		when "1000111100100110" => data_out <= rom_array(36646);
		when "1000111100100111" => data_out <= rom_array(36647);
		when "1000111100101000" => data_out <= rom_array(36648);
		when "1000111100101001" => data_out <= rom_array(36649);
		when "1000111100101010" => data_out <= rom_array(36650);
		when "1000111100101011" => data_out <= rom_array(36651);
		when "1000111100101100" => data_out <= rom_array(36652);
		when "1000111100101101" => data_out <= rom_array(36653);
		when "1000111100101110" => data_out <= rom_array(36654);
		when "1000111100101111" => data_out <= rom_array(36655);
		when "1000111100110000" => data_out <= rom_array(36656);
		when "1000111100110001" => data_out <= rom_array(36657);
		when "1000111100110010" => data_out <= rom_array(36658);
		when "1000111100110011" => data_out <= rom_array(36659);
		when "1000111100110100" => data_out <= rom_array(36660);
		when "1000111100110101" => data_out <= rom_array(36661);
		when "1000111100110110" => data_out <= rom_array(36662);
		when "1000111100110111" => data_out <= rom_array(36663);
		when "1000111100111000" => data_out <= rom_array(36664);
		when "1000111100111001" => data_out <= rom_array(36665);
		when "1000111100111010" => data_out <= rom_array(36666);
		when "1000111100111011" => data_out <= rom_array(36667);
		when "1000111100111100" => data_out <= rom_array(36668);
		when "1000111100111101" => data_out <= rom_array(36669);
		when "1000111100111110" => data_out <= rom_array(36670);
		when "1000111100111111" => data_out <= rom_array(36671);
		when "1000111101000000" => data_out <= rom_array(36672);
		when "1000111101000001" => data_out <= rom_array(36673);
		when "1000111101000010" => data_out <= rom_array(36674);
		when "1000111101000011" => data_out <= rom_array(36675);
		when "1000111101000100" => data_out <= rom_array(36676);
		when "1000111101000101" => data_out <= rom_array(36677);
		when "1000111101000110" => data_out <= rom_array(36678);
		when "1000111101000111" => data_out <= rom_array(36679);
		when "1000111101001000" => data_out <= rom_array(36680);
		when "1000111101001001" => data_out <= rom_array(36681);
		when "1000111101001010" => data_out <= rom_array(36682);
		when "1000111101001011" => data_out <= rom_array(36683);
		when "1000111101001100" => data_out <= rom_array(36684);
		when "1000111101001101" => data_out <= rom_array(36685);
		when "1000111101001110" => data_out <= rom_array(36686);
		when "1000111101001111" => data_out <= rom_array(36687);
		when "1000111101010000" => data_out <= rom_array(36688);
		when "1000111101010001" => data_out <= rom_array(36689);
		when "1000111101010010" => data_out <= rom_array(36690);
		when "1000111101010011" => data_out <= rom_array(36691);
		when "1000111101010100" => data_out <= rom_array(36692);
		when "1000111101010101" => data_out <= rom_array(36693);
		when "1000111101010110" => data_out <= rom_array(36694);
		when "1000111101010111" => data_out <= rom_array(36695);
		when "1000111101011000" => data_out <= rom_array(36696);
		when "1000111101011001" => data_out <= rom_array(36697);
		when "1000111101011010" => data_out <= rom_array(36698);
		when "1000111101011011" => data_out <= rom_array(36699);
		when "1000111101011100" => data_out <= rom_array(36700);
		when "1000111101011101" => data_out <= rom_array(36701);
		when "1000111101011110" => data_out <= rom_array(36702);
		when "1000111101011111" => data_out <= rom_array(36703);
		when "1000111101100000" => data_out <= rom_array(36704);
		when "1000111101100001" => data_out <= rom_array(36705);
		when "1000111101100010" => data_out <= rom_array(36706);
		when "1000111101100011" => data_out <= rom_array(36707);
		when "1000111101100100" => data_out <= rom_array(36708);
		when "1000111101100101" => data_out <= rom_array(36709);
		when "1000111101100110" => data_out <= rom_array(36710);
		when "1000111101100111" => data_out <= rom_array(36711);
		when "1000111101101000" => data_out <= rom_array(36712);
		when "1000111101101001" => data_out <= rom_array(36713);
		when "1000111101101010" => data_out <= rom_array(36714);
		when "1000111101101011" => data_out <= rom_array(36715);
		when "1000111101101100" => data_out <= rom_array(36716);
		when "1000111101101101" => data_out <= rom_array(36717);
		when "1000111101101110" => data_out <= rom_array(36718);
		when "1000111101101111" => data_out <= rom_array(36719);
		when "1000111101110000" => data_out <= rom_array(36720);
		when "1000111101110001" => data_out <= rom_array(36721);
		when "1000111101110010" => data_out <= rom_array(36722);
		when "1000111101110011" => data_out <= rom_array(36723);
		when "1000111101110100" => data_out <= rom_array(36724);
		when "1000111101110101" => data_out <= rom_array(36725);
		when "1000111101110110" => data_out <= rom_array(36726);
		when "1000111101110111" => data_out <= rom_array(36727);
		when "1000111101111000" => data_out <= rom_array(36728);
		when "1000111101111001" => data_out <= rom_array(36729);
		when "1000111101111010" => data_out <= rom_array(36730);
		when "1000111101111011" => data_out <= rom_array(36731);
		when "1000111101111100" => data_out <= rom_array(36732);
		when "1000111101111101" => data_out <= rom_array(36733);
		when "1000111101111110" => data_out <= rom_array(36734);
		when "1000111101111111" => data_out <= rom_array(36735);
		when "1000111110000000" => data_out <= rom_array(36736);
		when "1000111110000001" => data_out <= rom_array(36737);
		when "1000111110000010" => data_out <= rom_array(36738);
		when "1000111110000011" => data_out <= rom_array(36739);
		when "1000111110000100" => data_out <= rom_array(36740);
		when "1000111110000101" => data_out <= rom_array(36741);
		when "1000111110000110" => data_out <= rom_array(36742);
		when "1000111110000111" => data_out <= rom_array(36743);
		when "1000111110001000" => data_out <= rom_array(36744);
		when "1000111110001001" => data_out <= rom_array(36745);
		when "1000111110001010" => data_out <= rom_array(36746);
		when "1000111110001011" => data_out <= rom_array(36747);
		when "1000111110001100" => data_out <= rom_array(36748);
		when "1000111110001101" => data_out <= rom_array(36749);
		when "1000111110001110" => data_out <= rom_array(36750);
		when "1000111110001111" => data_out <= rom_array(36751);
		when "1000111110010000" => data_out <= rom_array(36752);
		when "1000111110010001" => data_out <= rom_array(36753);
		when "1000111110010010" => data_out <= rom_array(36754);
		when "1000111110010011" => data_out <= rom_array(36755);
		when "1000111110010100" => data_out <= rom_array(36756);
		when "1000111110010101" => data_out <= rom_array(36757);
		when "1000111110010110" => data_out <= rom_array(36758);
		when "1000111110010111" => data_out <= rom_array(36759);
		when "1000111110011000" => data_out <= rom_array(36760);
		when "1000111110011001" => data_out <= rom_array(36761);
		when "1000111110011010" => data_out <= rom_array(36762);
		when "1000111110011011" => data_out <= rom_array(36763);
		when "1000111110011100" => data_out <= rom_array(36764);
		when "1000111110011101" => data_out <= rom_array(36765);
		when "1000111110011110" => data_out <= rom_array(36766);
		when "1000111110011111" => data_out <= rom_array(36767);
		when "1000111110100000" => data_out <= rom_array(36768);
		when "1000111110100001" => data_out <= rom_array(36769);
		when "1000111110100010" => data_out <= rom_array(36770);
		when "1000111110100011" => data_out <= rom_array(36771);
		when "1000111110100100" => data_out <= rom_array(36772);
		when "1000111110100101" => data_out <= rom_array(36773);
		when "1000111110100110" => data_out <= rom_array(36774);
		when "1000111110100111" => data_out <= rom_array(36775);
		when "1000111110101000" => data_out <= rom_array(36776);
		when "1000111110101001" => data_out <= rom_array(36777);
		when "1000111110101010" => data_out <= rom_array(36778);
		when "1000111110101011" => data_out <= rom_array(36779);
		when "1000111110101100" => data_out <= rom_array(36780);
		when "1000111110101101" => data_out <= rom_array(36781);
		when "1000111110101110" => data_out <= rom_array(36782);
		when "1000111110101111" => data_out <= rom_array(36783);
		when "1000111110110000" => data_out <= rom_array(36784);
		when "1000111110110001" => data_out <= rom_array(36785);
		when "1000111110110010" => data_out <= rom_array(36786);
		when "1000111110110011" => data_out <= rom_array(36787);
		when "1000111110110100" => data_out <= rom_array(36788);
		when "1000111110110101" => data_out <= rom_array(36789);
		when "1000111110110110" => data_out <= rom_array(36790);
		when "1000111110110111" => data_out <= rom_array(36791);
		when "1000111110111000" => data_out <= rom_array(36792);
		when "1000111110111001" => data_out <= rom_array(36793);
		when "1000111110111010" => data_out <= rom_array(36794);
		when "1000111110111011" => data_out <= rom_array(36795);
		when "1000111110111100" => data_out <= rom_array(36796);
		when "1000111110111101" => data_out <= rom_array(36797);
		when "1000111110111110" => data_out <= rom_array(36798);
		when "1000111110111111" => data_out <= rom_array(36799);
		when "1000111111000000" => data_out <= rom_array(36800);
		when "1000111111000001" => data_out <= rom_array(36801);
		when "1000111111000010" => data_out <= rom_array(36802);
		when "1000111111000011" => data_out <= rom_array(36803);
		when "1000111111000100" => data_out <= rom_array(36804);
		when "1000111111000101" => data_out <= rom_array(36805);
		when "1000111111000110" => data_out <= rom_array(36806);
		when "1000111111000111" => data_out <= rom_array(36807);
		when "1000111111001000" => data_out <= rom_array(36808);
		when "1000111111001001" => data_out <= rom_array(36809);
		when "1000111111001010" => data_out <= rom_array(36810);
		when "1000111111001011" => data_out <= rom_array(36811);
		when "1000111111001100" => data_out <= rom_array(36812);
		when "1000111111001101" => data_out <= rom_array(36813);
		when "1000111111001110" => data_out <= rom_array(36814);
		when "1000111111001111" => data_out <= rom_array(36815);
		when "1000111111010000" => data_out <= rom_array(36816);
		when "1000111111010001" => data_out <= rom_array(36817);
		when "1000111111010010" => data_out <= rom_array(36818);
		when "1000111111010011" => data_out <= rom_array(36819);
		when "1000111111010100" => data_out <= rom_array(36820);
		when "1000111111010101" => data_out <= rom_array(36821);
		when "1000111111010110" => data_out <= rom_array(36822);
		when "1000111111010111" => data_out <= rom_array(36823);
		when "1000111111011000" => data_out <= rom_array(36824);
		when "1000111111011001" => data_out <= rom_array(36825);
		when "1000111111011010" => data_out <= rom_array(36826);
		when "1000111111011011" => data_out <= rom_array(36827);
		when "1000111111011100" => data_out <= rom_array(36828);
		when "1000111111011101" => data_out <= rom_array(36829);
		when "1000111111011110" => data_out <= rom_array(36830);
		when "1000111111011111" => data_out <= rom_array(36831);
		when "1000111111100000" => data_out <= rom_array(36832);
		when "1000111111100001" => data_out <= rom_array(36833);
		when "1000111111100010" => data_out <= rom_array(36834);
		when "1000111111100011" => data_out <= rom_array(36835);
		when "1000111111100100" => data_out <= rom_array(36836);
		when "1000111111100101" => data_out <= rom_array(36837);
		when "1000111111100110" => data_out <= rom_array(36838);
		when "1000111111100111" => data_out <= rom_array(36839);
		when "1000111111101000" => data_out <= rom_array(36840);
		when "1000111111101001" => data_out <= rom_array(36841);
		when "1000111111101010" => data_out <= rom_array(36842);
		when "1000111111101011" => data_out <= rom_array(36843);
		when "1000111111101100" => data_out <= rom_array(36844);
		when "1000111111101101" => data_out <= rom_array(36845);
		when "1000111111101110" => data_out <= rom_array(36846);
		when "1000111111101111" => data_out <= rom_array(36847);
		when "1000111111110000" => data_out <= rom_array(36848);
		when "1000111111110001" => data_out <= rom_array(36849);
		when "1000111111110010" => data_out <= rom_array(36850);
		when "1000111111110011" => data_out <= rom_array(36851);
		when "1000111111110100" => data_out <= rom_array(36852);
		when "1000111111110101" => data_out <= rom_array(36853);
		when "1000111111110110" => data_out <= rom_array(36854);
		when "1000111111110111" => data_out <= rom_array(36855);
		when "1000111111111000" => data_out <= rom_array(36856);
		when "1000111111111001" => data_out <= rom_array(36857);
		when "1000111111111010" => data_out <= rom_array(36858);
		when "1000111111111011" => data_out <= rom_array(36859);
		when "1000111111111100" => data_out <= rom_array(36860);
		when "1000111111111101" => data_out <= rom_array(36861);
		when "1000111111111110" => data_out <= rom_array(36862);
		when "1000111111111111" => data_out <= rom_array(36863);
		when "1001000000000000" => data_out <= rom_array(36864);
		when "1001000000000001" => data_out <= rom_array(36865);
		when "1001000000000010" => data_out <= rom_array(36866);
		when "1001000000000011" => data_out <= rom_array(36867);
		when "1001000000000100" => data_out <= rom_array(36868);
		when "1001000000000101" => data_out <= rom_array(36869);
		when "1001000000000110" => data_out <= rom_array(36870);
		when "1001000000000111" => data_out <= rom_array(36871);
		when "1001000000001000" => data_out <= rom_array(36872);
		when "1001000000001001" => data_out <= rom_array(36873);
		when "1001000000001010" => data_out <= rom_array(36874);
		when "1001000000001011" => data_out <= rom_array(36875);
		when "1001000000001100" => data_out <= rom_array(36876);
		when "1001000000001101" => data_out <= rom_array(36877);
		when "1001000000001110" => data_out <= rom_array(36878);
		when "1001000000001111" => data_out <= rom_array(36879);
		when "1001000000010000" => data_out <= rom_array(36880);
		when "1001000000010001" => data_out <= rom_array(36881);
		when "1001000000010010" => data_out <= rom_array(36882);
		when "1001000000010011" => data_out <= rom_array(36883);
		when "1001000000010100" => data_out <= rom_array(36884);
		when "1001000000010101" => data_out <= rom_array(36885);
		when "1001000000010110" => data_out <= rom_array(36886);
		when "1001000000010111" => data_out <= rom_array(36887);
		when "1001000000011000" => data_out <= rom_array(36888);
		when "1001000000011001" => data_out <= rom_array(36889);
		when "1001000000011010" => data_out <= rom_array(36890);
		when "1001000000011011" => data_out <= rom_array(36891);
		when "1001000000011100" => data_out <= rom_array(36892);
		when "1001000000011101" => data_out <= rom_array(36893);
		when "1001000000011110" => data_out <= rom_array(36894);
		when "1001000000011111" => data_out <= rom_array(36895);
		when "1001000000100000" => data_out <= rom_array(36896);
		when "1001000000100001" => data_out <= rom_array(36897);
		when "1001000000100010" => data_out <= rom_array(36898);
		when "1001000000100011" => data_out <= rom_array(36899);
		when "1001000000100100" => data_out <= rom_array(36900);
		when "1001000000100101" => data_out <= rom_array(36901);
		when "1001000000100110" => data_out <= rom_array(36902);
		when "1001000000100111" => data_out <= rom_array(36903);
		when "1001000000101000" => data_out <= rom_array(36904);
		when "1001000000101001" => data_out <= rom_array(36905);
		when "1001000000101010" => data_out <= rom_array(36906);
		when "1001000000101011" => data_out <= rom_array(36907);
		when "1001000000101100" => data_out <= rom_array(36908);
		when "1001000000101101" => data_out <= rom_array(36909);
		when "1001000000101110" => data_out <= rom_array(36910);
		when "1001000000101111" => data_out <= rom_array(36911);
		when "1001000000110000" => data_out <= rom_array(36912);
		when "1001000000110001" => data_out <= rom_array(36913);
		when "1001000000110010" => data_out <= rom_array(36914);
		when "1001000000110011" => data_out <= rom_array(36915);
		when "1001000000110100" => data_out <= rom_array(36916);
		when "1001000000110101" => data_out <= rom_array(36917);
		when "1001000000110110" => data_out <= rom_array(36918);
		when "1001000000110111" => data_out <= rom_array(36919);
		when "1001000000111000" => data_out <= rom_array(36920);
		when "1001000000111001" => data_out <= rom_array(36921);
		when "1001000000111010" => data_out <= rom_array(36922);
		when "1001000000111011" => data_out <= rom_array(36923);
		when "1001000000111100" => data_out <= rom_array(36924);
		when "1001000000111101" => data_out <= rom_array(36925);
		when "1001000000111110" => data_out <= rom_array(36926);
		when "1001000000111111" => data_out <= rom_array(36927);
		when "1001000001000000" => data_out <= rom_array(36928);
		when "1001000001000001" => data_out <= rom_array(36929);
		when "1001000001000010" => data_out <= rom_array(36930);
		when "1001000001000011" => data_out <= rom_array(36931);
		when "1001000001000100" => data_out <= rom_array(36932);
		when "1001000001000101" => data_out <= rom_array(36933);
		when "1001000001000110" => data_out <= rom_array(36934);
		when "1001000001000111" => data_out <= rom_array(36935);
		when "1001000001001000" => data_out <= rom_array(36936);
		when "1001000001001001" => data_out <= rom_array(36937);
		when "1001000001001010" => data_out <= rom_array(36938);
		when "1001000001001011" => data_out <= rom_array(36939);
		when "1001000001001100" => data_out <= rom_array(36940);
		when "1001000001001101" => data_out <= rom_array(36941);
		when "1001000001001110" => data_out <= rom_array(36942);
		when "1001000001001111" => data_out <= rom_array(36943);
		when "1001000001010000" => data_out <= rom_array(36944);
		when "1001000001010001" => data_out <= rom_array(36945);
		when "1001000001010010" => data_out <= rom_array(36946);
		when "1001000001010011" => data_out <= rom_array(36947);
		when "1001000001010100" => data_out <= rom_array(36948);
		when "1001000001010101" => data_out <= rom_array(36949);
		when "1001000001010110" => data_out <= rom_array(36950);
		when "1001000001010111" => data_out <= rom_array(36951);
		when "1001000001011000" => data_out <= rom_array(36952);
		when "1001000001011001" => data_out <= rom_array(36953);
		when "1001000001011010" => data_out <= rom_array(36954);
		when "1001000001011011" => data_out <= rom_array(36955);
		when "1001000001011100" => data_out <= rom_array(36956);
		when "1001000001011101" => data_out <= rom_array(36957);
		when "1001000001011110" => data_out <= rom_array(36958);
		when "1001000001011111" => data_out <= rom_array(36959);
		when "1001000001100000" => data_out <= rom_array(36960);
		when "1001000001100001" => data_out <= rom_array(36961);
		when "1001000001100010" => data_out <= rom_array(36962);
		when "1001000001100011" => data_out <= rom_array(36963);
		when "1001000001100100" => data_out <= rom_array(36964);
		when "1001000001100101" => data_out <= rom_array(36965);
		when "1001000001100110" => data_out <= rom_array(36966);
		when "1001000001100111" => data_out <= rom_array(36967);
		when "1001000001101000" => data_out <= rom_array(36968);
		when "1001000001101001" => data_out <= rom_array(36969);
		when "1001000001101010" => data_out <= rom_array(36970);
		when "1001000001101011" => data_out <= rom_array(36971);
		when "1001000001101100" => data_out <= rom_array(36972);
		when "1001000001101101" => data_out <= rom_array(36973);
		when "1001000001101110" => data_out <= rom_array(36974);
		when "1001000001101111" => data_out <= rom_array(36975);
		when "1001000001110000" => data_out <= rom_array(36976);
		when "1001000001110001" => data_out <= rom_array(36977);
		when "1001000001110010" => data_out <= rom_array(36978);
		when "1001000001110011" => data_out <= rom_array(36979);
		when "1001000001110100" => data_out <= rom_array(36980);
		when "1001000001110101" => data_out <= rom_array(36981);
		when "1001000001110110" => data_out <= rom_array(36982);
		when "1001000001110111" => data_out <= rom_array(36983);
		when "1001000001111000" => data_out <= rom_array(36984);
		when "1001000001111001" => data_out <= rom_array(36985);
		when "1001000001111010" => data_out <= rom_array(36986);
		when "1001000001111011" => data_out <= rom_array(36987);
		when "1001000001111100" => data_out <= rom_array(36988);
		when "1001000001111101" => data_out <= rom_array(36989);
		when "1001000001111110" => data_out <= rom_array(36990);
		when "1001000001111111" => data_out <= rom_array(36991);
		when "1001000010000000" => data_out <= rom_array(36992);
		when "1001000010000001" => data_out <= rom_array(36993);
		when "1001000010000010" => data_out <= rom_array(36994);
		when "1001000010000011" => data_out <= rom_array(36995);
		when "1001000010000100" => data_out <= rom_array(36996);
		when "1001000010000101" => data_out <= rom_array(36997);
		when "1001000010000110" => data_out <= rom_array(36998);
		when "1001000010000111" => data_out <= rom_array(36999);
		when "1001000010001000" => data_out <= rom_array(37000);
		when "1001000010001001" => data_out <= rom_array(37001);
		when "1001000010001010" => data_out <= rom_array(37002);
		when "1001000010001011" => data_out <= rom_array(37003);
		when "1001000010001100" => data_out <= rom_array(37004);
		when "1001000010001101" => data_out <= rom_array(37005);
		when "1001000010001110" => data_out <= rom_array(37006);
		when "1001000010001111" => data_out <= rom_array(37007);
		when "1001000010010000" => data_out <= rom_array(37008);
		when "1001000010010001" => data_out <= rom_array(37009);
		when "1001000010010010" => data_out <= rom_array(37010);
		when "1001000010010011" => data_out <= rom_array(37011);
		when "1001000010010100" => data_out <= rom_array(37012);
		when "1001000010010101" => data_out <= rom_array(37013);
		when "1001000010010110" => data_out <= rom_array(37014);
		when "1001000010010111" => data_out <= rom_array(37015);
		when "1001000010011000" => data_out <= rom_array(37016);
		when "1001000010011001" => data_out <= rom_array(37017);
		when "1001000010011010" => data_out <= rom_array(37018);
		when "1001000010011011" => data_out <= rom_array(37019);
		when "1001000010011100" => data_out <= rom_array(37020);
		when "1001000010011101" => data_out <= rom_array(37021);
		when "1001000010011110" => data_out <= rom_array(37022);
		when "1001000010011111" => data_out <= rom_array(37023);
		when "1001000010100000" => data_out <= rom_array(37024);
		when "1001000010100001" => data_out <= rom_array(37025);
		when "1001000010100010" => data_out <= rom_array(37026);
		when "1001000010100011" => data_out <= rom_array(37027);
		when "1001000010100100" => data_out <= rom_array(37028);
		when "1001000010100101" => data_out <= rom_array(37029);
		when "1001000010100110" => data_out <= rom_array(37030);
		when "1001000010100111" => data_out <= rom_array(37031);
		when "1001000010101000" => data_out <= rom_array(37032);
		when "1001000010101001" => data_out <= rom_array(37033);
		when "1001000010101010" => data_out <= rom_array(37034);
		when "1001000010101011" => data_out <= rom_array(37035);
		when "1001000010101100" => data_out <= rom_array(37036);
		when "1001000010101101" => data_out <= rom_array(37037);
		when "1001000010101110" => data_out <= rom_array(37038);
		when "1001000010101111" => data_out <= rom_array(37039);
		when "1001000010110000" => data_out <= rom_array(37040);
		when "1001000010110001" => data_out <= rom_array(37041);
		when "1001000010110010" => data_out <= rom_array(37042);
		when "1001000010110011" => data_out <= rom_array(37043);
		when "1001000010110100" => data_out <= rom_array(37044);
		when "1001000010110101" => data_out <= rom_array(37045);
		when "1001000010110110" => data_out <= rom_array(37046);
		when "1001000010110111" => data_out <= rom_array(37047);
		when "1001000010111000" => data_out <= rom_array(37048);
		when "1001000010111001" => data_out <= rom_array(37049);
		when "1001000010111010" => data_out <= rom_array(37050);
		when "1001000010111011" => data_out <= rom_array(37051);
		when "1001000010111100" => data_out <= rom_array(37052);
		when "1001000010111101" => data_out <= rom_array(37053);
		when "1001000010111110" => data_out <= rom_array(37054);
		when "1001000010111111" => data_out <= rom_array(37055);
		when "1001000011000000" => data_out <= rom_array(37056);
		when "1001000011000001" => data_out <= rom_array(37057);
		when "1001000011000010" => data_out <= rom_array(37058);
		when "1001000011000011" => data_out <= rom_array(37059);
		when "1001000011000100" => data_out <= rom_array(37060);
		when "1001000011000101" => data_out <= rom_array(37061);
		when "1001000011000110" => data_out <= rom_array(37062);
		when "1001000011000111" => data_out <= rom_array(37063);
		when "1001000011001000" => data_out <= rom_array(37064);
		when "1001000011001001" => data_out <= rom_array(37065);
		when "1001000011001010" => data_out <= rom_array(37066);
		when "1001000011001011" => data_out <= rom_array(37067);
		when "1001000011001100" => data_out <= rom_array(37068);
		when "1001000011001101" => data_out <= rom_array(37069);
		when "1001000011001110" => data_out <= rom_array(37070);
		when "1001000011001111" => data_out <= rom_array(37071);
		when "1001000011010000" => data_out <= rom_array(37072);
		when "1001000011010001" => data_out <= rom_array(37073);
		when "1001000011010010" => data_out <= rom_array(37074);
		when "1001000011010011" => data_out <= rom_array(37075);
		when "1001000011010100" => data_out <= rom_array(37076);
		when "1001000011010101" => data_out <= rom_array(37077);
		when "1001000011010110" => data_out <= rom_array(37078);
		when "1001000011010111" => data_out <= rom_array(37079);
		when "1001000011011000" => data_out <= rom_array(37080);
		when "1001000011011001" => data_out <= rom_array(37081);
		when "1001000011011010" => data_out <= rom_array(37082);
		when "1001000011011011" => data_out <= rom_array(37083);
		when "1001000011011100" => data_out <= rom_array(37084);
		when "1001000011011101" => data_out <= rom_array(37085);
		when "1001000011011110" => data_out <= rom_array(37086);
		when "1001000011011111" => data_out <= rom_array(37087);
		when "1001000011100000" => data_out <= rom_array(37088);
		when "1001000011100001" => data_out <= rom_array(37089);
		when "1001000011100010" => data_out <= rom_array(37090);
		when "1001000011100011" => data_out <= rom_array(37091);
		when "1001000011100100" => data_out <= rom_array(37092);
		when "1001000011100101" => data_out <= rom_array(37093);
		when "1001000011100110" => data_out <= rom_array(37094);
		when "1001000011100111" => data_out <= rom_array(37095);
		when "1001000011101000" => data_out <= rom_array(37096);
		when "1001000011101001" => data_out <= rom_array(37097);
		when "1001000011101010" => data_out <= rom_array(37098);
		when "1001000011101011" => data_out <= rom_array(37099);
		when "1001000011101100" => data_out <= rom_array(37100);
		when "1001000011101101" => data_out <= rom_array(37101);
		when "1001000011101110" => data_out <= rom_array(37102);
		when "1001000011101111" => data_out <= rom_array(37103);
		when "1001000011110000" => data_out <= rom_array(37104);
		when "1001000011110001" => data_out <= rom_array(37105);
		when "1001000011110010" => data_out <= rom_array(37106);
		when "1001000011110011" => data_out <= rom_array(37107);
		when "1001000011110100" => data_out <= rom_array(37108);
		when "1001000011110101" => data_out <= rom_array(37109);
		when "1001000011110110" => data_out <= rom_array(37110);
		when "1001000011110111" => data_out <= rom_array(37111);
		when "1001000011111000" => data_out <= rom_array(37112);
		when "1001000011111001" => data_out <= rom_array(37113);
		when "1001000011111010" => data_out <= rom_array(37114);
		when "1001000011111011" => data_out <= rom_array(37115);
		when "1001000011111100" => data_out <= rom_array(37116);
		when "1001000011111101" => data_out <= rom_array(37117);
		when "1001000011111110" => data_out <= rom_array(37118);
		when "1001000011111111" => data_out <= rom_array(37119);
		when "1001000100000000" => data_out <= rom_array(37120);
		when "1001000100000001" => data_out <= rom_array(37121);
		when "1001000100000010" => data_out <= rom_array(37122);
		when "1001000100000011" => data_out <= rom_array(37123);
		when "1001000100000100" => data_out <= rom_array(37124);
		when "1001000100000101" => data_out <= rom_array(37125);
		when "1001000100000110" => data_out <= rom_array(37126);
		when "1001000100000111" => data_out <= rom_array(37127);
		when "1001000100001000" => data_out <= rom_array(37128);
		when "1001000100001001" => data_out <= rom_array(37129);
		when "1001000100001010" => data_out <= rom_array(37130);
		when "1001000100001011" => data_out <= rom_array(37131);
		when "1001000100001100" => data_out <= rom_array(37132);
		when "1001000100001101" => data_out <= rom_array(37133);
		when "1001000100001110" => data_out <= rom_array(37134);
		when "1001000100001111" => data_out <= rom_array(37135);
		when "1001000100010000" => data_out <= rom_array(37136);
		when "1001000100010001" => data_out <= rom_array(37137);
		when "1001000100010010" => data_out <= rom_array(37138);
		when "1001000100010011" => data_out <= rom_array(37139);
		when "1001000100010100" => data_out <= rom_array(37140);
		when "1001000100010101" => data_out <= rom_array(37141);
		when "1001000100010110" => data_out <= rom_array(37142);
		when "1001000100010111" => data_out <= rom_array(37143);
		when "1001000100011000" => data_out <= rom_array(37144);
		when "1001000100011001" => data_out <= rom_array(37145);
		when "1001000100011010" => data_out <= rom_array(37146);
		when "1001000100011011" => data_out <= rom_array(37147);
		when "1001000100011100" => data_out <= rom_array(37148);
		when "1001000100011101" => data_out <= rom_array(37149);
		when "1001000100011110" => data_out <= rom_array(37150);
		when "1001000100011111" => data_out <= rom_array(37151);
		when "1001000100100000" => data_out <= rom_array(37152);
		when "1001000100100001" => data_out <= rom_array(37153);
		when "1001000100100010" => data_out <= rom_array(37154);
		when "1001000100100011" => data_out <= rom_array(37155);
		when "1001000100100100" => data_out <= rom_array(37156);
		when "1001000100100101" => data_out <= rom_array(37157);
		when "1001000100100110" => data_out <= rom_array(37158);
		when "1001000100100111" => data_out <= rom_array(37159);
		when "1001000100101000" => data_out <= rom_array(37160);
		when "1001000100101001" => data_out <= rom_array(37161);
		when "1001000100101010" => data_out <= rom_array(37162);
		when "1001000100101011" => data_out <= rom_array(37163);
		when "1001000100101100" => data_out <= rom_array(37164);
		when "1001000100101101" => data_out <= rom_array(37165);
		when "1001000100101110" => data_out <= rom_array(37166);
		when "1001000100101111" => data_out <= rom_array(37167);
		when "1001000100110000" => data_out <= rom_array(37168);
		when "1001000100110001" => data_out <= rom_array(37169);
		when "1001000100110010" => data_out <= rom_array(37170);
		when "1001000100110011" => data_out <= rom_array(37171);
		when "1001000100110100" => data_out <= rom_array(37172);
		when "1001000100110101" => data_out <= rom_array(37173);
		when "1001000100110110" => data_out <= rom_array(37174);
		when "1001000100110111" => data_out <= rom_array(37175);
		when "1001000100111000" => data_out <= rom_array(37176);
		when "1001000100111001" => data_out <= rom_array(37177);
		when "1001000100111010" => data_out <= rom_array(37178);
		when "1001000100111011" => data_out <= rom_array(37179);
		when "1001000100111100" => data_out <= rom_array(37180);
		when "1001000100111101" => data_out <= rom_array(37181);
		when "1001000100111110" => data_out <= rom_array(37182);
		when "1001000100111111" => data_out <= rom_array(37183);
		when "1001000101000000" => data_out <= rom_array(37184);
		when "1001000101000001" => data_out <= rom_array(37185);
		when "1001000101000010" => data_out <= rom_array(37186);
		when "1001000101000011" => data_out <= rom_array(37187);
		when "1001000101000100" => data_out <= rom_array(37188);
		when "1001000101000101" => data_out <= rom_array(37189);
		when "1001000101000110" => data_out <= rom_array(37190);
		when "1001000101000111" => data_out <= rom_array(37191);
		when "1001000101001000" => data_out <= rom_array(37192);
		when "1001000101001001" => data_out <= rom_array(37193);
		when "1001000101001010" => data_out <= rom_array(37194);
		when "1001000101001011" => data_out <= rom_array(37195);
		when "1001000101001100" => data_out <= rom_array(37196);
		when "1001000101001101" => data_out <= rom_array(37197);
		when "1001000101001110" => data_out <= rom_array(37198);
		when "1001000101001111" => data_out <= rom_array(37199);
		when "1001000101010000" => data_out <= rom_array(37200);
		when "1001000101010001" => data_out <= rom_array(37201);
		when "1001000101010010" => data_out <= rom_array(37202);
		when "1001000101010011" => data_out <= rom_array(37203);
		when "1001000101010100" => data_out <= rom_array(37204);
		when "1001000101010101" => data_out <= rom_array(37205);
		when "1001000101010110" => data_out <= rom_array(37206);
		when "1001000101010111" => data_out <= rom_array(37207);
		when "1001000101011000" => data_out <= rom_array(37208);
		when "1001000101011001" => data_out <= rom_array(37209);
		when "1001000101011010" => data_out <= rom_array(37210);
		when "1001000101011011" => data_out <= rom_array(37211);
		when "1001000101011100" => data_out <= rom_array(37212);
		when "1001000101011101" => data_out <= rom_array(37213);
		when "1001000101011110" => data_out <= rom_array(37214);
		when "1001000101011111" => data_out <= rom_array(37215);
		when "1001000101100000" => data_out <= rom_array(37216);
		when "1001000101100001" => data_out <= rom_array(37217);
		when "1001000101100010" => data_out <= rom_array(37218);
		when "1001000101100011" => data_out <= rom_array(37219);
		when "1001000101100100" => data_out <= rom_array(37220);
		when "1001000101100101" => data_out <= rom_array(37221);
		when "1001000101100110" => data_out <= rom_array(37222);
		when "1001000101100111" => data_out <= rom_array(37223);
		when "1001000101101000" => data_out <= rom_array(37224);
		when "1001000101101001" => data_out <= rom_array(37225);
		when "1001000101101010" => data_out <= rom_array(37226);
		when "1001000101101011" => data_out <= rom_array(37227);
		when "1001000101101100" => data_out <= rom_array(37228);
		when "1001000101101101" => data_out <= rom_array(37229);
		when "1001000101101110" => data_out <= rom_array(37230);
		when "1001000101101111" => data_out <= rom_array(37231);
		when "1001000101110000" => data_out <= rom_array(37232);
		when "1001000101110001" => data_out <= rom_array(37233);
		when "1001000101110010" => data_out <= rom_array(37234);
		when "1001000101110011" => data_out <= rom_array(37235);
		when "1001000101110100" => data_out <= rom_array(37236);
		when "1001000101110101" => data_out <= rom_array(37237);
		when "1001000101110110" => data_out <= rom_array(37238);
		when "1001000101110111" => data_out <= rom_array(37239);
		when "1001000101111000" => data_out <= rom_array(37240);
		when "1001000101111001" => data_out <= rom_array(37241);
		when "1001000101111010" => data_out <= rom_array(37242);
		when "1001000101111011" => data_out <= rom_array(37243);
		when "1001000101111100" => data_out <= rom_array(37244);
		when "1001000101111101" => data_out <= rom_array(37245);
		when "1001000101111110" => data_out <= rom_array(37246);
		when "1001000101111111" => data_out <= rom_array(37247);
		when "1001000110000000" => data_out <= rom_array(37248);
		when "1001000110000001" => data_out <= rom_array(37249);
		when "1001000110000010" => data_out <= rom_array(37250);
		when "1001000110000011" => data_out <= rom_array(37251);
		when "1001000110000100" => data_out <= rom_array(37252);
		when "1001000110000101" => data_out <= rom_array(37253);
		when "1001000110000110" => data_out <= rom_array(37254);
		when "1001000110000111" => data_out <= rom_array(37255);
		when "1001000110001000" => data_out <= rom_array(37256);
		when "1001000110001001" => data_out <= rom_array(37257);
		when "1001000110001010" => data_out <= rom_array(37258);
		when "1001000110001011" => data_out <= rom_array(37259);
		when "1001000110001100" => data_out <= rom_array(37260);
		when "1001000110001101" => data_out <= rom_array(37261);
		when "1001000110001110" => data_out <= rom_array(37262);
		when "1001000110001111" => data_out <= rom_array(37263);
		when "1001000110010000" => data_out <= rom_array(37264);
		when "1001000110010001" => data_out <= rom_array(37265);
		when "1001000110010010" => data_out <= rom_array(37266);
		when "1001000110010011" => data_out <= rom_array(37267);
		when "1001000110010100" => data_out <= rom_array(37268);
		when "1001000110010101" => data_out <= rom_array(37269);
		when "1001000110010110" => data_out <= rom_array(37270);
		when "1001000110010111" => data_out <= rom_array(37271);
		when "1001000110011000" => data_out <= rom_array(37272);
		when "1001000110011001" => data_out <= rom_array(37273);
		when "1001000110011010" => data_out <= rom_array(37274);
		when "1001000110011011" => data_out <= rom_array(37275);
		when "1001000110011100" => data_out <= rom_array(37276);
		when "1001000110011101" => data_out <= rom_array(37277);
		when "1001000110011110" => data_out <= rom_array(37278);
		when "1001000110011111" => data_out <= rom_array(37279);
		when "1001000110100000" => data_out <= rom_array(37280);
		when "1001000110100001" => data_out <= rom_array(37281);
		when "1001000110100010" => data_out <= rom_array(37282);
		when "1001000110100011" => data_out <= rom_array(37283);
		when "1001000110100100" => data_out <= rom_array(37284);
		when "1001000110100101" => data_out <= rom_array(37285);
		when "1001000110100110" => data_out <= rom_array(37286);
		when "1001000110100111" => data_out <= rom_array(37287);
		when "1001000110101000" => data_out <= rom_array(37288);
		when "1001000110101001" => data_out <= rom_array(37289);
		when "1001000110101010" => data_out <= rom_array(37290);
		when "1001000110101011" => data_out <= rom_array(37291);
		when "1001000110101100" => data_out <= rom_array(37292);
		when "1001000110101101" => data_out <= rom_array(37293);
		when "1001000110101110" => data_out <= rom_array(37294);
		when "1001000110101111" => data_out <= rom_array(37295);
		when "1001000110110000" => data_out <= rom_array(37296);
		when "1001000110110001" => data_out <= rom_array(37297);
		when "1001000110110010" => data_out <= rom_array(37298);
		when "1001000110110011" => data_out <= rom_array(37299);
		when "1001000110110100" => data_out <= rom_array(37300);
		when "1001000110110101" => data_out <= rom_array(37301);
		when "1001000110110110" => data_out <= rom_array(37302);
		when "1001000110110111" => data_out <= rom_array(37303);
		when "1001000110111000" => data_out <= rom_array(37304);
		when "1001000110111001" => data_out <= rom_array(37305);
		when "1001000110111010" => data_out <= rom_array(37306);
		when "1001000110111011" => data_out <= rom_array(37307);
		when "1001000110111100" => data_out <= rom_array(37308);
		when "1001000110111101" => data_out <= rom_array(37309);
		when "1001000110111110" => data_out <= rom_array(37310);
		when "1001000110111111" => data_out <= rom_array(37311);
		when "1001000111000000" => data_out <= rom_array(37312);
		when "1001000111000001" => data_out <= rom_array(37313);
		when "1001000111000010" => data_out <= rom_array(37314);
		when "1001000111000011" => data_out <= rom_array(37315);
		when "1001000111000100" => data_out <= rom_array(37316);
		when "1001000111000101" => data_out <= rom_array(37317);
		when "1001000111000110" => data_out <= rom_array(37318);
		when "1001000111000111" => data_out <= rom_array(37319);
		when "1001000111001000" => data_out <= rom_array(37320);
		when "1001000111001001" => data_out <= rom_array(37321);
		when "1001000111001010" => data_out <= rom_array(37322);
		when "1001000111001011" => data_out <= rom_array(37323);
		when "1001000111001100" => data_out <= rom_array(37324);
		when "1001000111001101" => data_out <= rom_array(37325);
		when "1001000111001110" => data_out <= rom_array(37326);
		when "1001000111001111" => data_out <= rom_array(37327);
		when "1001000111010000" => data_out <= rom_array(37328);
		when "1001000111010001" => data_out <= rom_array(37329);
		when "1001000111010010" => data_out <= rom_array(37330);
		when "1001000111010011" => data_out <= rom_array(37331);
		when "1001000111010100" => data_out <= rom_array(37332);
		when "1001000111010101" => data_out <= rom_array(37333);
		when "1001000111010110" => data_out <= rom_array(37334);
		when "1001000111010111" => data_out <= rom_array(37335);
		when "1001000111011000" => data_out <= rom_array(37336);
		when "1001000111011001" => data_out <= rom_array(37337);
		when "1001000111011010" => data_out <= rom_array(37338);
		when "1001000111011011" => data_out <= rom_array(37339);
		when "1001000111011100" => data_out <= rom_array(37340);
		when "1001000111011101" => data_out <= rom_array(37341);
		when "1001000111011110" => data_out <= rom_array(37342);
		when "1001000111011111" => data_out <= rom_array(37343);
		when "1001000111100000" => data_out <= rom_array(37344);
		when "1001000111100001" => data_out <= rom_array(37345);
		when "1001000111100010" => data_out <= rom_array(37346);
		when "1001000111100011" => data_out <= rom_array(37347);
		when "1001000111100100" => data_out <= rom_array(37348);
		when "1001000111100101" => data_out <= rom_array(37349);
		when "1001000111100110" => data_out <= rom_array(37350);
		when "1001000111100111" => data_out <= rom_array(37351);
		when "1001000111101000" => data_out <= rom_array(37352);
		when "1001000111101001" => data_out <= rom_array(37353);
		when "1001000111101010" => data_out <= rom_array(37354);
		when "1001000111101011" => data_out <= rom_array(37355);
		when "1001000111101100" => data_out <= rom_array(37356);
		when "1001000111101101" => data_out <= rom_array(37357);
		when "1001000111101110" => data_out <= rom_array(37358);
		when "1001000111101111" => data_out <= rom_array(37359);
		when "1001000111110000" => data_out <= rom_array(37360);
		when "1001000111110001" => data_out <= rom_array(37361);
		when "1001000111110010" => data_out <= rom_array(37362);
		when "1001000111110011" => data_out <= rom_array(37363);
		when "1001000111110100" => data_out <= rom_array(37364);
		when "1001000111110101" => data_out <= rom_array(37365);
		when "1001000111110110" => data_out <= rom_array(37366);
		when "1001000111110111" => data_out <= rom_array(37367);
		when "1001000111111000" => data_out <= rom_array(37368);
		when "1001000111111001" => data_out <= rom_array(37369);
		when "1001000111111010" => data_out <= rom_array(37370);
		when "1001000111111011" => data_out <= rom_array(37371);
		when "1001000111111100" => data_out <= rom_array(37372);
		when "1001000111111101" => data_out <= rom_array(37373);
		when "1001000111111110" => data_out <= rom_array(37374);
		when "1001000111111111" => data_out <= rom_array(37375);
		when "1001001000000000" => data_out <= rom_array(37376);
		when "1001001000000001" => data_out <= rom_array(37377);
		when "1001001000000010" => data_out <= rom_array(37378);
		when "1001001000000011" => data_out <= rom_array(37379);
		when "1001001000000100" => data_out <= rom_array(37380);
		when "1001001000000101" => data_out <= rom_array(37381);
		when "1001001000000110" => data_out <= rom_array(37382);
		when "1001001000000111" => data_out <= rom_array(37383);
		when "1001001000001000" => data_out <= rom_array(37384);
		when "1001001000001001" => data_out <= rom_array(37385);
		when "1001001000001010" => data_out <= rom_array(37386);
		when "1001001000001011" => data_out <= rom_array(37387);
		when "1001001000001100" => data_out <= rom_array(37388);
		when "1001001000001101" => data_out <= rom_array(37389);
		when "1001001000001110" => data_out <= rom_array(37390);
		when "1001001000001111" => data_out <= rom_array(37391);
		when "1001001000010000" => data_out <= rom_array(37392);
		when "1001001000010001" => data_out <= rom_array(37393);
		when "1001001000010010" => data_out <= rom_array(37394);
		when "1001001000010011" => data_out <= rom_array(37395);
		when "1001001000010100" => data_out <= rom_array(37396);
		when "1001001000010101" => data_out <= rom_array(37397);
		when "1001001000010110" => data_out <= rom_array(37398);
		when "1001001000010111" => data_out <= rom_array(37399);
		when "1001001000011000" => data_out <= rom_array(37400);
		when "1001001000011001" => data_out <= rom_array(37401);
		when "1001001000011010" => data_out <= rom_array(37402);
		when "1001001000011011" => data_out <= rom_array(37403);
		when "1001001000011100" => data_out <= rom_array(37404);
		when "1001001000011101" => data_out <= rom_array(37405);
		when "1001001000011110" => data_out <= rom_array(37406);
		when "1001001000011111" => data_out <= rom_array(37407);
		when "1001001000100000" => data_out <= rom_array(37408);
		when "1001001000100001" => data_out <= rom_array(37409);
		when "1001001000100010" => data_out <= rom_array(37410);
		when "1001001000100011" => data_out <= rom_array(37411);
		when "1001001000100100" => data_out <= rom_array(37412);
		when "1001001000100101" => data_out <= rom_array(37413);
		when "1001001000100110" => data_out <= rom_array(37414);
		when "1001001000100111" => data_out <= rom_array(37415);
		when "1001001000101000" => data_out <= rom_array(37416);
		when "1001001000101001" => data_out <= rom_array(37417);
		when "1001001000101010" => data_out <= rom_array(37418);
		when "1001001000101011" => data_out <= rom_array(37419);
		when "1001001000101100" => data_out <= rom_array(37420);
		when "1001001000101101" => data_out <= rom_array(37421);
		when "1001001000101110" => data_out <= rom_array(37422);
		when "1001001000101111" => data_out <= rom_array(37423);
		when "1001001000110000" => data_out <= rom_array(37424);
		when "1001001000110001" => data_out <= rom_array(37425);
		when "1001001000110010" => data_out <= rom_array(37426);
		when "1001001000110011" => data_out <= rom_array(37427);
		when "1001001000110100" => data_out <= rom_array(37428);
		when "1001001000110101" => data_out <= rom_array(37429);
		when "1001001000110110" => data_out <= rom_array(37430);
		when "1001001000110111" => data_out <= rom_array(37431);
		when "1001001000111000" => data_out <= rom_array(37432);
		when "1001001000111001" => data_out <= rom_array(37433);
		when "1001001000111010" => data_out <= rom_array(37434);
		when "1001001000111011" => data_out <= rom_array(37435);
		when "1001001000111100" => data_out <= rom_array(37436);
		when "1001001000111101" => data_out <= rom_array(37437);
		when "1001001000111110" => data_out <= rom_array(37438);
		when "1001001000111111" => data_out <= rom_array(37439);
		when "1001001001000000" => data_out <= rom_array(37440);
		when "1001001001000001" => data_out <= rom_array(37441);
		when "1001001001000010" => data_out <= rom_array(37442);
		when "1001001001000011" => data_out <= rom_array(37443);
		when "1001001001000100" => data_out <= rom_array(37444);
		when "1001001001000101" => data_out <= rom_array(37445);
		when "1001001001000110" => data_out <= rom_array(37446);
		when "1001001001000111" => data_out <= rom_array(37447);
		when "1001001001001000" => data_out <= rom_array(37448);
		when "1001001001001001" => data_out <= rom_array(37449);
		when "1001001001001010" => data_out <= rom_array(37450);
		when "1001001001001011" => data_out <= rom_array(37451);
		when "1001001001001100" => data_out <= rom_array(37452);
		when "1001001001001101" => data_out <= rom_array(37453);
		when "1001001001001110" => data_out <= rom_array(37454);
		when "1001001001001111" => data_out <= rom_array(37455);
		when "1001001001010000" => data_out <= rom_array(37456);
		when "1001001001010001" => data_out <= rom_array(37457);
		when "1001001001010010" => data_out <= rom_array(37458);
		when "1001001001010011" => data_out <= rom_array(37459);
		when "1001001001010100" => data_out <= rom_array(37460);
		when "1001001001010101" => data_out <= rom_array(37461);
		when "1001001001010110" => data_out <= rom_array(37462);
		when "1001001001010111" => data_out <= rom_array(37463);
		when "1001001001011000" => data_out <= rom_array(37464);
		when "1001001001011001" => data_out <= rom_array(37465);
		when "1001001001011010" => data_out <= rom_array(37466);
		when "1001001001011011" => data_out <= rom_array(37467);
		when "1001001001011100" => data_out <= rom_array(37468);
		when "1001001001011101" => data_out <= rom_array(37469);
		when "1001001001011110" => data_out <= rom_array(37470);
		when "1001001001011111" => data_out <= rom_array(37471);
		when "1001001001100000" => data_out <= rom_array(37472);
		when "1001001001100001" => data_out <= rom_array(37473);
		when "1001001001100010" => data_out <= rom_array(37474);
		when "1001001001100011" => data_out <= rom_array(37475);
		when "1001001001100100" => data_out <= rom_array(37476);
		when "1001001001100101" => data_out <= rom_array(37477);
		when "1001001001100110" => data_out <= rom_array(37478);
		when "1001001001100111" => data_out <= rom_array(37479);
		when "1001001001101000" => data_out <= rom_array(37480);
		when "1001001001101001" => data_out <= rom_array(37481);
		when "1001001001101010" => data_out <= rom_array(37482);
		when "1001001001101011" => data_out <= rom_array(37483);
		when "1001001001101100" => data_out <= rom_array(37484);
		when "1001001001101101" => data_out <= rom_array(37485);
		when "1001001001101110" => data_out <= rom_array(37486);
		when "1001001001101111" => data_out <= rom_array(37487);
		when "1001001001110000" => data_out <= rom_array(37488);
		when "1001001001110001" => data_out <= rom_array(37489);
		when "1001001001110010" => data_out <= rom_array(37490);
		when "1001001001110011" => data_out <= rom_array(37491);
		when "1001001001110100" => data_out <= rom_array(37492);
		when "1001001001110101" => data_out <= rom_array(37493);
		when "1001001001110110" => data_out <= rom_array(37494);
		when "1001001001110111" => data_out <= rom_array(37495);
		when "1001001001111000" => data_out <= rom_array(37496);
		when "1001001001111001" => data_out <= rom_array(37497);
		when "1001001001111010" => data_out <= rom_array(37498);
		when "1001001001111011" => data_out <= rom_array(37499);
		when "1001001001111100" => data_out <= rom_array(37500);
		when "1001001001111101" => data_out <= rom_array(37501);
		when "1001001001111110" => data_out <= rom_array(37502);
		when "1001001001111111" => data_out <= rom_array(37503);
		when "1001001010000000" => data_out <= rom_array(37504);
		when "1001001010000001" => data_out <= rom_array(37505);
		when "1001001010000010" => data_out <= rom_array(37506);
		when "1001001010000011" => data_out <= rom_array(37507);
		when "1001001010000100" => data_out <= rom_array(37508);
		when "1001001010000101" => data_out <= rom_array(37509);
		when "1001001010000110" => data_out <= rom_array(37510);
		when "1001001010000111" => data_out <= rom_array(37511);
		when "1001001010001000" => data_out <= rom_array(37512);
		when "1001001010001001" => data_out <= rom_array(37513);
		when "1001001010001010" => data_out <= rom_array(37514);
		when "1001001010001011" => data_out <= rom_array(37515);
		when "1001001010001100" => data_out <= rom_array(37516);
		when "1001001010001101" => data_out <= rom_array(37517);
		when "1001001010001110" => data_out <= rom_array(37518);
		when "1001001010001111" => data_out <= rom_array(37519);
		when "1001001010010000" => data_out <= rom_array(37520);
		when "1001001010010001" => data_out <= rom_array(37521);
		when "1001001010010010" => data_out <= rom_array(37522);
		when "1001001010010011" => data_out <= rom_array(37523);
		when "1001001010010100" => data_out <= rom_array(37524);
		when "1001001010010101" => data_out <= rom_array(37525);
		when "1001001010010110" => data_out <= rom_array(37526);
		when "1001001010010111" => data_out <= rom_array(37527);
		when "1001001010011000" => data_out <= rom_array(37528);
		when "1001001010011001" => data_out <= rom_array(37529);
		when "1001001010011010" => data_out <= rom_array(37530);
		when "1001001010011011" => data_out <= rom_array(37531);
		when "1001001010011100" => data_out <= rom_array(37532);
		when "1001001010011101" => data_out <= rom_array(37533);
		when "1001001010011110" => data_out <= rom_array(37534);
		when "1001001010011111" => data_out <= rom_array(37535);
		when "1001001010100000" => data_out <= rom_array(37536);
		when "1001001010100001" => data_out <= rom_array(37537);
		when "1001001010100010" => data_out <= rom_array(37538);
		when "1001001010100011" => data_out <= rom_array(37539);
		when "1001001010100100" => data_out <= rom_array(37540);
		when "1001001010100101" => data_out <= rom_array(37541);
		when "1001001010100110" => data_out <= rom_array(37542);
		when "1001001010100111" => data_out <= rom_array(37543);
		when "1001001010101000" => data_out <= rom_array(37544);
		when "1001001010101001" => data_out <= rom_array(37545);
		when "1001001010101010" => data_out <= rom_array(37546);
		when "1001001010101011" => data_out <= rom_array(37547);
		when "1001001010101100" => data_out <= rom_array(37548);
		when "1001001010101101" => data_out <= rom_array(37549);
		when "1001001010101110" => data_out <= rom_array(37550);
		when "1001001010101111" => data_out <= rom_array(37551);
		when "1001001010110000" => data_out <= rom_array(37552);
		when "1001001010110001" => data_out <= rom_array(37553);
		when "1001001010110010" => data_out <= rom_array(37554);
		when "1001001010110011" => data_out <= rom_array(37555);
		when "1001001010110100" => data_out <= rom_array(37556);
		when "1001001010110101" => data_out <= rom_array(37557);
		when "1001001010110110" => data_out <= rom_array(37558);
		when "1001001010110111" => data_out <= rom_array(37559);
		when "1001001010111000" => data_out <= rom_array(37560);
		when "1001001010111001" => data_out <= rom_array(37561);
		when "1001001010111010" => data_out <= rom_array(37562);
		when "1001001010111011" => data_out <= rom_array(37563);
		when "1001001010111100" => data_out <= rom_array(37564);
		when "1001001010111101" => data_out <= rom_array(37565);
		when "1001001010111110" => data_out <= rom_array(37566);
		when "1001001010111111" => data_out <= rom_array(37567);
		when "1001001011000000" => data_out <= rom_array(37568);
		when "1001001011000001" => data_out <= rom_array(37569);
		when "1001001011000010" => data_out <= rom_array(37570);
		when "1001001011000011" => data_out <= rom_array(37571);
		when "1001001011000100" => data_out <= rom_array(37572);
		when "1001001011000101" => data_out <= rom_array(37573);
		when "1001001011000110" => data_out <= rom_array(37574);
		when "1001001011000111" => data_out <= rom_array(37575);
		when "1001001011001000" => data_out <= rom_array(37576);
		when "1001001011001001" => data_out <= rom_array(37577);
		when "1001001011001010" => data_out <= rom_array(37578);
		when "1001001011001011" => data_out <= rom_array(37579);
		when "1001001011001100" => data_out <= rom_array(37580);
		when "1001001011001101" => data_out <= rom_array(37581);
		when "1001001011001110" => data_out <= rom_array(37582);
		when "1001001011001111" => data_out <= rom_array(37583);
		when "1001001011010000" => data_out <= rom_array(37584);
		when "1001001011010001" => data_out <= rom_array(37585);
		when "1001001011010010" => data_out <= rom_array(37586);
		when "1001001011010011" => data_out <= rom_array(37587);
		when "1001001011010100" => data_out <= rom_array(37588);
		when "1001001011010101" => data_out <= rom_array(37589);
		when "1001001011010110" => data_out <= rom_array(37590);
		when "1001001011010111" => data_out <= rom_array(37591);
		when "1001001011011000" => data_out <= rom_array(37592);
		when "1001001011011001" => data_out <= rom_array(37593);
		when "1001001011011010" => data_out <= rom_array(37594);
		when "1001001011011011" => data_out <= rom_array(37595);
		when "1001001011011100" => data_out <= rom_array(37596);
		when "1001001011011101" => data_out <= rom_array(37597);
		when "1001001011011110" => data_out <= rom_array(37598);
		when "1001001011011111" => data_out <= rom_array(37599);
		when "1001001011100000" => data_out <= rom_array(37600);
		when "1001001011100001" => data_out <= rom_array(37601);
		when "1001001011100010" => data_out <= rom_array(37602);
		when "1001001011100011" => data_out <= rom_array(37603);
		when "1001001011100100" => data_out <= rom_array(37604);
		when "1001001011100101" => data_out <= rom_array(37605);
		when "1001001011100110" => data_out <= rom_array(37606);
		when "1001001011100111" => data_out <= rom_array(37607);
		when "1001001011101000" => data_out <= rom_array(37608);
		when "1001001011101001" => data_out <= rom_array(37609);
		when "1001001011101010" => data_out <= rom_array(37610);
		when "1001001011101011" => data_out <= rom_array(37611);
		when "1001001011101100" => data_out <= rom_array(37612);
		when "1001001011101101" => data_out <= rom_array(37613);
		when "1001001011101110" => data_out <= rom_array(37614);
		when "1001001011101111" => data_out <= rom_array(37615);
		when "1001001011110000" => data_out <= rom_array(37616);
		when "1001001011110001" => data_out <= rom_array(37617);
		when "1001001011110010" => data_out <= rom_array(37618);
		when "1001001011110011" => data_out <= rom_array(37619);
		when "1001001011110100" => data_out <= rom_array(37620);
		when "1001001011110101" => data_out <= rom_array(37621);
		when "1001001011110110" => data_out <= rom_array(37622);
		when "1001001011110111" => data_out <= rom_array(37623);
		when "1001001011111000" => data_out <= rom_array(37624);
		when "1001001011111001" => data_out <= rom_array(37625);
		when "1001001011111010" => data_out <= rom_array(37626);
		when "1001001011111011" => data_out <= rom_array(37627);
		when "1001001011111100" => data_out <= rom_array(37628);
		when "1001001011111101" => data_out <= rom_array(37629);
		when "1001001011111110" => data_out <= rom_array(37630);
		when "1001001011111111" => data_out <= rom_array(37631);
		when "1001001100000000" => data_out <= rom_array(37632);
		when "1001001100000001" => data_out <= rom_array(37633);
		when "1001001100000010" => data_out <= rom_array(37634);
		when "1001001100000011" => data_out <= rom_array(37635);
		when "1001001100000100" => data_out <= rom_array(37636);
		when "1001001100000101" => data_out <= rom_array(37637);
		when "1001001100000110" => data_out <= rom_array(37638);
		when "1001001100000111" => data_out <= rom_array(37639);
		when "1001001100001000" => data_out <= rom_array(37640);
		when "1001001100001001" => data_out <= rom_array(37641);
		when "1001001100001010" => data_out <= rom_array(37642);
		when "1001001100001011" => data_out <= rom_array(37643);
		when "1001001100001100" => data_out <= rom_array(37644);
		when "1001001100001101" => data_out <= rom_array(37645);
		when "1001001100001110" => data_out <= rom_array(37646);
		when "1001001100001111" => data_out <= rom_array(37647);
		when "1001001100010000" => data_out <= rom_array(37648);
		when "1001001100010001" => data_out <= rom_array(37649);
		when "1001001100010010" => data_out <= rom_array(37650);
		when "1001001100010011" => data_out <= rom_array(37651);
		when "1001001100010100" => data_out <= rom_array(37652);
		when "1001001100010101" => data_out <= rom_array(37653);
		when "1001001100010110" => data_out <= rom_array(37654);
		when "1001001100010111" => data_out <= rom_array(37655);
		when "1001001100011000" => data_out <= rom_array(37656);
		when "1001001100011001" => data_out <= rom_array(37657);
		when "1001001100011010" => data_out <= rom_array(37658);
		when "1001001100011011" => data_out <= rom_array(37659);
		when "1001001100011100" => data_out <= rom_array(37660);
		when "1001001100011101" => data_out <= rom_array(37661);
		when "1001001100011110" => data_out <= rom_array(37662);
		when "1001001100011111" => data_out <= rom_array(37663);
		when "1001001100100000" => data_out <= rom_array(37664);
		when "1001001100100001" => data_out <= rom_array(37665);
		when "1001001100100010" => data_out <= rom_array(37666);
		when "1001001100100011" => data_out <= rom_array(37667);
		when "1001001100100100" => data_out <= rom_array(37668);
		when "1001001100100101" => data_out <= rom_array(37669);
		when "1001001100100110" => data_out <= rom_array(37670);
		when "1001001100100111" => data_out <= rom_array(37671);
		when "1001001100101000" => data_out <= rom_array(37672);
		when "1001001100101001" => data_out <= rom_array(37673);
		when "1001001100101010" => data_out <= rom_array(37674);
		when "1001001100101011" => data_out <= rom_array(37675);
		when "1001001100101100" => data_out <= rom_array(37676);
		when "1001001100101101" => data_out <= rom_array(37677);
		when "1001001100101110" => data_out <= rom_array(37678);
		when "1001001100101111" => data_out <= rom_array(37679);
		when "1001001100110000" => data_out <= rom_array(37680);
		when "1001001100110001" => data_out <= rom_array(37681);
		when "1001001100110010" => data_out <= rom_array(37682);
		when "1001001100110011" => data_out <= rom_array(37683);
		when "1001001100110100" => data_out <= rom_array(37684);
		when "1001001100110101" => data_out <= rom_array(37685);
		when "1001001100110110" => data_out <= rom_array(37686);
		when "1001001100110111" => data_out <= rom_array(37687);
		when "1001001100111000" => data_out <= rom_array(37688);
		when "1001001100111001" => data_out <= rom_array(37689);
		when "1001001100111010" => data_out <= rom_array(37690);
		when "1001001100111011" => data_out <= rom_array(37691);
		when "1001001100111100" => data_out <= rom_array(37692);
		when "1001001100111101" => data_out <= rom_array(37693);
		when "1001001100111110" => data_out <= rom_array(37694);
		when "1001001100111111" => data_out <= rom_array(37695);
		when "1001001101000000" => data_out <= rom_array(37696);
		when "1001001101000001" => data_out <= rom_array(37697);
		when "1001001101000010" => data_out <= rom_array(37698);
		when "1001001101000011" => data_out <= rom_array(37699);
		when "1001001101000100" => data_out <= rom_array(37700);
		when "1001001101000101" => data_out <= rom_array(37701);
		when "1001001101000110" => data_out <= rom_array(37702);
		when "1001001101000111" => data_out <= rom_array(37703);
		when "1001001101001000" => data_out <= rom_array(37704);
		when "1001001101001001" => data_out <= rom_array(37705);
		when "1001001101001010" => data_out <= rom_array(37706);
		when "1001001101001011" => data_out <= rom_array(37707);
		when "1001001101001100" => data_out <= rom_array(37708);
		when "1001001101001101" => data_out <= rom_array(37709);
		when "1001001101001110" => data_out <= rom_array(37710);
		when "1001001101001111" => data_out <= rom_array(37711);
		when "1001001101010000" => data_out <= rom_array(37712);
		when "1001001101010001" => data_out <= rom_array(37713);
		when "1001001101010010" => data_out <= rom_array(37714);
		when "1001001101010011" => data_out <= rom_array(37715);
		when "1001001101010100" => data_out <= rom_array(37716);
		when "1001001101010101" => data_out <= rom_array(37717);
		when "1001001101010110" => data_out <= rom_array(37718);
		when "1001001101010111" => data_out <= rom_array(37719);
		when "1001001101011000" => data_out <= rom_array(37720);
		when "1001001101011001" => data_out <= rom_array(37721);
		when "1001001101011010" => data_out <= rom_array(37722);
		when "1001001101011011" => data_out <= rom_array(37723);
		when "1001001101011100" => data_out <= rom_array(37724);
		when "1001001101011101" => data_out <= rom_array(37725);
		when "1001001101011110" => data_out <= rom_array(37726);
		when "1001001101011111" => data_out <= rom_array(37727);
		when "1001001101100000" => data_out <= rom_array(37728);
		when "1001001101100001" => data_out <= rom_array(37729);
		when "1001001101100010" => data_out <= rom_array(37730);
		when "1001001101100011" => data_out <= rom_array(37731);
		when "1001001101100100" => data_out <= rom_array(37732);
		when "1001001101100101" => data_out <= rom_array(37733);
		when "1001001101100110" => data_out <= rom_array(37734);
		when "1001001101100111" => data_out <= rom_array(37735);
		when "1001001101101000" => data_out <= rom_array(37736);
		when "1001001101101001" => data_out <= rom_array(37737);
		when "1001001101101010" => data_out <= rom_array(37738);
		when "1001001101101011" => data_out <= rom_array(37739);
		when "1001001101101100" => data_out <= rom_array(37740);
		when "1001001101101101" => data_out <= rom_array(37741);
		when "1001001101101110" => data_out <= rom_array(37742);
		when "1001001101101111" => data_out <= rom_array(37743);
		when "1001001101110000" => data_out <= rom_array(37744);
		when "1001001101110001" => data_out <= rom_array(37745);
		when "1001001101110010" => data_out <= rom_array(37746);
		when "1001001101110011" => data_out <= rom_array(37747);
		when "1001001101110100" => data_out <= rom_array(37748);
		when "1001001101110101" => data_out <= rom_array(37749);
		when "1001001101110110" => data_out <= rom_array(37750);
		when "1001001101110111" => data_out <= rom_array(37751);
		when "1001001101111000" => data_out <= rom_array(37752);
		when "1001001101111001" => data_out <= rom_array(37753);
		when "1001001101111010" => data_out <= rom_array(37754);
		when "1001001101111011" => data_out <= rom_array(37755);
		when "1001001101111100" => data_out <= rom_array(37756);
		when "1001001101111101" => data_out <= rom_array(37757);
		when "1001001101111110" => data_out <= rom_array(37758);
		when "1001001101111111" => data_out <= rom_array(37759);
		when "1001001110000000" => data_out <= rom_array(37760);
		when "1001001110000001" => data_out <= rom_array(37761);
		when "1001001110000010" => data_out <= rom_array(37762);
		when "1001001110000011" => data_out <= rom_array(37763);
		when "1001001110000100" => data_out <= rom_array(37764);
		when "1001001110000101" => data_out <= rom_array(37765);
		when "1001001110000110" => data_out <= rom_array(37766);
		when "1001001110000111" => data_out <= rom_array(37767);
		when "1001001110001000" => data_out <= rom_array(37768);
		when "1001001110001001" => data_out <= rom_array(37769);
		when "1001001110001010" => data_out <= rom_array(37770);
		when "1001001110001011" => data_out <= rom_array(37771);
		when "1001001110001100" => data_out <= rom_array(37772);
		when "1001001110001101" => data_out <= rom_array(37773);
		when "1001001110001110" => data_out <= rom_array(37774);
		when "1001001110001111" => data_out <= rom_array(37775);
		when "1001001110010000" => data_out <= rom_array(37776);
		when "1001001110010001" => data_out <= rom_array(37777);
		when "1001001110010010" => data_out <= rom_array(37778);
		when "1001001110010011" => data_out <= rom_array(37779);
		when "1001001110010100" => data_out <= rom_array(37780);
		when "1001001110010101" => data_out <= rom_array(37781);
		when "1001001110010110" => data_out <= rom_array(37782);
		when "1001001110010111" => data_out <= rom_array(37783);
		when "1001001110011000" => data_out <= rom_array(37784);
		when "1001001110011001" => data_out <= rom_array(37785);
		when "1001001110011010" => data_out <= rom_array(37786);
		when "1001001110011011" => data_out <= rom_array(37787);
		when "1001001110011100" => data_out <= rom_array(37788);
		when "1001001110011101" => data_out <= rom_array(37789);
		when "1001001110011110" => data_out <= rom_array(37790);
		when "1001001110011111" => data_out <= rom_array(37791);
		when "1001001110100000" => data_out <= rom_array(37792);
		when "1001001110100001" => data_out <= rom_array(37793);
		when "1001001110100010" => data_out <= rom_array(37794);
		when "1001001110100011" => data_out <= rom_array(37795);
		when "1001001110100100" => data_out <= rom_array(37796);
		when "1001001110100101" => data_out <= rom_array(37797);
		when "1001001110100110" => data_out <= rom_array(37798);
		when "1001001110100111" => data_out <= rom_array(37799);
		when "1001001110101000" => data_out <= rom_array(37800);
		when "1001001110101001" => data_out <= rom_array(37801);
		when "1001001110101010" => data_out <= rom_array(37802);
		when "1001001110101011" => data_out <= rom_array(37803);
		when "1001001110101100" => data_out <= rom_array(37804);
		when "1001001110101101" => data_out <= rom_array(37805);
		when "1001001110101110" => data_out <= rom_array(37806);
		when "1001001110101111" => data_out <= rom_array(37807);
		when "1001001110110000" => data_out <= rom_array(37808);
		when "1001001110110001" => data_out <= rom_array(37809);
		when "1001001110110010" => data_out <= rom_array(37810);
		when "1001001110110011" => data_out <= rom_array(37811);
		when "1001001110110100" => data_out <= rom_array(37812);
		when "1001001110110101" => data_out <= rom_array(37813);
		when "1001001110110110" => data_out <= rom_array(37814);
		when "1001001110110111" => data_out <= rom_array(37815);
		when "1001001110111000" => data_out <= rom_array(37816);
		when "1001001110111001" => data_out <= rom_array(37817);
		when "1001001110111010" => data_out <= rom_array(37818);
		when "1001001110111011" => data_out <= rom_array(37819);
		when "1001001110111100" => data_out <= rom_array(37820);
		when "1001001110111101" => data_out <= rom_array(37821);
		when "1001001110111110" => data_out <= rom_array(37822);
		when "1001001110111111" => data_out <= rom_array(37823);
		when "1001001111000000" => data_out <= rom_array(37824);
		when "1001001111000001" => data_out <= rom_array(37825);
		when "1001001111000010" => data_out <= rom_array(37826);
		when "1001001111000011" => data_out <= rom_array(37827);
		when "1001001111000100" => data_out <= rom_array(37828);
		when "1001001111000101" => data_out <= rom_array(37829);
		when "1001001111000110" => data_out <= rom_array(37830);
		when "1001001111000111" => data_out <= rom_array(37831);
		when "1001001111001000" => data_out <= rom_array(37832);
		when "1001001111001001" => data_out <= rom_array(37833);
		when "1001001111001010" => data_out <= rom_array(37834);
		when "1001001111001011" => data_out <= rom_array(37835);
		when "1001001111001100" => data_out <= rom_array(37836);
		when "1001001111001101" => data_out <= rom_array(37837);
		when "1001001111001110" => data_out <= rom_array(37838);
		when "1001001111001111" => data_out <= rom_array(37839);
		when "1001001111010000" => data_out <= rom_array(37840);
		when "1001001111010001" => data_out <= rom_array(37841);
		when "1001001111010010" => data_out <= rom_array(37842);
		when "1001001111010011" => data_out <= rom_array(37843);
		when "1001001111010100" => data_out <= rom_array(37844);
		when "1001001111010101" => data_out <= rom_array(37845);
		when "1001001111010110" => data_out <= rom_array(37846);
		when "1001001111010111" => data_out <= rom_array(37847);
		when "1001001111011000" => data_out <= rom_array(37848);
		when "1001001111011001" => data_out <= rom_array(37849);
		when "1001001111011010" => data_out <= rom_array(37850);
		when "1001001111011011" => data_out <= rom_array(37851);
		when "1001001111011100" => data_out <= rom_array(37852);
		when "1001001111011101" => data_out <= rom_array(37853);
		when "1001001111011110" => data_out <= rom_array(37854);
		when "1001001111011111" => data_out <= rom_array(37855);
		when "1001001111100000" => data_out <= rom_array(37856);
		when "1001001111100001" => data_out <= rom_array(37857);
		when "1001001111100010" => data_out <= rom_array(37858);
		when "1001001111100011" => data_out <= rom_array(37859);
		when "1001001111100100" => data_out <= rom_array(37860);
		when "1001001111100101" => data_out <= rom_array(37861);
		when "1001001111100110" => data_out <= rom_array(37862);
		when "1001001111100111" => data_out <= rom_array(37863);
		when "1001001111101000" => data_out <= rom_array(37864);
		when "1001001111101001" => data_out <= rom_array(37865);
		when "1001001111101010" => data_out <= rom_array(37866);
		when "1001001111101011" => data_out <= rom_array(37867);
		when "1001001111101100" => data_out <= rom_array(37868);
		when "1001001111101101" => data_out <= rom_array(37869);
		when "1001001111101110" => data_out <= rom_array(37870);
		when "1001001111101111" => data_out <= rom_array(37871);
		when "1001001111110000" => data_out <= rom_array(37872);
		when "1001001111110001" => data_out <= rom_array(37873);
		when "1001001111110010" => data_out <= rom_array(37874);
		when "1001001111110011" => data_out <= rom_array(37875);
		when "1001001111110100" => data_out <= rom_array(37876);
		when "1001001111110101" => data_out <= rom_array(37877);
		when "1001001111110110" => data_out <= rom_array(37878);
		when "1001001111110111" => data_out <= rom_array(37879);
		when "1001001111111000" => data_out <= rom_array(37880);
		when "1001001111111001" => data_out <= rom_array(37881);
		when "1001001111111010" => data_out <= rom_array(37882);
		when "1001001111111011" => data_out <= rom_array(37883);
		when "1001001111111100" => data_out <= rom_array(37884);
		when "1001001111111101" => data_out <= rom_array(37885);
		when "1001001111111110" => data_out <= rom_array(37886);
		when "1001001111111111" => data_out <= rom_array(37887);
		when "1001010000000000" => data_out <= rom_array(37888);
		when "1001010000000001" => data_out <= rom_array(37889);
		when "1001010000000010" => data_out <= rom_array(37890);
		when "1001010000000011" => data_out <= rom_array(37891);
		when "1001010000000100" => data_out <= rom_array(37892);
		when "1001010000000101" => data_out <= rom_array(37893);
		when "1001010000000110" => data_out <= rom_array(37894);
		when "1001010000000111" => data_out <= rom_array(37895);
		when "1001010000001000" => data_out <= rom_array(37896);
		when "1001010000001001" => data_out <= rom_array(37897);
		when "1001010000001010" => data_out <= rom_array(37898);
		when "1001010000001011" => data_out <= rom_array(37899);
		when "1001010000001100" => data_out <= rom_array(37900);
		when "1001010000001101" => data_out <= rom_array(37901);
		when "1001010000001110" => data_out <= rom_array(37902);
		when "1001010000001111" => data_out <= rom_array(37903);
		when "1001010000010000" => data_out <= rom_array(37904);
		when "1001010000010001" => data_out <= rom_array(37905);
		when "1001010000010010" => data_out <= rom_array(37906);
		when "1001010000010011" => data_out <= rom_array(37907);
		when "1001010000010100" => data_out <= rom_array(37908);
		when "1001010000010101" => data_out <= rom_array(37909);
		when "1001010000010110" => data_out <= rom_array(37910);
		when "1001010000010111" => data_out <= rom_array(37911);
		when "1001010000011000" => data_out <= rom_array(37912);
		when "1001010000011001" => data_out <= rom_array(37913);
		when "1001010000011010" => data_out <= rom_array(37914);
		when "1001010000011011" => data_out <= rom_array(37915);
		when "1001010000011100" => data_out <= rom_array(37916);
		when "1001010000011101" => data_out <= rom_array(37917);
		when "1001010000011110" => data_out <= rom_array(37918);
		when "1001010000011111" => data_out <= rom_array(37919);
		when "1001010000100000" => data_out <= rom_array(37920);
		when "1001010000100001" => data_out <= rom_array(37921);
		when "1001010000100010" => data_out <= rom_array(37922);
		when "1001010000100011" => data_out <= rom_array(37923);
		when "1001010000100100" => data_out <= rom_array(37924);
		when "1001010000100101" => data_out <= rom_array(37925);
		when "1001010000100110" => data_out <= rom_array(37926);
		when "1001010000100111" => data_out <= rom_array(37927);
		when "1001010000101000" => data_out <= rom_array(37928);
		when "1001010000101001" => data_out <= rom_array(37929);
		when "1001010000101010" => data_out <= rom_array(37930);
		when "1001010000101011" => data_out <= rom_array(37931);
		when "1001010000101100" => data_out <= rom_array(37932);
		when "1001010000101101" => data_out <= rom_array(37933);
		when "1001010000101110" => data_out <= rom_array(37934);
		when "1001010000101111" => data_out <= rom_array(37935);
		when "1001010000110000" => data_out <= rom_array(37936);
		when "1001010000110001" => data_out <= rom_array(37937);
		when "1001010000110010" => data_out <= rom_array(37938);
		when "1001010000110011" => data_out <= rom_array(37939);
		when "1001010000110100" => data_out <= rom_array(37940);
		when "1001010000110101" => data_out <= rom_array(37941);
		when "1001010000110110" => data_out <= rom_array(37942);
		when "1001010000110111" => data_out <= rom_array(37943);
		when "1001010000111000" => data_out <= rom_array(37944);
		when "1001010000111001" => data_out <= rom_array(37945);
		when "1001010000111010" => data_out <= rom_array(37946);
		when "1001010000111011" => data_out <= rom_array(37947);
		when "1001010000111100" => data_out <= rom_array(37948);
		when "1001010000111101" => data_out <= rom_array(37949);
		when "1001010000111110" => data_out <= rom_array(37950);
		when "1001010000111111" => data_out <= rom_array(37951);
		when "1001010001000000" => data_out <= rom_array(37952);
		when "1001010001000001" => data_out <= rom_array(37953);
		when "1001010001000010" => data_out <= rom_array(37954);
		when "1001010001000011" => data_out <= rom_array(37955);
		when "1001010001000100" => data_out <= rom_array(37956);
		when "1001010001000101" => data_out <= rom_array(37957);
		when "1001010001000110" => data_out <= rom_array(37958);
		when "1001010001000111" => data_out <= rom_array(37959);
		when "1001010001001000" => data_out <= rom_array(37960);
		when "1001010001001001" => data_out <= rom_array(37961);
		when "1001010001001010" => data_out <= rom_array(37962);
		when "1001010001001011" => data_out <= rom_array(37963);
		when "1001010001001100" => data_out <= rom_array(37964);
		when "1001010001001101" => data_out <= rom_array(37965);
		when "1001010001001110" => data_out <= rom_array(37966);
		when "1001010001001111" => data_out <= rom_array(37967);
		when "1001010001010000" => data_out <= rom_array(37968);
		when "1001010001010001" => data_out <= rom_array(37969);
		when "1001010001010010" => data_out <= rom_array(37970);
		when "1001010001010011" => data_out <= rom_array(37971);
		when "1001010001010100" => data_out <= rom_array(37972);
		when "1001010001010101" => data_out <= rom_array(37973);
		when "1001010001010110" => data_out <= rom_array(37974);
		when "1001010001010111" => data_out <= rom_array(37975);
		when "1001010001011000" => data_out <= rom_array(37976);
		when "1001010001011001" => data_out <= rom_array(37977);
		when "1001010001011010" => data_out <= rom_array(37978);
		when "1001010001011011" => data_out <= rom_array(37979);
		when "1001010001011100" => data_out <= rom_array(37980);
		when "1001010001011101" => data_out <= rom_array(37981);
		when "1001010001011110" => data_out <= rom_array(37982);
		when "1001010001011111" => data_out <= rom_array(37983);
		when "1001010001100000" => data_out <= rom_array(37984);
		when "1001010001100001" => data_out <= rom_array(37985);
		when "1001010001100010" => data_out <= rom_array(37986);
		when "1001010001100011" => data_out <= rom_array(37987);
		when "1001010001100100" => data_out <= rom_array(37988);
		when "1001010001100101" => data_out <= rom_array(37989);
		when "1001010001100110" => data_out <= rom_array(37990);
		when "1001010001100111" => data_out <= rom_array(37991);
		when "1001010001101000" => data_out <= rom_array(37992);
		when "1001010001101001" => data_out <= rom_array(37993);
		when "1001010001101010" => data_out <= rom_array(37994);
		when "1001010001101011" => data_out <= rom_array(37995);
		when "1001010001101100" => data_out <= rom_array(37996);
		when "1001010001101101" => data_out <= rom_array(37997);
		when "1001010001101110" => data_out <= rom_array(37998);
		when "1001010001101111" => data_out <= rom_array(37999);
		when "1001010001110000" => data_out <= rom_array(38000);
		when "1001010001110001" => data_out <= rom_array(38001);
		when "1001010001110010" => data_out <= rom_array(38002);
		when "1001010001110011" => data_out <= rom_array(38003);
		when "1001010001110100" => data_out <= rom_array(38004);
		when "1001010001110101" => data_out <= rom_array(38005);
		when "1001010001110110" => data_out <= rom_array(38006);
		when "1001010001110111" => data_out <= rom_array(38007);
		when "1001010001111000" => data_out <= rom_array(38008);
		when "1001010001111001" => data_out <= rom_array(38009);
		when "1001010001111010" => data_out <= rom_array(38010);
		when "1001010001111011" => data_out <= rom_array(38011);
		when "1001010001111100" => data_out <= rom_array(38012);
		when "1001010001111101" => data_out <= rom_array(38013);
		when "1001010001111110" => data_out <= rom_array(38014);
		when "1001010001111111" => data_out <= rom_array(38015);
		when "1001010010000000" => data_out <= rom_array(38016);
		when "1001010010000001" => data_out <= rom_array(38017);
		when "1001010010000010" => data_out <= rom_array(38018);
		when "1001010010000011" => data_out <= rom_array(38019);
		when "1001010010000100" => data_out <= rom_array(38020);
		when "1001010010000101" => data_out <= rom_array(38021);
		when "1001010010000110" => data_out <= rom_array(38022);
		when "1001010010000111" => data_out <= rom_array(38023);
		when "1001010010001000" => data_out <= rom_array(38024);
		when "1001010010001001" => data_out <= rom_array(38025);
		when "1001010010001010" => data_out <= rom_array(38026);
		when "1001010010001011" => data_out <= rom_array(38027);
		when "1001010010001100" => data_out <= rom_array(38028);
		when "1001010010001101" => data_out <= rom_array(38029);
		when "1001010010001110" => data_out <= rom_array(38030);
		when "1001010010001111" => data_out <= rom_array(38031);
		when "1001010010010000" => data_out <= rom_array(38032);
		when "1001010010010001" => data_out <= rom_array(38033);
		when "1001010010010010" => data_out <= rom_array(38034);
		when "1001010010010011" => data_out <= rom_array(38035);
		when "1001010010010100" => data_out <= rom_array(38036);
		when "1001010010010101" => data_out <= rom_array(38037);
		when "1001010010010110" => data_out <= rom_array(38038);
		when "1001010010010111" => data_out <= rom_array(38039);
		when "1001010010011000" => data_out <= rom_array(38040);
		when "1001010010011001" => data_out <= rom_array(38041);
		when "1001010010011010" => data_out <= rom_array(38042);
		when "1001010010011011" => data_out <= rom_array(38043);
		when "1001010010011100" => data_out <= rom_array(38044);
		when "1001010010011101" => data_out <= rom_array(38045);
		when "1001010010011110" => data_out <= rom_array(38046);
		when "1001010010011111" => data_out <= rom_array(38047);
		when "1001010010100000" => data_out <= rom_array(38048);
		when "1001010010100001" => data_out <= rom_array(38049);
		when "1001010010100010" => data_out <= rom_array(38050);
		when "1001010010100011" => data_out <= rom_array(38051);
		when "1001010010100100" => data_out <= rom_array(38052);
		when "1001010010100101" => data_out <= rom_array(38053);
		when "1001010010100110" => data_out <= rom_array(38054);
		when "1001010010100111" => data_out <= rom_array(38055);
		when "1001010010101000" => data_out <= rom_array(38056);
		when "1001010010101001" => data_out <= rom_array(38057);
		when "1001010010101010" => data_out <= rom_array(38058);
		when "1001010010101011" => data_out <= rom_array(38059);
		when "1001010010101100" => data_out <= rom_array(38060);
		when "1001010010101101" => data_out <= rom_array(38061);
		when "1001010010101110" => data_out <= rom_array(38062);
		when "1001010010101111" => data_out <= rom_array(38063);
		when "1001010010110000" => data_out <= rom_array(38064);
		when "1001010010110001" => data_out <= rom_array(38065);
		when "1001010010110010" => data_out <= rom_array(38066);
		when "1001010010110011" => data_out <= rom_array(38067);
		when "1001010010110100" => data_out <= rom_array(38068);
		when "1001010010110101" => data_out <= rom_array(38069);
		when "1001010010110110" => data_out <= rom_array(38070);
		when "1001010010110111" => data_out <= rom_array(38071);
		when "1001010010111000" => data_out <= rom_array(38072);
		when "1001010010111001" => data_out <= rom_array(38073);
		when "1001010010111010" => data_out <= rom_array(38074);
		when "1001010010111011" => data_out <= rom_array(38075);
		when "1001010010111100" => data_out <= rom_array(38076);
		when "1001010010111101" => data_out <= rom_array(38077);
		when "1001010010111110" => data_out <= rom_array(38078);
		when "1001010010111111" => data_out <= rom_array(38079);
		when "1001010011000000" => data_out <= rom_array(38080);
		when "1001010011000001" => data_out <= rom_array(38081);
		when "1001010011000010" => data_out <= rom_array(38082);
		when "1001010011000011" => data_out <= rom_array(38083);
		when "1001010011000100" => data_out <= rom_array(38084);
		when "1001010011000101" => data_out <= rom_array(38085);
		when "1001010011000110" => data_out <= rom_array(38086);
		when "1001010011000111" => data_out <= rom_array(38087);
		when "1001010011001000" => data_out <= rom_array(38088);
		when "1001010011001001" => data_out <= rom_array(38089);
		when "1001010011001010" => data_out <= rom_array(38090);
		when "1001010011001011" => data_out <= rom_array(38091);
		when "1001010011001100" => data_out <= rom_array(38092);
		when "1001010011001101" => data_out <= rom_array(38093);
		when "1001010011001110" => data_out <= rom_array(38094);
		when "1001010011001111" => data_out <= rom_array(38095);
		when "1001010011010000" => data_out <= rom_array(38096);
		when "1001010011010001" => data_out <= rom_array(38097);
		when "1001010011010010" => data_out <= rom_array(38098);
		when "1001010011010011" => data_out <= rom_array(38099);
		when "1001010011010100" => data_out <= rom_array(38100);
		when "1001010011010101" => data_out <= rom_array(38101);
		when "1001010011010110" => data_out <= rom_array(38102);
		when "1001010011010111" => data_out <= rom_array(38103);
		when "1001010011011000" => data_out <= rom_array(38104);
		when "1001010011011001" => data_out <= rom_array(38105);
		when "1001010011011010" => data_out <= rom_array(38106);
		when "1001010011011011" => data_out <= rom_array(38107);
		when "1001010011011100" => data_out <= rom_array(38108);
		when "1001010011011101" => data_out <= rom_array(38109);
		when "1001010011011110" => data_out <= rom_array(38110);
		when "1001010011011111" => data_out <= rom_array(38111);
		when "1001010011100000" => data_out <= rom_array(38112);
		when "1001010011100001" => data_out <= rom_array(38113);
		when "1001010011100010" => data_out <= rom_array(38114);
		when "1001010011100011" => data_out <= rom_array(38115);
		when "1001010011100100" => data_out <= rom_array(38116);
		when "1001010011100101" => data_out <= rom_array(38117);
		when "1001010011100110" => data_out <= rom_array(38118);
		when "1001010011100111" => data_out <= rom_array(38119);
		when "1001010011101000" => data_out <= rom_array(38120);
		when "1001010011101001" => data_out <= rom_array(38121);
		when "1001010011101010" => data_out <= rom_array(38122);
		when "1001010011101011" => data_out <= rom_array(38123);
		when "1001010011101100" => data_out <= rom_array(38124);
		when "1001010011101101" => data_out <= rom_array(38125);
		when "1001010011101110" => data_out <= rom_array(38126);
		when "1001010011101111" => data_out <= rom_array(38127);
		when "1001010011110000" => data_out <= rom_array(38128);
		when "1001010011110001" => data_out <= rom_array(38129);
		when "1001010011110010" => data_out <= rom_array(38130);
		when "1001010011110011" => data_out <= rom_array(38131);
		when "1001010011110100" => data_out <= rom_array(38132);
		when "1001010011110101" => data_out <= rom_array(38133);
		when "1001010011110110" => data_out <= rom_array(38134);
		when "1001010011110111" => data_out <= rom_array(38135);
		when "1001010011111000" => data_out <= rom_array(38136);
		when "1001010011111001" => data_out <= rom_array(38137);
		when "1001010011111010" => data_out <= rom_array(38138);
		when "1001010011111011" => data_out <= rom_array(38139);
		when "1001010011111100" => data_out <= rom_array(38140);
		when "1001010011111101" => data_out <= rom_array(38141);
		when "1001010011111110" => data_out <= rom_array(38142);
		when "1001010011111111" => data_out <= rom_array(38143);
		when "1001010100000000" => data_out <= rom_array(38144);
		when "1001010100000001" => data_out <= rom_array(38145);
		when "1001010100000010" => data_out <= rom_array(38146);
		when "1001010100000011" => data_out <= rom_array(38147);
		when "1001010100000100" => data_out <= rom_array(38148);
		when "1001010100000101" => data_out <= rom_array(38149);
		when "1001010100000110" => data_out <= rom_array(38150);
		when "1001010100000111" => data_out <= rom_array(38151);
		when "1001010100001000" => data_out <= rom_array(38152);
		when "1001010100001001" => data_out <= rom_array(38153);
		when "1001010100001010" => data_out <= rom_array(38154);
		when "1001010100001011" => data_out <= rom_array(38155);
		when "1001010100001100" => data_out <= rom_array(38156);
		when "1001010100001101" => data_out <= rom_array(38157);
		when "1001010100001110" => data_out <= rom_array(38158);
		when "1001010100001111" => data_out <= rom_array(38159);
		when "1001010100010000" => data_out <= rom_array(38160);
		when "1001010100010001" => data_out <= rom_array(38161);
		when "1001010100010010" => data_out <= rom_array(38162);
		when "1001010100010011" => data_out <= rom_array(38163);
		when "1001010100010100" => data_out <= rom_array(38164);
		when "1001010100010101" => data_out <= rom_array(38165);
		when "1001010100010110" => data_out <= rom_array(38166);
		when "1001010100010111" => data_out <= rom_array(38167);
		when "1001010100011000" => data_out <= rom_array(38168);
		when "1001010100011001" => data_out <= rom_array(38169);
		when "1001010100011010" => data_out <= rom_array(38170);
		when "1001010100011011" => data_out <= rom_array(38171);
		when "1001010100011100" => data_out <= rom_array(38172);
		when "1001010100011101" => data_out <= rom_array(38173);
		when "1001010100011110" => data_out <= rom_array(38174);
		when "1001010100011111" => data_out <= rom_array(38175);
		when "1001010100100000" => data_out <= rom_array(38176);
		when "1001010100100001" => data_out <= rom_array(38177);
		when "1001010100100010" => data_out <= rom_array(38178);
		when "1001010100100011" => data_out <= rom_array(38179);
		when "1001010100100100" => data_out <= rom_array(38180);
		when "1001010100100101" => data_out <= rom_array(38181);
		when "1001010100100110" => data_out <= rom_array(38182);
		when "1001010100100111" => data_out <= rom_array(38183);
		when "1001010100101000" => data_out <= rom_array(38184);
		when "1001010100101001" => data_out <= rom_array(38185);
		when "1001010100101010" => data_out <= rom_array(38186);
		when "1001010100101011" => data_out <= rom_array(38187);
		when "1001010100101100" => data_out <= rom_array(38188);
		when "1001010100101101" => data_out <= rom_array(38189);
		when "1001010100101110" => data_out <= rom_array(38190);
		when "1001010100101111" => data_out <= rom_array(38191);
		when "1001010100110000" => data_out <= rom_array(38192);
		when "1001010100110001" => data_out <= rom_array(38193);
		when "1001010100110010" => data_out <= rom_array(38194);
		when "1001010100110011" => data_out <= rom_array(38195);
		when "1001010100110100" => data_out <= rom_array(38196);
		when "1001010100110101" => data_out <= rom_array(38197);
		when "1001010100110110" => data_out <= rom_array(38198);
		when "1001010100110111" => data_out <= rom_array(38199);
		when "1001010100111000" => data_out <= rom_array(38200);
		when "1001010100111001" => data_out <= rom_array(38201);
		when "1001010100111010" => data_out <= rom_array(38202);
		when "1001010100111011" => data_out <= rom_array(38203);
		when "1001010100111100" => data_out <= rom_array(38204);
		when "1001010100111101" => data_out <= rom_array(38205);
		when "1001010100111110" => data_out <= rom_array(38206);
		when "1001010100111111" => data_out <= rom_array(38207);
		when "1001010101000000" => data_out <= rom_array(38208);
		when "1001010101000001" => data_out <= rom_array(38209);
		when "1001010101000010" => data_out <= rom_array(38210);
		when "1001010101000011" => data_out <= rom_array(38211);
		when "1001010101000100" => data_out <= rom_array(38212);
		when "1001010101000101" => data_out <= rom_array(38213);
		when "1001010101000110" => data_out <= rom_array(38214);
		when "1001010101000111" => data_out <= rom_array(38215);
		when "1001010101001000" => data_out <= rom_array(38216);
		when "1001010101001001" => data_out <= rom_array(38217);
		when "1001010101001010" => data_out <= rom_array(38218);
		when "1001010101001011" => data_out <= rom_array(38219);
		when "1001010101001100" => data_out <= rom_array(38220);
		when "1001010101001101" => data_out <= rom_array(38221);
		when "1001010101001110" => data_out <= rom_array(38222);
		when "1001010101001111" => data_out <= rom_array(38223);
		when "1001010101010000" => data_out <= rom_array(38224);
		when "1001010101010001" => data_out <= rom_array(38225);
		when "1001010101010010" => data_out <= rom_array(38226);
		when "1001010101010011" => data_out <= rom_array(38227);
		when "1001010101010100" => data_out <= rom_array(38228);
		when "1001010101010101" => data_out <= rom_array(38229);
		when "1001010101010110" => data_out <= rom_array(38230);
		when "1001010101010111" => data_out <= rom_array(38231);
		when "1001010101011000" => data_out <= rom_array(38232);
		when "1001010101011001" => data_out <= rom_array(38233);
		when "1001010101011010" => data_out <= rom_array(38234);
		when "1001010101011011" => data_out <= rom_array(38235);
		when "1001010101011100" => data_out <= rom_array(38236);
		when "1001010101011101" => data_out <= rom_array(38237);
		when "1001010101011110" => data_out <= rom_array(38238);
		when "1001010101011111" => data_out <= rom_array(38239);
		when "1001010101100000" => data_out <= rom_array(38240);
		when "1001010101100001" => data_out <= rom_array(38241);
		when "1001010101100010" => data_out <= rom_array(38242);
		when "1001010101100011" => data_out <= rom_array(38243);
		when "1001010101100100" => data_out <= rom_array(38244);
		when "1001010101100101" => data_out <= rom_array(38245);
		when "1001010101100110" => data_out <= rom_array(38246);
		when "1001010101100111" => data_out <= rom_array(38247);
		when "1001010101101000" => data_out <= rom_array(38248);
		when "1001010101101001" => data_out <= rom_array(38249);
		when "1001010101101010" => data_out <= rom_array(38250);
		when "1001010101101011" => data_out <= rom_array(38251);
		when "1001010101101100" => data_out <= rom_array(38252);
		when "1001010101101101" => data_out <= rom_array(38253);
		when "1001010101101110" => data_out <= rom_array(38254);
		when "1001010101101111" => data_out <= rom_array(38255);
		when "1001010101110000" => data_out <= rom_array(38256);
		when "1001010101110001" => data_out <= rom_array(38257);
		when "1001010101110010" => data_out <= rom_array(38258);
		when "1001010101110011" => data_out <= rom_array(38259);
		when "1001010101110100" => data_out <= rom_array(38260);
		when "1001010101110101" => data_out <= rom_array(38261);
		when "1001010101110110" => data_out <= rom_array(38262);
		when "1001010101110111" => data_out <= rom_array(38263);
		when "1001010101111000" => data_out <= rom_array(38264);
		when "1001010101111001" => data_out <= rom_array(38265);
		when "1001010101111010" => data_out <= rom_array(38266);
		when "1001010101111011" => data_out <= rom_array(38267);
		when "1001010101111100" => data_out <= rom_array(38268);
		when "1001010101111101" => data_out <= rom_array(38269);
		when "1001010101111110" => data_out <= rom_array(38270);
		when "1001010101111111" => data_out <= rom_array(38271);
		when "1001010110000000" => data_out <= rom_array(38272);
		when "1001010110000001" => data_out <= rom_array(38273);
		when "1001010110000010" => data_out <= rom_array(38274);
		when "1001010110000011" => data_out <= rom_array(38275);
		when "1001010110000100" => data_out <= rom_array(38276);
		when "1001010110000101" => data_out <= rom_array(38277);
		when "1001010110000110" => data_out <= rom_array(38278);
		when "1001010110000111" => data_out <= rom_array(38279);
		when "1001010110001000" => data_out <= rom_array(38280);
		when "1001010110001001" => data_out <= rom_array(38281);
		when "1001010110001010" => data_out <= rom_array(38282);
		when "1001010110001011" => data_out <= rom_array(38283);
		when "1001010110001100" => data_out <= rom_array(38284);
		when "1001010110001101" => data_out <= rom_array(38285);
		when "1001010110001110" => data_out <= rom_array(38286);
		when "1001010110001111" => data_out <= rom_array(38287);
		when "1001010110010000" => data_out <= rom_array(38288);
		when "1001010110010001" => data_out <= rom_array(38289);
		when "1001010110010010" => data_out <= rom_array(38290);
		when "1001010110010011" => data_out <= rom_array(38291);
		when "1001010110010100" => data_out <= rom_array(38292);
		when "1001010110010101" => data_out <= rom_array(38293);
		when "1001010110010110" => data_out <= rom_array(38294);
		when "1001010110010111" => data_out <= rom_array(38295);
		when "1001010110011000" => data_out <= rom_array(38296);
		when "1001010110011001" => data_out <= rom_array(38297);
		when "1001010110011010" => data_out <= rom_array(38298);
		when "1001010110011011" => data_out <= rom_array(38299);
		when "1001010110011100" => data_out <= rom_array(38300);
		when "1001010110011101" => data_out <= rom_array(38301);
		when "1001010110011110" => data_out <= rom_array(38302);
		when "1001010110011111" => data_out <= rom_array(38303);
		when "1001010110100000" => data_out <= rom_array(38304);
		when "1001010110100001" => data_out <= rom_array(38305);
		when "1001010110100010" => data_out <= rom_array(38306);
		when "1001010110100011" => data_out <= rom_array(38307);
		when "1001010110100100" => data_out <= rom_array(38308);
		when "1001010110100101" => data_out <= rom_array(38309);
		when "1001010110100110" => data_out <= rom_array(38310);
		when "1001010110100111" => data_out <= rom_array(38311);
		when "1001010110101000" => data_out <= rom_array(38312);
		when "1001010110101001" => data_out <= rom_array(38313);
		when "1001010110101010" => data_out <= rom_array(38314);
		when "1001010110101011" => data_out <= rom_array(38315);
		when "1001010110101100" => data_out <= rom_array(38316);
		when "1001010110101101" => data_out <= rom_array(38317);
		when "1001010110101110" => data_out <= rom_array(38318);
		when "1001010110101111" => data_out <= rom_array(38319);
		when "1001010110110000" => data_out <= rom_array(38320);
		when "1001010110110001" => data_out <= rom_array(38321);
		when "1001010110110010" => data_out <= rom_array(38322);
		when "1001010110110011" => data_out <= rom_array(38323);
		when "1001010110110100" => data_out <= rom_array(38324);
		when "1001010110110101" => data_out <= rom_array(38325);
		when "1001010110110110" => data_out <= rom_array(38326);
		when "1001010110110111" => data_out <= rom_array(38327);
		when "1001010110111000" => data_out <= rom_array(38328);
		when "1001010110111001" => data_out <= rom_array(38329);
		when "1001010110111010" => data_out <= rom_array(38330);
		when "1001010110111011" => data_out <= rom_array(38331);
		when "1001010110111100" => data_out <= rom_array(38332);
		when "1001010110111101" => data_out <= rom_array(38333);
		when "1001010110111110" => data_out <= rom_array(38334);
		when "1001010110111111" => data_out <= rom_array(38335);
		when "1001010111000000" => data_out <= rom_array(38336);
		when "1001010111000001" => data_out <= rom_array(38337);
		when "1001010111000010" => data_out <= rom_array(38338);
		when "1001010111000011" => data_out <= rom_array(38339);
		when "1001010111000100" => data_out <= rom_array(38340);
		when "1001010111000101" => data_out <= rom_array(38341);
		when "1001010111000110" => data_out <= rom_array(38342);
		when "1001010111000111" => data_out <= rom_array(38343);
		when "1001010111001000" => data_out <= rom_array(38344);
		when "1001010111001001" => data_out <= rom_array(38345);
		when "1001010111001010" => data_out <= rom_array(38346);
		when "1001010111001011" => data_out <= rom_array(38347);
		when "1001010111001100" => data_out <= rom_array(38348);
		when "1001010111001101" => data_out <= rom_array(38349);
		when "1001010111001110" => data_out <= rom_array(38350);
		when "1001010111001111" => data_out <= rom_array(38351);
		when "1001010111010000" => data_out <= rom_array(38352);
		when "1001010111010001" => data_out <= rom_array(38353);
		when "1001010111010010" => data_out <= rom_array(38354);
		when "1001010111010011" => data_out <= rom_array(38355);
		when "1001010111010100" => data_out <= rom_array(38356);
		when "1001010111010101" => data_out <= rom_array(38357);
		when "1001010111010110" => data_out <= rom_array(38358);
		when "1001010111010111" => data_out <= rom_array(38359);
		when "1001010111011000" => data_out <= rom_array(38360);
		when "1001010111011001" => data_out <= rom_array(38361);
		when "1001010111011010" => data_out <= rom_array(38362);
		when "1001010111011011" => data_out <= rom_array(38363);
		when "1001010111011100" => data_out <= rom_array(38364);
		when "1001010111011101" => data_out <= rom_array(38365);
		when "1001010111011110" => data_out <= rom_array(38366);
		when "1001010111011111" => data_out <= rom_array(38367);
		when "1001010111100000" => data_out <= rom_array(38368);
		when "1001010111100001" => data_out <= rom_array(38369);
		when "1001010111100010" => data_out <= rom_array(38370);
		when "1001010111100011" => data_out <= rom_array(38371);
		when "1001010111100100" => data_out <= rom_array(38372);
		when "1001010111100101" => data_out <= rom_array(38373);
		when "1001010111100110" => data_out <= rom_array(38374);
		when "1001010111100111" => data_out <= rom_array(38375);
		when "1001010111101000" => data_out <= rom_array(38376);
		when "1001010111101001" => data_out <= rom_array(38377);
		when "1001010111101010" => data_out <= rom_array(38378);
		when "1001010111101011" => data_out <= rom_array(38379);
		when "1001010111101100" => data_out <= rom_array(38380);
		when "1001010111101101" => data_out <= rom_array(38381);
		when "1001010111101110" => data_out <= rom_array(38382);
		when "1001010111101111" => data_out <= rom_array(38383);
		when "1001010111110000" => data_out <= rom_array(38384);
		when "1001010111110001" => data_out <= rom_array(38385);
		when "1001010111110010" => data_out <= rom_array(38386);
		when "1001010111110011" => data_out <= rom_array(38387);
		when "1001010111110100" => data_out <= rom_array(38388);
		when "1001010111110101" => data_out <= rom_array(38389);
		when "1001010111110110" => data_out <= rom_array(38390);
		when "1001010111110111" => data_out <= rom_array(38391);
		when "1001010111111000" => data_out <= rom_array(38392);
		when "1001010111111001" => data_out <= rom_array(38393);
		when "1001010111111010" => data_out <= rom_array(38394);
		when "1001010111111011" => data_out <= rom_array(38395);
		when "1001010111111100" => data_out <= rom_array(38396);
		when "1001010111111101" => data_out <= rom_array(38397);
		when "1001010111111110" => data_out <= rom_array(38398);
		when "1001010111111111" => data_out <= rom_array(38399);
		when "1001011000000000" => data_out <= rom_array(38400);
		when "1001011000000001" => data_out <= rom_array(38401);
		when "1001011000000010" => data_out <= rom_array(38402);
		when "1001011000000011" => data_out <= rom_array(38403);
		when "1001011000000100" => data_out <= rom_array(38404);
		when "1001011000000101" => data_out <= rom_array(38405);
		when "1001011000000110" => data_out <= rom_array(38406);
		when "1001011000000111" => data_out <= rom_array(38407);
		when "1001011000001000" => data_out <= rom_array(38408);
		when "1001011000001001" => data_out <= rom_array(38409);
		when "1001011000001010" => data_out <= rom_array(38410);
		when "1001011000001011" => data_out <= rom_array(38411);
		when "1001011000001100" => data_out <= rom_array(38412);
		when "1001011000001101" => data_out <= rom_array(38413);
		when "1001011000001110" => data_out <= rom_array(38414);
		when "1001011000001111" => data_out <= rom_array(38415);
		when "1001011000010000" => data_out <= rom_array(38416);
		when "1001011000010001" => data_out <= rom_array(38417);
		when "1001011000010010" => data_out <= rom_array(38418);
		when "1001011000010011" => data_out <= rom_array(38419);
		when "1001011000010100" => data_out <= rom_array(38420);
		when "1001011000010101" => data_out <= rom_array(38421);
		when "1001011000010110" => data_out <= rom_array(38422);
		when "1001011000010111" => data_out <= rom_array(38423);
		when "1001011000011000" => data_out <= rom_array(38424);
		when "1001011000011001" => data_out <= rom_array(38425);
		when "1001011000011010" => data_out <= rom_array(38426);
		when "1001011000011011" => data_out <= rom_array(38427);
		when "1001011000011100" => data_out <= rom_array(38428);
		when "1001011000011101" => data_out <= rom_array(38429);
		when "1001011000011110" => data_out <= rom_array(38430);
		when "1001011000011111" => data_out <= rom_array(38431);
		when "1001011000100000" => data_out <= rom_array(38432);
		when "1001011000100001" => data_out <= rom_array(38433);
		when "1001011000100010" => data_out <= rom_array(38434);
		when "1001011000100011" => data_out <= rom_array(38435);
		when "1001011000100100" => data_out <= rom_array(38436);
		when "1001011000100101" => data_out <= rom_array(38437);
		when "1001011000100110" => data_out <= rom_array(38438);
		when "1001011000100111" => data_out <= rom_array(38439);
		when "1001011000101000" => data_out <= rom_array(38440);
		when "1001011000101001" => data_out <= rom_array(38441);
		when "1001011000101010" => data_out <= rom_array(38442);
		when "1001011000101011" => data_out <= rom_array(38443);
		when "1001011000101100" => data_out <= rom_array(38444);
		when "1001011000101101" => data_out <= rom_array(38445);
		when "1001011000101110" => data_out <= rom_array(38446);
		when "1001011000101111" => data_out <= rom_array(38447);
		when "1001011000110000" => data_out <= rom_array(38448);
		when "1001011000110001" => data_out <= rom_array(38449);
		when "1001011000110010" => data_out <= rom_array(38450);
		when "1001011000110011" => data_out <= rom_array(38451);
		when "1001011000110100" => data_out <= rom_array(38452);
		when "1001011000110101" => data_out <= rom_array(38453);
		when "1001011000110110" => data_out <= rom_array(38454);
		when "1001011000110111" => data_out <= rom_array(38455);
		when "1001011000111000" => data_out <= rom_array(38456);
		when "1001011000111001" => data_out <= rom_array(38457);
		when "1001011000111010" => data_out <= rom_array(38458);
		when "1001011000111011" => data_out <= rom_array(38459);
		when "1001011000111100" => data_out <= rom_array(38460);
		when "1001011000111101" => data_out <= rom_array(38461);
		when "1001011000111110" => data_out <= rom_array(38462);
		when "1001011000111111" => data_out <= rom_array(38463);
		when "1001011001000000" => data_out <= rom_array(38464);
		when "1001011001000001" => data_out <= rom_array(38465);
		when "1001011001000010" => data_out <= rom_array(38466);
		when "1001011001000011" => data_out <= rom_array(38467);
		when "1001011001000100" => data_out <= rom_array(38468);
		when "1001011001000101" => data_out <= rom_array(38469);
		when "1001011001000110" => data_out <= rom_array(38470);
		when "1001011001000111" => data_out <= rom_array(38471);
		when "1001011001001000" => data_out <= rom_array(38472);
		when "1001011001001001" => data_out <= rom_array(38473);
		when "1001011001001010" => data_out <= rom_array(38474);
		when "1001011001001011" => data_out <= rom_array(38475);
		when "1001011001001100" => data_out <= rom_array(38476);
		when "1001011001001101" => data_out <= rom_array(38477);
		when "1001011001001110" => data_out <= rom_array(38478);
		when "1001011001001111" => data_out <= rom_array(38479);
		when "1001011001010000" => data_out <= rom_array(38480);
		when "1001011001010001" => data_out <= rom_array(38481);
		when "1001011001010010" => data_out <= rom_array(38482);
		when "1001011001010011" => data_out <= rom_array(38483);
		when "1001011001010100" => data_out <= rom_array(38484);
		when "1001011001010101" => data_out <= rom_array(38485);
		when "1001011001010110" => data_out <= rom_array(38486);
		when "1001011001010111" => data_out <= rom_array(38487);
		when "1001011001011000" => data_out <= rom_array(38488);
		when "1001011001011001" => data_out <= rom_array(38489);
		when "1001011001011010" => data_out <= rom_array(38490);
		when "1001011001011011" => data_out <= rom_array(38491);
		when "1001011001011100" => data_out <= rom_array(38492);
		when "1001011001011101" => data_out <= rom_array(38493);
		when "1001011001011110" => data_out <= rom_array(38494);
		when "1001011001011111" => data_out <= rom_array(38495);
		when "1001011001100000" => data_out <= rom_array(38496);
		when "1001011001100001" => data_out <= rom_array(38497);
		when "1001011001100010" => data_out <= rom_array(38498);
		when "1001011001100011" => data_out <= rom_array(38499);
		when "1001011001100100" => data_out <= rom_array(38500);
		when "1001011001100101" => data_out <= rom_array(38501);
		when "1001011001100110" => data_out <= rom_array(38502);
		when "1001011001100111" => data_out <= rom_array(38503);
		when "1001011001101000" => data_out <= rom_array(38504);
		when "1001011001101001" => data_out <= rom_array(38505);
		when "1001011001101010" => data_out <= rom_array(38506);
		when "1001011001101011" => data_out <= rom_array(38507);
		when "1001011001101100" => data_out <= rom_array(38508);
		when "1001011001101101" => data_out <= rom_array(38509);
		when "1001011001101110" => data_out <= rom_array(38510);
		when "1001011001101111" => data_out <= rom_array(38511);
		when "1001011001110000" => data_out <= rom_array(38512);
		when "1001011001110001" => data_out <= rom_array(38513);
		when "1001011001110010" => data_out <= rom_array(38514);
		when "1001011001110011" => data_out <= rom_array(38515);
		when "1001011001110100" => data_out <= rom_array(38516);
		when "1001011001110101" => data_out <= rom_array(38517);
		when "1001011001110110" => data_out <= rom_array(38518);
		when "1001011001110111" => data_out <= rom_array(38519);
		when "1001011001111000" => data_out <= rom_array(38520);
		when "1001011001111001" => data_out <= rom_array(38521);
		when "1001011001111010" => data_out <= rom_array(38522);
		when "1001011001111011" => data_out <= rom_array(38523);
		when "1001011001111100" => data_out <= rom_array(38524);
		when "1001011001111101" => data_out <= rom_array(38525);
		when "1001011001111110" => data_out <= rom_array(38526);
		when "1001011001111111" => data_out <= rom_array(38527);
		when "1001011010000000" => data_out <= rom_array(38528);
		when "1001011010000001" => data_out <= rom_array(38529);
		when "1001011010000010" => data_out <= rom_array(38530);
		when "1001011010000011" => data_out <= rom_array(38531);
		when "1001011010000100" => data_out <= rom_array(38532);
		when "1001011010000101" => data_out <= rom_array(38533);
		when "1001011010000110" => data_out <= rom_array(38534);
		when "1001011010000111" => data_out <= rom_array(38535);
		when "1001011010001000" => data_out <= rom_array(38536);
		when "1001011010001001" => data_out <= rom_array(38537);
		when "1001011010001010" => data_out <= rom_array(38538);
		when "1001011010001011" => data_out <= rom_array(38539);
		when "1001011010001100" => data_out <= rom_array(38540);
		when "1001011010001101" => data_out <= rom_array(38541);
		when "1001011010001110" => data_out <= rom_array(38542);
		when "1001011010001111" => data_out <= rom_array(38543);
		when "1001011010010000" => data_out <= rom_array(38544);
		when "1001011010010001" => data_out <= rom_array(38545);
		when "1001011010010010" => data_out <= rom_array(38546);
		when "1001011010010011" => data_out <= rom_array(38547);
		when "1001011010010100" => data_out <= rom_array(38548);
		when "1001011010010101" => data_out <= rom_array(38549);
		when "1001011010010110" => data_out <= rom_array(38550);
		when "1001011010010111" => data_out <= rom_array(38551);
		when "1001011010011000" => data_out <= rom_array(38552);
		when "1001011010011001" => data_out <= rom_array(38553);
		when "1001011010011010" => data_out <= rom_array(38554);
		when "1001011010011011" => data_out <= rom_array(38555);
		when "1001011010011100" => data_out <= rom_array(38556);
		when "1001011010011101" => data_out <= rom_array(38557);
		when "1001011010011110" => data_out <= rom_array(38558);
		when "1001011010011111" => data_out <= rom_array(38559);
		when "1001011010100000" => data_out <= rom_array(38560);
		when "1001011010100001" => data_out <= rom_array(38561);
		when "1001011010100010" => data_out <= rom_array(38562);
		when "1001011010100011" => data_out <= rom_array(38563);
		when "1001011010100100" => data_out <= rom_array(38564);
		when "1001011010100101" => data_out <= rom_array(38565);
		when "1001011010100110" => data_out <= rom_array(38566);
		when "1001011010100111" => data_out <= rom_array(38567);
		when "1001011010101000" => data_out <= rom_array(38568);
		when "1001011010101001" => data_out <= rom_array(38569);
		when "1001011010101010" => data_out <= rom_array(38570);
		when "1001011010101011" => data_out <= rom_array(38571);
		when "1001011010101100" => data_out <= rom_array(38572);
		when "1001011010101101" => data_out <= rom_array(38573);
		when "1001011010101110" => data_out <= rom_array(38574);
		when "1001011010101111" => data_out <= rom_array(38575);
		when "1001011010110000" => data_out <= rom_array(38576);
		when "1001011010110001" => data_out <= rom_array(38577);
		when "1001011010110010" => data_out <= rom_array(38578);
		when "1001011010110011" => data_out <= rom_array(38579);
		when "1001011010110100" => data_out <= rom_array(38580);
		when "1001011010110101" => data_out <= rom_array(38581);
		when "1001011010110110" => data_out <= rom_array(38582);
		when "1001011010110111" => data_out <= rom_array(38583);
		when "1001011010111000" => data_out <= rom_array(38584);
		when "1001011010111001" => data_out <= rom_array(38585);
		when "1001011010111010" => data_out <= rom_array(38586);
		when "1001011010111011" => data_out <= rom_array(38587);
		when "1001011010111100" => data_out <= rom_array(38588);
		when "1001011010111101" => data_out <= rom_array(38589);
		when "1001011010111110" => data_out <= rom_array(38590);
		when "1001011010111111" => data_out <= rom_array(38591);
		when "1001011011000000" => data_out <= rom_array(38592);
		when "1001011011000001" => data_out <= rom_array(38593);
		when "1001011011000010" => data_out <= rom_array(38594);
		when "1001011011000011" => data_out <= rom_array(38595);
		when "1001011011000100" => data_out <= rom_array(38596);
		when "1001011011000101" => data_out <= rom_array(38597);
		when "1001011011000110" => data_out <= rom_array(38598);
		when "1001011011000111" => data_out <= rom_array(38599);
		when "1001011011001000" => data_out <= rom_array(38600);
		when "1001011011001001" => data_out <= rom_array(38601);
		when "1001011011001010" => data_out <= rom_array(38602);
		when "1001011011001011" => data_out <= rom_array(38603);
		when "1001011011001100" => data_out <= rom_array(38604);
		when "1001011011001101" => data_out <= rom_array(38605);
		when "1001011011001110" => data_out <= rom_array(38606);
		when "1001011011001111" => data_out <= rom_array(38607);
		when "1001011011010000" => data_out <= rom_array(38608);
		when "1001011011010001" => data_out <= rom_array(38609);
		when "1001011011010010" => data_out <= rom_array(38610);
		when "1001011011010011" => data_out <= rom_array(38611);
		when "1001011011010100" => data_out <= rom_array(38612);
		when "1001011011010101" => data_out <= rom_array(38613);
		when "1001011011010110" => data_out <= rom_array(38614);
		when "1001011011010111" => data_out <= rom_array(38615);
		when "1001011011011000" => data_out <= rom_array(38616);
		when "1001011011011001" => data_out <= rom_array(38617);
		when "1001011011011010" => data_out <= rom_array(38618);
		when "1001011011011011" => data_out <= rom_array(38619);
		when "1001011011011100" => data_out <= rom_array(38620);
		when "1001011011011101" => data_out <= rom_array(38621);
		when "1001011011011110" => data_out <= rom_array(38622);
		when "1001011011011111" => data_out <= rom_array(38623);
		when "1001011011100000" => data_out <= rom_array(38624);
		when "1001011011100001" => data_out <= rom_array(38625);
		when "1001011011100010" => data_out <= rom_array(38626);
		when "1001011011100011" => data_out <= rom_array(38627);
		when "1001011011100100" => data_out <= rom_array(38628);
		when "1001011011100101" => data_out <= rom_array(38629);
		when "1001011011100110" => data_out <= rom_array(38630);
		when "1001011011100111" => data_out <= rom_array(38631);
		when "1001011011101000" => data_out <= rom_array(38632);
		when "1001011011101001" => data_out <= rom_array(38633);
		when "1001011011101010" => data_out <= rom_array(38634);
		when "1001011011101011" => data_out <= rom_array(38635);
		when "1001011011101100" => data_out <= rom_array(38636);
		when "1001011011101101" => data_out <= rom_array(38637);
		when "1001011011101110" => data_out <= rom_array(38638);
		when "1001011011101111" => data_out <= rom_array(38639);
		when "1001011011110000" => data_out <= rom_array(38640);
		when "1001011011110001" => data_out <= rom_array(38641);
		when "1001011011110010" => data_out <= rom_array(38642);
		when "1001011011110011" => data_out <= rom_array(38643);
		when "1001011011110100" => data_out <= rom_array(38644);
		when "1001011011110101" => data_out <= rom_array(38645);
		when "1001011011110110" => data_out <= rom_array(38646);
		when "1001011011110111" => data_out <= rom_array(38647);
		when "1001011011111000" => data_out <= rom_array(38648);
		when "1001011011111001" => data_out <= rom_array(38649);
		when "1001011011111010" => data_out <= rom_array(38650);
		when "1001011011111011" => data_out <= rom_array(38651);
		when "1001011011111100" => data_out <= rom_array(38652);
		when "1001011011111101" => data_out <= rom_array(38653);
		when "1001011011111110" => data_out <= rom_array(38654);
		when "1001011011111111" => data_out <= rom_array(38655);
		when "1001011100000000" => data_out <= rom_array(38656);
		when "1001011100000001" => data_out <= rom_array(38657);
		when "1001011100000010" => data_out <= rom_array(38658);
		when "1001011100000011" => data_out <= rom_array(38659);
		when "1001011100000100" => data_out <= rom_array(38660);
		when "1001011100000101" => data_out <= rom_array(38661);
		when "1001011100000110" => data_out <= rom_array(38662);
		when "1001011100000111" => data_out <= rom_array(38663);
		when "1001011100001000" => data_out <= rom_array(38664);
		when "1001011100001001" => data_out <= rom_array(38665);
		when "1001011100001010" => data_out <= rom_array(38666);
		when "1001011100001011" => data_out <= rom_array(38667);
		when "1001011100001100" => data_out <= rom_array(38668);
		when "1001011100001101" => data_out <= rom_array(38669);
		when "1001011100001110" => data_out <= rom_array(38670);
		when "1001011100001111" => data_out <= rom_array(38671);
		when "1001011100010000" => data_out <= rom_array(38672);
		when "1001011100010001" => data_out <= rom_array(38673);
		when "1001011100010010" => data_out <= rom_array(38674);
		when "1001011100010011" => data_out <= rom_array(38675);
		when "1001011100010100" => data_out <= rom_array(38676);
		when "1001011100010101" => data_out <= rom_array(38677);
		when "1001011100010110" => data_out <= rom_array(38678);
		when "1001011100010111" => data_out <= rom_array(38679);
		when "1001011100011000" => data_out <= rom_array(38680);
		when "1001011100011001" => data_out <= rom_array(38681);
		when "1001011100011010" => data_out <= rom_array(38682);
		when "1001011100011011" => data_out <= rom_array(38683);
		when "1001011100011100" => data_out <= rom_array(38684);
		when "1001011100011101" => data_out <= rom_array(38685);
		when "1001011100011110" => data_out <= rom_array(38686);
		when "1001011100011111" => data_out <= rom_array(38687);
		when "1001011100100000" => data_out <= rom_array(38688);
		when "1001011100100001" => data_out <= rom_array(38689);
		when "1001011100100010" => data_out <= rom_array(38690);
		when "1001011100100011" => data_out <= rom_array(38691);
		when "1001011100100100" => data_out <= rom_array(38692);
		when "1001011100100101" => data_out <= rom_array(38693);
		when "1001011100100110" => data_out <= rom_array(38694);
		when "1001011100100111" => data_out <= rom_array(38695);
		when "1001011100101000" => data_out <= rom_array(38696);
		when "1001011100101001" => data_out <= rom_array(38697);
		when "1001011100101010" => data_out <= rom_array(38698);
		when "1001011100101011" => data_out <= rom_array(38699);
		when "1001011100101100" => data_out <= rom_array(38700);
		when "1001011100101101" => data_out <= rom_array(38701);
		when "1001011100101110" => data_out <= rom_array(38702);
		when "1001011100101111" => data_out <= rom_array(38703);
		when "1001011100110000" => data_out <= rom_array(38704);
		when "1001011100110001" => data_out <= rom_array(38705);
		when "1001011100110010" => data_out <= rom_array(38706);
		when "1001011100110011" => data_out <= rom_array(38707);
		when "1001011100110100" => data_out <= rom_array(38708);
		when "1001011100110101" => data_out <= rom_array(38709);
		when "1001011100110110" => data_out <= rom_array(38710);
		when "1001011100110111" => data_out <= rom_array(38711);
		when "1001011100111000" => data_out <= rom_array(38712);
		when "1001011100111001" => data_out <= rom_array(38713);
		when "1001011100111010" => data_out <= rom_array(38714);
		when "1001011100111011" => data_out <= rom_array(38715);
		when "1001011100111100" => data_out <= rom_array(38716);
		when "1001011100111101" => data_out <= rom_array(38717);
		when "1001011100111110" => data_out <= rom_array(38718);
		when "1001011100111111" => data_out <= rom_array(38719);
		when "1001011101000000" => data_out <= rom_array(38720);
		when "1001011101000001" => data_out <= rom_array(38721);
		when "1001011101000010" => data_out <= rom_array(38722);
		when "1001011101000011" => data_out <= rom_array(38723);
		when "1001011101000100" => data_out <= rom_array(38724);
		when "1001011101000101" => data_out <= rom_array(38725);
		when "1001011101000110" => data_out <= rom_array(38726);
		when "1001011101000111" => data_out <= rom_array(38727);
		when "1001011101001000" => data_out <= rom_array(38728);
		when "1001011101001001" => data_out <= rom_array(38729);
		when "1001011101001010" => data_out <= rom_array(38730);
		when "1001011101001011" => data_out <= rom_array(38731);
		when "1001011101001100" => data_out <= rom_array(38732);
		when "1001011101001101" => data_out <= rom_array(38733);
		when "1001011101001110" => data_out <= rom_array(38734);
		when "1001011101001111" => data_out <= rom_array(38735);
		when "1001011101010000" => data_out <= rom_array(38736);
		when "1001011101010001" => data_out <= rom_array(38737);
		when "1001011101010010" => data_out <= rom_array(38738);
		when "1001011101010011" => data_out <= rom_array(38739);
		when "1001011101010100" => data_out <= rom_array(38740);
		when "1001011101010101" => data_out <= rom_array(38741);
		when "1001011101010110" => data_out <= rom_array(38742);
		when "1001011101010111" => data_out <= rom_array(38743);
		when "1001011101011000" => data_out <= rom_array(38744);
		when "1001011101011001" => data_out <= rom_array(38745);
		when "1001011101011010" => data_out <= rom_array(38746);
		when "1001011101011011" => data_out <= rom_array(38747);
		when "1001011101011100" => data_out <= rom_array(38748);
		when "1001011101011101" => data_out <= rom_array(38749);
		when "1001011101011110" => data_out <= rom_array(38750);
		when "1001011101011111" => data_out <= rom_array(38751);
		when "1001011101100000" => data_out <= rom_array(38752);
		when "1001011101100001" => data_out <= rom_array(38753);
		when "1001011101100010" => data_out <= rom_array(38754);
		when "1001011101100011" => data_out <= rom_array(38755);
		when "1001011101100100" => data_out <= rom_array(38756);
		when "1001011101100101" => data_out <= rom_array(38757);
		when "1001011101100110" => data_out <= rom_array(38758);
		when "1001011101100111" => data_out <= rom_array(38759);
		when "1001011101101000" => data_out <= rom_array(38760);
		when "1001011101101001" => data_out <= rom_array(38761);
		when "1001011101101010" => data_out <= rom_array(38762);
		when "1001011101101011" => data_out <= rom_array(38763);
		when "1001011101101100" => data_out <= rom_array(38764);
		when "1001011101101101" => data_out <= rom_array(38765);
		when "1001011101101110" => data_out <= rom_array(38766);
		when "1001011101101111" => data_out <= rom_array(38767);
		when "1001011101110000" => data_out <= rom_array(38768);
		when "1001011101110001" => data_out <= rom_array(38769);
		when "1001011101110010" => data_out <= rom_array(38770);
		when "1001011101110011" => data_out <= rom_array(38771);
		when "1001011101110100" => data_out <= rom_array(38772);
		when "1001011101110101" => data_out <= rom_array(38773);
		when "1001011101110110" => data_out <= rom_array(38774);
		when "1001011101110111" => data_out <= rom_array(38775);
		when "1001011101111000" => data_out <= rom_array(38776);
		when "1001011101111001" => data_out <= rom_array(38777);
		when "1001011101111010" => data_out <= rom_array(38778);
		when "1001011101111011" => data_out <= rom_array(38779);
		when "1001011101111100" => data_out <= rom_array(38780);
		when "1001011101111101" => data_out <= rom_array(38781);
		when "1001011101111110" => data_out <= rom_array(38782);
		when "1001011101111111" => data_out <= rom_array(38783);
		when "1001011110000000" => data_out <= rom_array(38784);
		when "1001011110000001" => data_out <= rom_array(38785);
		when "1001011110000010" => data_out <= rom_array(38786);
		when "1001011110000011" => data_out <= rom_array(38787);
		when "1001011110000100" => data_out <= rom_array(38788);
		when "1001011110000101" => data_out <= rom_array(38789);
		when "1001011110000110" => data_out <= rom_array(38790);
		when "1001011110000111" => data_out <= rom_array(38791);
		when "1001011110001000" => data_out <= rom_array(38792);
		when "1001011110001001" => data_out <= rom_array(38793);
		when "1001011110001010" => data_out <= rom_array(38794);
		when "1001011110001011" => data_out <= rom_array(38795);
		when "1001011110001100" => data_out <= rom_array(38796);
		when "1001011110001101" => data_out <= rom_array(38797);
		when "1001011110001110" => data_out <= rom_array(38798);
		when "1001011110001111" => data_out <= rom_array(38799);
		when "1001011110010000" => data_out <= rom_array(38800);
		when "1001011110010001" => data_out <= rom_array(38801);
		when "1001011110010010" => data_out <= rom_array(38802);
		when "1001011110010011" => data_out <= rom_array(38803);
		when "1001011110010100" => data_out <= rom_array(38804);
		when "1001011110010101" => data_out <= rom_array(38805);
		when "1001011110010110" => data_out <= rom_array(38806);
		when "1001011110010111" => data_out <= rom_array(38807);
		when "1001011110011000" => data_out <= rom_array(38808);
		when "1001011110011001" => data_out <= rom_array(38809);
		when "1001011110011010" => data_out <= rom_array(38810);
		when "1001011110011011" => data_out <= rom_array(38811);
		when "1001011110011100" => data_out <= rom_array(38812);
		when "1001011110011101" => data_out <= rom_array(38813);
		when "1001011110011110" => data_out <= rom_array(38814);
		when "1001011110011111" => data_out <= rom_array(38815);
		when "1001011110100000" => data_out <= rom_array(38816);
		when "1001011110100001" => data_out <= rom_array(38817);
		when "1001011110100010" => data_out <= rom_array(38818);
		when "1001011110100011" => data_out <= rom_array(38819);
		when "1001011110100100" => data_out <= rom_array(38820);
		when "1001011110100101" => data_out <= rom_array(38821);
		when "1001011110100110" => data_out <= rom_array(38822);
		when "1001011110100111" => data_out <= rom_array(38823);
		when "1001011110101000" => data_out <= rom_array(38824);
		when "1001011110101001" => data_out <= rom_array(38825);
		when "1001011110101010" => data_out <= rom_array(38826);
		when "1001011110101011" => data_out <= rom_array(38827);
		when "1001011110101100" => data_out <= rom_array(38828);
		when "1001011110101101" => data_out <= rom_array(38829);
		when "1001011110101110" => data_out <= rom_array(38830);
		when "1001011110101111" => data_out <= rom_array(38831);
		when "1001011110110000" => data_out <= rom_array(38832);
		when "1001011110110001" => data_out <= rom_array(38833);
		when "1001011110110010" => data_out <= rom_array(38834);
		when "1001011110110011" => data_out <= rom_array(38835);
		when "1001011110110100" => data_out <= rom_array(38836);
		when "1001011110110101" => data_out <= rom_array(38837);
		when "1001011110110110" => data_out <= rom_array(38838);
		when "1001011110110111" => data_out <= rom_array(38839);
		when "1001011110111000" => data_out <= rom_array(38840);
		when "1001011110111001" => data_out <= rom_array(38841);
		when "1001011110111010" => data_out <= rom_array(38842);
		when "1001011110111011" => data_out <= rom_array(38843);
		when "1001011110111100" => data_out <= rom_array(38844);
		when "1001011110111101" => data_out <= rom_array(38845);
		when "1001011110111110" => data_out <= rom_array(38846);
		when "1001011110111111" => data_out <= rom_array(38847);
		when "1001011111000000" => data_out <= rom_array(38848);
		when "1001011111000001" => data_out <= rom_array(38849);
		when "1001011111000010" => data_out <= rom_array(38850);
		when "1001011111000011" => data_out <= rom_array(38851);
		when "1001011111000100" => data_out <= rom_array(38852);
		when "1001011111000101" => data_out <= rom_array(38853);
		when "1001011111000110" => data_out <= rom_array(38854);
		when "1001011111000111" => data_out <= rom_array(38855);
		when "1001011111001000" => data_out <= rom_array(38856);
		when "1001011111001001" => data_out <= rom_array(38857);
		when "1001011111001010" => data_out <= rom_array(38858);
		when "1001011111001011" => data_out <= rom_array(38859);
		when "1001011111001100" => data_out <= rom_array(38860);
		when "1001011111001101" => data_out <= rom_array(38861);
		when "1001011111001110" => data_out <= rom_array(38862);
		when "1001011111001111" => data_out <= rom_array(38863);
		when "1001011111010000" => data_out <= rom_array(38864);
		when "1001011111010001" => data_out <= rom_array(38865);
		when "1001011111010010" => data_out <= rom_array(38866);
		when "1001011111010011" => data_out <= rom_array(38867);
		when "1001011111010100" => data_out <= rom_array(38868);
		when "1001011111010101" => data_out <= rom_array(38869);
		when "1001011111010110" => data_out <= rom_array(38870);
		when "1001011111010111" => data_out <= rom_array(38871);
		when "1001011111011000" => data_out <= rom_array(38872);
		when "1001011111011001" => data_out <= rom_array(38873);
		when "1001011111011010" => data_out <= rom_array(38874);
		when "1001011111011011" => data_out <= rom_array(38875);
		when "1001011111011100" => data_out <= rom_array(38876);
		when "1001011111011101" => data_out <= rom_array(38877);
		when "1001011111011110" => data_out <= rom_array(38878);
		when "1001011111011111" => data_out <= rom_array(38879);
		when "1001011111100000" => data_out <= rom_array(38880);
		when "1001011111100001" => data_out <= rom_array(38881);
		when "1001011111100010" => data_out <= rom_array(38882);
		when "1001011111100011" => data_out <= rom_array(38883);
		when "1001011111100100" => data_out <= rom_array(38884);
		when "1001011111100101" => data_out <= rom_array(38885);
		when "1001011111100110" => data_out <= rom_array(38886);
		when "1001011111100111" => data_out <= rom_array(38887);
		when "1001011111101000" => data_out <= rom_array(38888);
		when "1001011111101001" => data_out <= rom_array(38889);
		when "1001011111101010" => data_out <= rom_array(38890);
		when "1001011111101011" => data_out <= rom_array(38891);
		when "1001011111101100" => data_out <= rom_array(38892);
		when "1001011111101101" => data_out <= rom_array(38893);
		when "1001011111101110" => data_out <= rom_array(38894);
		when "1001011111101111" => data_out <= rom_array(38895);
		when "1001011111110000" => data_out <= rom_array(38896);
		when "1001011111110001" => data_out <= rom_array(38897);
		when "1001011111110010" => data_out <= rom_array(38898);
		when "1001011111110011" => data_out <= rom_array(38899);
		when "1001011111110100" => data_out <= rom_array(38900);
		when "1001011111110101" => data_out <= rom_array(38901);
		when "1001011111110110" => data_out <= rom_array(38902);
		when "1001011111110111" => data_out <= rom_array(38903);
		when "1001011111111000" => data_out <= rom_array(38904);
		when "1001011111111001" => data_out <= rom_array(38905);
		when "1001011111111010" => data_out <= rom_array(38906);
		when "1001011111111011" => data_out <= rom_array(38907);
		when "1001011111111100" => data_out <= rom_array(38908);
		when "1001011111111101" => data_out <= rom_array(38909);
		when "1001011111111110" => data_out <= rom_array(38910);
		when "1001011111111111" => data_out <= rom_array(38911);
		when "1001100000000000" => data_out <= rom_array(38912);
		when "1001100000000001" => data_out <= rom_array(38913);
		when "1001100000000010" => data_out <= rom_array(38914);
		when "1001100000000011" => data_out <= rom_array(38915);
		when "1001100000000100" => data_out <= rom_array(38916);
		when "1001100000000101" => data_out <= rom_array(38917);
		when "1001100000000110" => data_out <= rom_array(38918);
		when "1001100000000111" => data_out <= rom_array(38919);
		when "1001100000001000" => data_out <= rom_array(38920);
		when "1001100000001001" => data_out <= rom_array(38921);
		when "1001100000001010" => data_out <= rom_array(38922);
		when "1001100000001011" => data_out <= rom_array(38923);
		when "1001100000001100" => data_out <= rom_array(38924);
		when "1001100000001101" => data_out <= rom_array(38925);
		when "1001100000001110" => data_out <= rom_array(38926);
		when "1001100000001111" => data_out <= rom_array(38927);
		when "1001100000010000" => data_out <= rom_array(38928);
		when "1001100000010001" => data_out <= rom_array(38929);
		when "1001100000010010" => data_out <= rom_array(38930);
		when "1001100000010011" => data_out <= rom_array(38931);
		when "1001100000010100" => data_out <= rom_array(38932);
		when "1001100000010101" => data_out <= rom_array(38933);
		when "1001100000010110" => data_out <= rom_array(38934);
		when "1001100000010111" => data_out <= rom_array(38935);
		when "1001100000011000" => data_out <= rom_array(38936);
		when "1001100000011001" => data_out <= rom_array(38937);
		when "1001100000011010" => data_out <= rom_array(38938);
		when "1001100000011011" => data_out <= rom_array(38939);
		when "1001100000011100" => data_out <= rom_array(38940);
		when "1001100000011101" => data_out <= rom_array(38941);
		when "1001100000011110" => data_out <= rom_array(38942);
		when "1001100000011111" => data_out <= rom_array(38943);
		when "1001100000100000" => data_out <= rom_array(38944);
		when "1001100000100001" => data_out <= rom_array(38945);
		when "1001100000100010" => data_out <= rom_array(38946);
		when "1001100000100011" => data_out <= rom_array(38947);
		when "1001100000100100" => data_out <= rom_array(38948);
		when "1001100000100101" => data_out <= rom_array(38949);
		when "1001100000100110" => data_out <= rom_array(38950);
		when "1001100000100111" => data_out <= rom_array(38951);
		when "1001100000101000" => data_out <= rom_array(38952);
		when "1001100000101001" => data_out <= rom_array(38953);
		when "1001100000101010" => data_out <= rom_array(38954);
		when "1001100000101011" => data_out <= rom_array(38955);
		when "1001100000101100" => data_out <= rom_array(38956);
		when "1001100000101101" => data_out <= rom_array(38957);
		when "1001100000101110" => data_out <= rom_array(38958);
		when "1001100000101111" => data_out <= rom_array(38959);
		when "1001100000110000" => data_out <= rom_array(38960);
		when "1001100000110001" => data_out <= rom_array(38961);
		when "1001100000110010" => data_out <= rom_array(38962);
		when "1001100000110011" => data_out <= rom_array(38963);
		when "1001100000110100" => data_out <= rom_array(38964);
		when "1001100000110101" => data_out <= rom_array(38965);
		when "1001100000110110" => data_out <= rom_array(38966);
		when "1001100000110111" => data_out <= rom_array(38967);
		when "1001100000111000" => data_out <= rom_array(38968);
		when "1001100000111001" => data_out <= rom_array(38969);
		when "1001100000111010" => data_out <= rom_array(38970);
		when "1001100000111011" => data_out <= rom_array(38971);
		when "1001100000111100" => data_out <= rom_array(38972);
		when "1001100000111101" => data_out <= rom_array(38973);
		when "1001100000111110" => data_out <= rom_array(38974);
		when "1001100000111111" => data_out <= rom_array(38975);
		when "1001100001000000" => data_out <= rom_array(38976);
		when "1001100001000001" => data_out <= rom_array(38977);
		when "1001100001000010" => data_out <= rom_array(38978);
		when "1001100001000011" => data_out <= rom_array(38979);
		when "1001100001000100" => data_out <= rom_array(38980);
		when "1001100001000101" => data_out <= rom_array(38981);
		when "1001100001000110" => data_out <= rom_array(38982);
		when "1001100001000111" => data_out <= rom_array(38983);
		when "1001100001001000" => data_out <= rom_array(38984);
		when "1001100001001001" => data_out <= rom_array(38985);
		when "1001100001001010" => data_out <= rom_array(38986);
		when "1001100001001011" => data_out <= rom_array(38987);
		when "1001100001001100" => data_out <= rom_array(38988);
		when "1001100001001101" => data_out <= rom_array(38989);
		when "1001100001001110" => data_out <= rom_array(38990);
		when "1001100001001111" => data_out <= rom_array(38991);
		when "1001100001010000" => data_out <= rom_array(38992);
		when "1001100001010001" => data_out <= rom_array(38993);
		when "1001100001010010" => data_out <= rom_array(38994);
		when "1001100001010011" => data_out <= rom_array(38995);
		when "1001100001010100" => data_out <= rom_array(38996);
		when "1001100001010101" => data_out <= rom_array(38997);
		when "1001100001010110" => data_out <= rom_array(38998);
		when "1001100001010111" => data_out <= rom_array(38999);
		when "1001100001011000" => data_out <= rom_array(39000);
		when "1001100001011001" => data_out <= rom_array(39001);
		when "1001100001011010" => data_out <= rom_array(39002);
		when "1001100001011011" => data_out <= rom_array(39003);
		when "1001100001011100" => data_out <= rom_array(39004);
		when "1001100001011101" => data_out <= rom_array(39005);
		when "1001100001011110" => data_out <= rom_array(39006);
		when "1001100001011111" => data_out <= rom_array(39007);
		when "1001100001100000" => data_out <= rom_array(39008);
		when "1001100001100001" => data_out <= rom_array(39009);
		when "1001100001100010" => data_out <= rom_array(39010);
		when "1001100001100011" => data_out <= rom_array(39011);
		when "1001100001100100" => data_out <= rom_array(39012);
		when "1001100001100101" => data_out <= rom_array(39013);
		when "1001100001100110" => data_out <= rom_array(39014);
		when "1001100001100111" => data_out <= rom_array(39015);
		when "1001100001101000" => data_out <= rom_array(39016);
		when "1001100001101001" => data_out <= rom_array(39017);
		when "1001100001101010" => data_out <= rom_array(39018);
		when "1001100001101011" => data_out <= rom_array(39019);
		when "1001100001101100" => data_out <= rom_array(39020);
		when "1001100001101101" => data_out <= rom_array(39021);
		when "1001100001101110" => data_out <= rom_array(39022);
		when "1001100001101111" => data_out <= rom_array(39023);
		when "1001100001110000" => data_out <= rom_array(39024);
		when "1001100001110001" => data_out <= rom_array(39025);
		when "1001100001110010" => data_out <= rom_array(39026);
		when "1001100001110011" => data_out <= rom_array(39027);
		when "1001100001110100" => data_out <= rom_array(39028);
		when "1001100001110101" => data_out <= rom_array(39029);
		when "1001100001110110" => data_out <= rom_array(39030);
		when "1001100001110111" => data_out <= rom_array(39031);
		when "1001100001111000" => data_out <= rom_array(39032);
		when "1001100001111001" => data_out <= rom_array(39033);
		when "1001100001111010" => data_out <= rom_array(39034);
		when "1001100001111011" => data_out <= rom_array(39035);
		when "1001100001111100" => data_out <= rom_array(39036);
		when "1001100001111101" => data_out <= rom_array(39037);
		when "1001100001111110" => data_out <= rom_array(39038);
		when "1001100001111111" => data_out <= rom_array(39039);
		when "1001100010000000" => data_out <= rom_array(39040);
		when "1001100010000001" => data_out <= rom_array(39041);
		when "1001100010000010" => data_out <= rom_array(39042);
		when "1001100010000011" => data_out <= rom_array(39043);
		when "1001100010000100" => data_out <= rom_array(39044);
		when "1001100010000101" => data_out <= rom_array(39045);
		when "1001100010000110" => data_out <= rom_array(39046);
		when "1001100010000111" => data_out <= rom_array(39047);
		when "1001100010001000" => data_out <= rom_array(39048);
		when "1001100010001001" => data_out <= rom_array(39049);
		when "1001100010001010" => data_out <= rom_array(39050);
		when "1001100010001011" => data_out <= rom_array(39051);
		when "1001100010001100" => data_out <= rom_array(39052);
		when "1001100010001101" => data_out <= rom_array(39053);
		when "1001100010001110" => data_out <= rom_array(39054);
		when "1001100010001111" => data_out <= rom_array(39055);
		when "1001100010010000" => data_out <= rom_array(39056);
		when "1001100010010001" => data_out <= rom_array(39057);
		when "1001100010010010" => data_out <= rom_array(39058);
		when "1001100010010011" => data_out <= rom_array(39059);
		when "1001100010010100" => data_out <= rom_array(39060);
		when "1001100010010101" => data_out <= rom_array(39061);
		when "1001100010010110" => data_out <= rom_array(39062);
		when "1001100010010111" => data_out <= rom_array(39063);
		when "1001100010011000" => data_out <= rom_array(39064);
		when "1001100010011001" => data_out <= rom_array(39065);
		when "1001100010011010" => data_out <= rom_array(39066);
		when "1001100010011011" => data_out <= rom_array(39067);
		when "1001100010011100" => data_out <= rom_array(39068);
		when "1001100010011101" => data_out <= rom_array(39069);
		when "1001100010011110" => data_out <= rom_array(39070);
		when "1001100010011111" => data_out <= rom_array(39071);
		when "1001100010100000" => data_out <= rom_array(39072);
		when "1001100010100001" => data_out <= rom_array(39073);
		when "1001100010100010" => data_out <= rom_array(39074);
		when "1001100010100011" => data_out <= rom_array(39075);
		when "1001100010100100" => data_out <= rom_array(39076);
		when "1001100010100101" => data_out <= rom_array(39077);
		when "1001100010100110" => data_out <= rom_array(39078);
		when "1001100010100111" => data_out <= rom_array(39079);
		when "1001100010101000" => data_out <= rom_array(39080);
		when "1001100010101001" => data_out <= rom_array(39081);
		when "1001100010101010" => data_out <= rom_array(39082);
		when "1001100010101011" => data_out <= rom_array(39083);
		when "1001100010101100" => data_out <= rom_array(39084);
		when "1001100010101101" => data_out <= rom_array(39085);
		when "1001100010101110" => data_out <= rom_array(39086);
		when "1001100010101111" => data_out <= rom_array(39087);
		when "1001100010110000" => data_out <= rom_array(39088);
		when "1001100010110001" => data_out <= rom_array(39089);
		when "1001100010110010" => data_out <= rom_array(39090);
		when "1001100010110011" => data_out <= rom_array(39091);
		when "1001100010110100" => data_out <= rom_array(39092);
		when "1001100010110101" => data_out <= rom_array(39093);
		when "1001100010110110" => data_out <= rom_array(39094);
		when "1001100010110111" => data_out <= rom_array(39095);
		when "1001100010111000" => data_out <= rom_array(39096);
		when "1001100010111001" => data_out <= rom_array(39097);
		when "1001100010111010" => data_out <= rom_array(39098);
		when "1001100010111011" => data_out <= rom_array(39099);
		when "1001100010111100" => data_out <= rom_array(39100);
		when "1001100010111101" => data_out <= rom_array(39101);
		when "1001100010111110" => data_out <= rom_array(39102);
		when "1001100010111111" => data_out <= rom_array(39103);
		when "1001100011000000" => data_out <= rom_array(39104);
		when "1001100011000001" => data_out <= rom_array(39105);
		when "1001100011000010" => data_out <= rom_array(39106);
		when "1001100011000011" => data_out <= rom_array(39107);
		when "1001100011000100" => data_out <= rom_array(39108);
		when "1001100011000101" => data_out <= rom_array(39109);
		when "1001100011000110" => data_out <= rom_array(39110);
		when "1001100011000111" => data_out <= rom_array(39111);
		when "1001100011001000" => data_out <= rom_array(39112);
		when "1001100011001001" => data_out <= rom_array(39113);
		when "1001100011001010" => data_out <= rom_array(39114);
		when "1001100011001011" => data_out <= rom_array(39115);
		when "1001100011001100" => data_out <= rom_array(39116);
		when "1001100011001101" => data_out <= rom_array(39117);
		when "1001100011001110" => data_out <= rom_array(39118);
		when "1001100011001111" => data_out <= rom_array(39119);
		when "1001100011010000" => data_out <= rom_array(39120);
		when "1001100011010001" => data_out <= rom_array(39121);
		when "1001100011010010" => data_out <= rom_array(39122);
		when "1001100011010011" => data_out <= rom_array(39123);
		when "1001100011010100" => data_out <= rom_array(39124);
		when "1001100011010101" => data_out <= rom_array(39125);
		when "1001100011010110" => data_out <= rom_array(39126);
		when "1001100011010111" => data_out <= rom_array(39127);
		when "1001100011011000" => data_out <= rom_array(39128);
		when "1001100011011001" => data_out <= rom_array(39129);
		when "1001100011011010" => data_out <= rom_array(39130);
		when "1001100011011011" => data_out <= rom_array(39131);
		when "1001100011011100" => data_out <= rom_array(39132);
		when "1001100011011101" => data_out <= rom_array(39133);
		when "1001100011011110" => data_out <= rom_array(39134);
		when "1001100011011111" => data_out <= rom_array(39135);
		when "1001100011100000" => data_out <= rom_array(39136);
		when "1001100011100001" => data_out <= rom_array(39137);
		when "1001100011100010" => data_out <= rom_array(39138);
		when "1001100011100011" => data_out <= rom_array(39139);
		when "1001100011100100" => data_out <= rom_array(39140);
		when "1001100011100101" => data_out <= rom_array(39141);
		when "1001100011100110" => data_out <= rom_array(39142);
		when "1001100011100111" => data_out <= rom_array(39143);
		when "1001100011101000" => data_out <= rom_array(39144);
		when "1001100011101001" => data_out <= rom_array(39145);
		when "1001100011101010" => data_out <= rom_array(39146);
		when "1001100011101011" => data_out <= rom_array(39147);
		when "1001100011101100" => data_out <= rom_array(39148);
		when "1001100011101101" => data_out <= rom_array(39149);
		when "1001100011101110" => data_out <= rom_array(39150);
		when "1001100011101111" => data_out <= rom_array(39151);
		when "1001100011110000" => data_out <= rom_array(39152);
		when "1001100011110001" => data_out <= rom_array(39153);
		when "1001100011110010" => data_out <= rom_array(39154);
		when "1001100011110011" => data_out <= rom_array(39155);
		when "1001100011110100" => data_out <= rom_array(39156);
		when "1001100011110101" => data_out <= rom_array(39157);
		when "1001100011110110" => data_out <= rom_array(39158);
		when "1001100011110111" => data_out <= rom_array(39159);
		when "1001100011111000" => data_out <= rom_array(39160);
		when "1001100011111001" => data_out <= rom_array(39161);
		when "1001100011111010" => data_out <= rom_array(39162);
		when "1001100011111011" => data_out <= rom_array(39163);
		when "1001100011111100" => data_out <= rom_array(39164);
		when "1001100011111101" => data_out <= rom_array(39165);
		when "1001100011111110" => data_out <= rom_array(39166);
		when "1001100011111111" => data_out <= rom_array(39167);
		when "1001100100000000" => data_out <= rom_array(39168);
		when "1001100100000001" => data_out <= rom_array(39169);
		when "1001100100000010" => data_out <= rom_array(39170);
		when "1001100100000011" => data_out <= rom_array(39171);
		when "1001100100000100" => data_out <= rom_array(39172);
		when "1001100100000101" => data_out <= rom_array(39173);
		when "1001100100000110" => data_out <= rom_array(39174);
		when "1001100100000111" => data_out <= rom_array(39175);
		when "1001100100001000" => data_out <= rom_array(39176);
		when "1001100100001001" => data_out <= rom_array(39177);
		when "1001100100001010" => data_out <= rom_array(39178);
		when "1001100100001011" => data_out <= rom_array(39179);
		when "1001100100001100" => data_out <= rom_array(39180);
		when "1001100100001101" => data_out <= rom_array(39181);
		when "1001100100001110" => data_out <= rom_array(39182);
		when "1001100100001111" => data_out <= rom_array(39183);
		when "1001100100010000" => data_out <= rom_array(39184);
		when "1001100100010001" => data_out <= rom_array(39185);
		when "1001100100010010" => data_out <= rom_array(39186);
		when "1001100100010011" => data_out <= rom_array(39187);
		when "1001100100010100" => data_out <= rom_array(39188);
		when "1001100100010101" => data_out <= rom_array(39189);
		when "1001100100010110" => data_out <= rom_array(39190);
		when "1001100100010111" => data_out <= rom_array(39191);
		when "1001100100011000" => data_out <= rom_array(39192);
		when "1001100100011001" => data_out <= rom_array(39193);
		when "1001100100011010" => data_out <= rom_array(39194);
		when "1001100100011011" => data_out <= rom_array(39195);
		when "1001100100011100" => data_out <= rom_array(39196);
		when "1001100100011101" => data_out <= rom_array(39197);
		when "1001100100011110" => data_out <= rom_array(39198);
		when "1001100100011111" => data_out <= rom_array(39199);
		when "1001100100100000" => data_out <= rom_array(39200);
		when "1001100100100001" => data_out <= rom_array(39201);
		when "1001100100100010" => data_out <= rom_array(39202);
		when "1001100100100011" => data_out <= rom_array(39203);
		when "1001100100100100" => data_out <= rom_array(39204);
		when "1001100100100101" => data_out <= rom_array(39205);
		when "1001100100100110" => data_out <= rom_array(39206);
		when "1001100100100111" => data_out <= rom_array(39207);
		when "1001100100101000" => data_out <= rom_array(39208);
		when "1001100100101001" => data_out <= rom_array(39209);
		when "1001100100101010" => data_out <= rom_array(39210);
		when "1001100100101011" => data_out <= rom_array(39211);
		when "1001100100101100" => data_out <= rom_array(39212);
		when "1001100100101101" => data_out <= rom_array(39213);
		when "1001100100101110" => data_out <= rom_array(39214);
		when "1001100100101111" => data_out <= rom_array(39215);
		when "1001100100110000" => data_out <= rom_array(39216);
		when "1001100100110001" => data_out <= rom_array(39217);
		when "1001100100110010" => data_out <= rom_array(39218);
		when "1001100100110011" => data_out <= rom_array(39219);
		when "1001100100110100" => data_out <= rom_array(39220);
		when "1001100100110101" => data_out <= rom_array(39221);
		when "1001100100110110" => data_out <= rom_array(39222);
		when "1001100100110111" => data_out <= rom_array(39223);
		when "1001100100111000" => data_out <= rom_array(39224);
		when "1001100100111001" => data_out <= rom_array(39225);
		when "1001100100111010" => data_out <= rom_array(39226);
		when "1001100100111011" => data_out <= rom_array(39227);
		when "1001100100111100" => data_out <= rom_array(39228);
		when "1001100100111101" => data_out <= rom_array(39229);
		when "1001100100111110" => data_out <= rom_array(39230);
		when "1001100100111111" => data_out <= rom_array(39231);
		when "1001100101000000" => data_out <= rom_array(39232);
		when "1001100101000001" => data_out <= rom_array(39233);
		when "1001100101000010" => data_out <= rom_array(39234);
		when "1001100101000011" => data_out <= rom_array(39235);
		when "1001100101000100" => data_out <= rom_array(39236);
		when "1001100101000101" => data_out <= rom_array(39237);
		when "1001100101000110" => data_out <= rom_array(39238);
		when "1001100101000111" => data_out <= rom_array(39239);
		when "1001100101001000" => data_out <= rom_array(39240);
		when "1001100101001001" => data_out <= rom_array(39241);
		when "1001100101001010" => data_out <= rom_array(39242);
		when "1001100101001011" => data_out <= rom_array(39243);
		when "1001100101001100" => data_out <= rom_array(39244);
		when "1001100101001101" => data_out <= rom_array(39245);
		when "1001100101001110" => data_out <= rom_array(39246);
		when "1001100101001111" => data_out <= rom_array(39247);
		when "1001100101010000" => data_out <= rom_array(39248);
		when "1001100101010001" => data_out <= rom_array(39249);
		when "1001100101010010" => data_out <= rom_array(39250);
		when "1001100101010011" => data_out <= rom_array(39251);
		when "1001100101010100" => data_out <= rom_array(39252);
		when "1001100101010101" => data_out <= rom_array(39253);
		when "1001100101010110" => data_out <= rom_array(39254);
		when "1001100101010111" => data_out <= rom_array(39255);
		when "1001100101011000" => data_out <= rom_array(39256);
		when "1001100101011001" => data_out <= rom_array(39257);
		when "1001100101011010" => data_out <= rom_array(39258);
		when "1001100101011011" => data_out <= rom_array(39259);
		when "1001100101011100" => data_out <= rom_array(39260);
		when "1001100101011101" => data_out <= rom_array(39261);
		when "1001100101011110" => data_out <= rom_array(39262);
		when "1001100101011111" => data_out <= rom_array(39263);
		when "1001100101100000" => data_out <= rom_array(39264);
		when "1001100101100001" => data_out <= rom_array(39265);
		when "1001100101100010" => data_out <= rom_array(39266);
		when "1001100101100011" => data_out <= rom_array(39267);
		when "1001100101100100" => data_out <= rom_array(39268);
		when "1001100101100101" => data_out <= rom_array(39269);
		when "1001100101100110" => data_out <= rom_array(39270);
		when "1001100101100111" => data_out <= rom_array(39271);
		when "1001100101101000" => data_out <= rom_array(39272);
		when "1001100101101001" => data_out <= rom_array(39273);
		when "1001100101101010" => data_out <= rom_array(39274);
		when "1001100101101011" => data_out <= rom_array(39275);
		when "1001100101101100" => data_out <= rom_array(39276);
		when "1001100101101101" => data_out <= rom_array(39277);
		when "1001100101101110" => data_out <= rom_array(39278);
		when "1001100101101111" => data_out <= rom_array(39279);
		when "1001100101110000" => data_out <= rom_array(39280);
		when "1001100101110001" => data_out <= rom_array(39281);
		when "1001100101110010" => data_out <= rom_array(39282);
		when "1001100101110011" => data_out <= rom_array(39283);
		when "1001100101110100" => data_out <= rom_array(39284);
		when "1001100101110101" => data_out <= rom_array(39285);
		when "1001100101110110" => data_out <= rom_array(39286);
		when "1001100101110111" => data_out <= rom_array(39287);
		when "1001100101111000" => data_out <= rom_array(39288);
		when "1001100101111001" => data_out <= rom_array(39289);
		when "1001100101111010" => data_out <= rom_array(39290);
		when "1001100101111011" => data_out <= rom_array(39291);
		when "1001100101111100" => data_out <= rom_array(39292);
		when "1001100101111101" => data_out <= rom_array(39293);
		when "1001100101111110" => data_out <= rom_array(39294);
		when "1001100101111111" => data_out <= rom_array(39295);
		when "1001100110000000" => data_out <= rom_array(39296);
		when "1001100110000001" => data_out <= rom_array(39297);
		when "1001100110000010" => data_out <= rom_array(39298);
		when "1001100110000011" => data_out <= rom_array(39299);
		when "1001100110000100" => data_out <= rom_array(39300);
		when "1001100110000101" => data_out <= rom_array(39301);
		when "1001100110000110" => data_out <= rom_array(39302);
		when "1001100110000111" => data_out <= rom_array(39303);
		when "1001100110001000" => data_out <= rom_array(39304);
		when "1001100110001001" => data_out <= rom_array(39305);
		when "1001100110001010" => data_out <= rom_array(39306);
		when "1001100110001011" => data_out <= rom_array(39307);
		when "1001100110001100" => data_out <= rom_array(39308);
		when "1001100110001101" => data_out <= rom_array(39309);
		when "1001100110001110" => data_out <= rom_array(39310);
		when "1001100110001111" => data_out <= rom_array(39311);
		when "1001100110010000" => data_out <= rom_array(39312);
		when "1001100110010001" => data_out <= rom_array(39313);
		when "1001100110010010" => data_out <= rom_array(39314);
		when "1001100110010011" => data_out <= rom_array(39315);
		when "1001100110010100" => data_out <= rom_array(39316);
		when "1001100110010101" => data_out <= rom_array(39317);
		when "1001100110010110" => data_out <= rom_array(39318);
		when "1001100110010111" => data_out <= rom_array(39319);
		when "1001100110011000" => data_out <= rom_array(39320);
		when "1001100110011001" => data_out <= rom_array(39321);
		when "1001100110011010" => data_out <= rom_array(39322);
		when "1001100110011011" => data_out <= rom_array(39323);
		when "1001100110011100" => data_out <= rom_array(39324);
		when "1001100110011101" => data_out <= rom_array(39325);
		when "1001100110011110" => data_out <= rom_array(39326);
		when "1001100110011111" => data_out <= rom_array(39327);
		when "1001100110100000" => data_out <= rom_array(39328);
		when "1001100110100001" => data_out <= rom_array(39329);
		when "1001100110100010" => data_out <= rom_array(39330);
		when "1001100110100011" => data_out <= rom_array(39331);
		when "1001100110100100" => data_out <= rom_array(39332);
		when "1001100110100101" => data_out <= rom_array(39333);
		when "1001100110100110" => data_out <= rom_array(39334);
		when "1001100110100111" => data_out <= rom_array(39335);
		when "1001100110101000" => data_out <= rom_array(39336);
		when "1001100110101001" => data_out <= rom_array(39337);
		when "1001100110101010" => data_out <= rom_array(39338);
		when "1001100110101011" => data_out <= rom_array(39339);
		when "1001100110101100" => data_out <= rom_array(39340);
		when "1001100110101101" => data_out <= rom_array(39341);
		when "1001100110101110" => data_out <= rom_array(39342);
		when "1001100110101111" => data_out <= rom_array(39343);
		when "1001100110110000" => data_out <= rom_array(39344);
		when "1001100110110001" => data_out <= rom_array(39345);
		when "1001100110110010" => data_out <= rom_array(39346);
		when "1001100110110011" => data_out <= rom_array(39347);
		when "1001100110110100" => data_out <= rom_array(39348);
		when "1001100110110101" => data_out <= rom_array(39349);
		when "1001100110110110" => data_out <= rom_array(39350);
		when "1001100110110111" => data_out <= rom_array(39351);
		when "1001100110111000" => data_out <= rom_array(39352);
		when "1001100110111001" => data_out <= rom_array(39353);
		when "1001100110111010" => data_out <= rom_array(39354);
		when "1001100110111011" => data_out <= rom_array(39355);
		when "1001100110111100" => data_out <= rom_array(39356);
		when "1001100110111101" => data_out <= rom_array(39357);
		when "1001100110111110" => data_out <= rom_array(39358);
		when "1001100110111111" => data_out <= rom_array(39359);
		when "1001100111000000" => data_out <= rom_array(39360);
		when "1001100111000001" => data_out <= rom_array(39361);
		when "1001100111000010" => data_out <= rom_array(39362);
		when "1001100111000011" => data_out <= rom_array(39363);
		when "1001100111000100" => data_out <= rom_array(39364);
		when "1001100111000101" => data_out <= rom_array(39365);
		when "1001100111000110" => data_out <= rom_array(39366);
		when "1001100111000111" => data_out <= rom_array(39367);
		when "1001100111001000" => data_out <= rom_array(39368);
		when "1001100111001001" => data_out <= rom_array(39369);
		when "1001100111001010" => data_out <= rom_array(39370);
		when "1001100111001011" => data_out <= rom_array(39371);
		when "1001100111001100" => data_out <= rom_array(39372);
		when "1001100111001101" => data_out <= rom_array(39373);
		when "1001100111001110" => data_out <= rom_array(39374);
		when "1001100111001111" => data_out <= rom_array(39375);
		when "1001100111010000" => data_out <= rom_array(39376);
		when "1001100111010001" => data_out <= rom_array(39377);
		when "1001100111010010" => data_out <= rom_array(39378);
		when "1001100111010011" => data_out <= rom_array(39379);
		when "1001100111010100" => data_out <= rom_array(39380);
		when "1001100111010101" => data_out <= rom_array(39381);
		when "1001100111010110" => data_out <= rom_array(39382);
		when "1001100111010111" => data_out <= rom_array(39383);
		when "1001100111011000" => data_out <= rom_array(39384);
		when "1001100111011001" => data_out <= rom_array(39385);
		when "1001100111011010" => data_out <= rom_array(39386);
		when "1001100111011011" => data_out <= rom_array(39387);
		when "1001100111011100" => data_out <= rom_array(39388);
		when "1001100111011101" => data_out <= rom_array(39389);
		when "1001100111011110" => data_out <= rom_array(39390);
		when "1001100111011111" => data_out <= rom_array(39391);
		when "1001100111100000" => data_out <= rom_array(39392);
		when "1001100111100001" => data_out <= rom_array(39393);
		when "1001100111100010" => data_out <= rom_array(39394);
		when "1001100111100011" => data_out <= rom_array(39395);
		when "1001100111100100" => data_out <= rom_array(39396);
		when "1001100111100101" => data_out <= rom_array(39397);
		when "1001100111100110" => data_out <= rom_array(39398);
		when "1001100111100111" => data_out <= rom_array(39399);
		when "1001100111101000" => data_out <= rom_array(39400);
		when "1001100111101001" => data_out <= rom_array(39401);
		when "1001100111101010" => data_out <= rom_array(39402);
		when "1001100111101011" => data_out <= rom_array(39403);
		when "1001100111101100" => data_out <= rom_array(39404);
		when "1001100111101101" => data_out <= rom_array(39405);
		when "1001100111101110" => data_out <= rom_array(39406);
		when "1001100111101111" => data_out <= rom_array(39407);
		when "1001100111110000" => data_out <= rom_array(39408);
		when "1001100111110001" => data_out <= rom_array(39409);
		when "1001100111110010" => data_out <= rom_array(39410);
		when "1001100111110011" => data_out <= rom_array(39411);
		when "1001100111110100" => data_out <= rom_array(39412);
		when "1001100111110101" => data_out <= rom_array(39413);
		when "1001100111110110" => data_out <= rom_array(39414);
		when "1001100111110111" => data_out <= rom_array(39415);
		when "1001100111111000" => data_out <= rom_array(39416);
		when "1001100111111001" => data_out <= rom_array(39417);
		when "1001100111111010" => data_out <= rom_array(39418);
		when "1001100111111011" => data_out <= rom_array(39419);
		when "1001100111111100" => data_out <= rom_array(39420);
		when "1001100111111101" => data_out <= rom_array(39421);
		when "1001100111111110" => data_out <= rom_array(39422);
		when "1001100111111111" => data_out <= rom_array(39423);
		when "1001101000000000" => data_out <= rom_array(39424);
		when "1001101000000001" => data_out <= rom_array(39425);
		when "1001101000000010" => data_out <= rom_array(39426);
		when "1001101000000011" => data_out <= rom_array(39427);
		when "1001101000000100" => data_out <= rom_array(39428);
		when "1001101000000101" => data_out <= rom_array(39429);
		when "1001101000000110" => data_out <= rom_array(39430);
		when "1001101000000111" => data_out <= rom_array(39431);
		when "1001101000001000" => data_out <= rom_array(39432);
		when "1001101000001001" => data_out <= rom_array(39433);
		when "1001101000001010" => data_out <= rom_array(39434);
		when "1001101000001011" => data_out <= rom_array(39435);
		when "1001101000001100" => data_out <= rom_array(39436);
		when "1001101000001101" => data_out <= rom_array(39437);
		when "1001101000001110" => data_out <= rom_array(39438);
		when "1001101000001111" => data_out <= rom_array(39439);
		when "1001101000010000" => data_out <= rom_array(39440);
		when "1001101000010001" => data_out <= rom_array(39441);
		when "1001101000010010" => data_out <= rom_array(39442);
		when "1001101000010011" => data_out <= rom_array(39443);
		when "1001101000010100" => data_out <= rom_array(39444);
		when "1001101000010101" => data_out <= rom_array(39445);
		when "1001101000010110" => data_out <= rom_array(39446);
		when "1001101000010111" => data_out <= rom_array(39447);
		when "1001101000011000" => data_out <= rom_array(39448);
		when "1001101000011001" => data_out <= rom_array(39449);
		when "1001101000011010" => data_out <= rom_array(39450);
		when "1001101000011011" => data_out <= rom_array(39451);
		when "1001101000011100" => data_out <= rom_array(39452);
		when "1001101000011101" => data_out <= rom_array(39453);
		when "1001101000011110" => data_out <= rom_array(39454);
		when "1001101000011111" => data_out <= rom_array(39455);
		when "1001101000100000" => data_out <= rom_array(39456);
		when "1001101000100001" => data_out <= rom_array(39457);
		when "1001101000100010" => data_out <= rom_array(39458);
		when "1001101000100011" => data_out <= rom_array(39459);
		when "1001101000100100" => data_out <= rom_array(39460);
		when "1001101000100101" => data_out <= rom_array(39461);
		when "1001101000100110" => data_out <= rom_array(39462);
		when "1001101000100111" => data_out <= rom_array(39463);
		when "1001101000101000" => data_out <= rom_array(39464);
		when "1001101000101001" => data_out <= rom_array(39465);
		when "1001101000101010" => data_out <= rom_array(39466);
		when "1001101000101011" => data_out <= rom_array(39467);
		when "1001101000101100" => data_out <= rom_array(39468);
		when "1001101000101101" => data_out <= rom_array(39469);
		when "1001101000101110" => data_out <= rom_array(39470);
		when "1001101000101111" => data_out <= rom_array(39471);
		when "1001101000110000" => data_out <= rom_array(39472);
		when "1001101000110001" => data_out <= rom_array(39473);
		when "1001101000110010" => data_out <= rom_array(39474);
		when "1001101000110011" => data_out <= rom_array(39475);
		when "1001101000110100" => data_out <= rom_array(39476);
		when "1001101000110101" => data_out <= rom_array(39477);
		when "1001101000110110" => data_out <= rom_array(39478);
		when "1001101000110111" => data_out <= rom_array(39479);
		when "1001101000111000" => data_out <= rom_array(39480);
		when "1001101000111001" => data_out <= rom_array(39481);
		when "1001101000111010" => data_out <= rom_array(39482);
		when "1001101000111011" => data_out <= rom_array(39483);
		when "1001101000111100" => data_out <= rom_array(39484);
		when "1001101000111101" => data_out <= rom_array(39485);
		when "1001101000111110" => data_out <= rom_array(39486);
		when "1001101000111111" => data_out <= rom_array(39487);
		when "1001101001000000" => data_out <= rom_array(39488);
		when "1001101001000001" => data_out <= rom_array(39489);
		when "1001101001000010" => data_out <= rom_array(39490);
		when "1001101001000011" => data_out <= rom_array(39491);
		when "1001101001000100" => data_out <= rom_array(39492);
		when "1001101001000101" => data_out <= rom_array(39493);
		when "1001101001000110" => data_out <= rom_array(39494);
		when "1001101001000111" => data_out <= rom_array(39495);
		when "1001101001001000" => data_out <= rom_array(39496);
		when "1001101001001001" => data_out <= rom_array(39497);
		when "1001101001001010" => data_out <= rom_array(39498);
		when "1001101001001011" => data_out <= rom_array(39499);
		when "1001101001001100" => data_out <= rom_array(39500);
		when "1001101001001101" => data_out <= rom_array(39501);
		when "1001101001001110" => data_out <= rom_array(39502);
		when "1001101001001111" => data_out <= rom_array(39503);
		when "1001101001010000" => data_out <= rom_array(39504);
		when "1001101001010001" => data_out <= rom_array(39505);
		when "1001101001010010" => data_out <= rom_array(39506);
		when "1001101001010011" => data_out <= rom_array(39507);
		when "1001101001010100" => data_out <= rom_array(39508);
		when "1001101001010101" => data_out <= rom_array(39509);
		when "1001101001010110" => data_out <= rom_array(39510);
		when "1001101001010111" => data_out <= rom_array(39511);
		when "1001101001011000" => data_out <= rom_array(39512);
		when "1001101001011001" => data_out <= rom_array(39513);
		when "1001101001011010" => data_out <= rom_array(39514);
		when "1001101001011011" => data_out <= rom_array(39515);
		when "1001101001011100" => data_out <= rom_array(39516);
		when "1001101001011101" => data_out <= rom_array(39517);
		when "1001101001011110" => data_out <= rom_array(39518);
		when "1001101001011111" => data_out <= rom_array(39519);
		when "1001101001100000" => data_out <= rom_array(39520);
		when "1001101001100001" => data_out <= rom_array(39521);
		when "1001101001100010" => data_out <= rom_array(39522);
		when "1001101001100011" => data_out <= rom_array(39523);
		when "1001101001100100" => data_out <= rom_array(39524);
		when "1001101001100101" => data_out <= rom_array(39525);
		when "1001101001100110" => data_out <= rom_array(39526);
		when "1001101001100111" => data_out <= rom_array(39527);
		when "1001101001101000" => data_out <= rom_array(39528);
		when "1001101001101001" => data_out <= rom_array(39529);
		when "1001101001101010" => data_out <= rom_array(39530);
		when "1001101001101011" => data_out <= rom_array(39531);
		when "1001101001101100" => data_out <= rom_array(39532);
		when "1001101001101101" => data_out <= rom_array(39533);
		when "1001101001101110" => data_out <= rom_array(39534);
		when "1001101001101111" => data_out <= rom_array(39535);
		when "1001101001110000" => data_out <= rom_array(39536);
		when "1001101001110001" => data_out <= rom_array(39537);
		when "1001101001110010" => data_out <= rom_array(39538);
		when "1001101001110011" => data_out <= rom_array(39539);
		when "1001101001110100" => data_out <= rom_array(39540);
		when "1001101001110101" => data_out <= rom_array(39541);
		when "1001101001110110" => data_out <= rom_array(39542);
		when "1001101001110111" => data_out <= rom_array(39543);
		when "1001101001111000" => data_out <= rom_array(39544);
		when "1001101001111001" => data_out <= rom_array(39545);
		when "1001101001111010" => data_out <= rom_array(39546);
		when "1001101001111011" => data_out <= rom_array(39547);
		when "1001101001111100" => data_out <= rom_array(39548);
		when "1001101001111101" => data_out <= rom_array(39549);
		when "1001101001111110" => data_out <= rom_array(39550);
		when "1001101001111111" => data_out <= rom_array(39551);
		when "1001101010000000" => data_out <= rom_array(39552);
		when "1001101010000001" => data_out <= rom_array(39553);
		when "1001101010000010" => data_out <= rom_array(39554);
		when "1001101010000011" => data_out <= rom_array(39555);
		when "1001101010000100" => data_out <= rom_array(39556);
		when "1001101010000101" => data_out <= rom_array(39557);
		when "1001101010000110" => data_out <= rom_array(39558);
		when "1001101010000111" => data_out <= rom_array(39559);
		when "1001101010001000" => data_out <= rom_array(39560);
		when "1001101010001001" => data_out <= rom_array(39561);
		when "1001101010001010" => data_out <= rom_array(39562);
		when "1001101010001011" => data_out <= rom_array(39563);
		when "1001101010001100" => data_out <= rom_array(39564);
		when "1001101010001101" => data_out <= rom_array(39565);
		when "1001101010001110" => data_out <= rom_array(39566);
		when "1001101010001111" => data_out <= rom_array(39567);
		when "1001101010010000" => data_out <= rom_array(39568);
		when "1001101010010001" => data_out <= rom_array(39569);
		when "1001101010010010" => data_out <= rom_array(39570);
		when "1001101010010011" => data_out <= rom_array(39571);
		when "1001101010010100" => data_out <= rom_array(39572);
		when "1001101010010101" => data_out <= rom_array(39573);
		when "1001101010010110" => data_out <= rom_array(39574);
		when "1001101010010111" => data_out <= rom_array(39575);
		when "1001101010011000" => data_out <= rom_array(39576);
		when "1001101010011001" => data_out <= rom_array(39577);
		when "1001101010011010" => data_out <= rom_array(39578);
		when "1001101010011011" => data_out <= rom_array(39579);
		when "1001101010011100" => data_out <= rom_array(39580);
		when "1001101010011101" => data_out <= rom_array(39581);
		when "1001101010011110" => data_out <= rom_array(39582);
		when "1001101010011111" => data_out <= rom_array(39583);
		when "1001101010100000" => data_out <= rom_array(39584);
		when "1001101010100001" => data_out <= rom_array(39585);
		when "1001101010100010" => data_out <= rom_array(39586);
		when "1001101010100011" => data_out <= rom_array(39587);
		when "1001101010100100" => data_out <= rom_array(39588);
		when "1001101010100101" => data_out <= rom_array(39589);
		when "1001101010100110" => data_out <= rom_array(39590);
		when "1001101010100111" => data_out <= rom_array(39591);
		when "1001101010101000" => data_out <= rom_array(39592);
		when "1001101010101001" => data_out <= rom_array(39593);
		when "1001101010101010" => data_out <= rom_array(39594);
		when "1001101010101011" => data_out <= rom_array(39595);
		when "1001101010101100" => data_out <= rom_array(39596);
		when "1001101010101101" => data_out <= rom_array(39597);
		when "1001101010101110" => data_out <= rom_array(39598);
		when "1001101010101111" => data_out <= rom_array(39599);
		when "1001101010110000" => data_out <= rom_array(39600);
		when "1001101010110001" => data_out <= rom_array(39601);
		when "1001101010110010" => data_out <= rom_array(39602);
		when "1001101010110011" => data_out <= rom_array(39603);
		when "1001101010110100" => data_out <= rom_array(39604);
		when "1001101010110101" => data_out <= rom_array(39605);
		when "1001101010110110" => data_out <= rom_array(39606);
		when "1001101010110111" => data_out <= rom_array(39607);
		when "1001101010111000" => data_out <= rom_array(39608);
		when "1001101010111001" => data_out <= rom_array(39609);
		when "1001101010111010" => data_out <= rom_array(39610);
		when "1001101010111011" => data_out <= rom_array(39611);
		when "1001101010111100" => data_out <= rom_array(39612);
		when "1001101010111101" => data_out <= rom_array(39613);
		when "1001101010111110" => data_out <= rom_array(39614);
		when "1001101010111111" => data_out <= rom_array(39615);
		when "1001101011000000" => data_out <= rom_array(39616);
		when "1001101011000001" => data_out <= rom_array(39617);
		when "1001101011000010" => data_out <= rom_array(39618);
		when "1001101011000011" => data_out <= rom_array(39619);
		when "1001101011000100" => data_out <= rom_array(39620);
		when "1001101011000101" => data_out <= rom_array(39621);
		when "1001101011000110" => data_out <= rom_array(39622);
		when "1001101011000111" => data_out <= rom_array(39623);
		when "1001101011001000" => data_out <= rom_array(39624);
		when "1001101011001001" => data_out <= rom_array(39625);
		when "1001101011001010" => data_out <= rom_array(39626);
		when "1001101011001011" => data_out <= rom_array(39627);
		when "1001101011001100" => data_out <= rom_array(39628);
		when "1001101011001101" => data_out <= rom_array(39629);
		when "1001101011001110" => data_out <= rom_array(39630);
		when "1001101011001111" => data_out <= rom_array(39631);
		when "1001101011010000" => data_out <= rom_array(39632);
		when "1001101011010001" => data_out <= rom_array(39633);
		when "1001101011010010" => data_out <= rom_array(39634);
		when "1001101011010011" => data_out <= rom_array(39635);
		when "1001101011010100" => data_out <= rom_array(39636);
		when "1001101011010101" => data_out <= rom_array(39637);
		when "1001101011010110" => data_out <= rom_array(39638);
		when "1001101011010111" => data_out <= rom_array(39639);
		when "1001101011011000" => data_out <= rom_array(39640);
		when "1001101011011001" => data_out <= rom_array(39641);
		when "1001101011011010" => data_out <= rom_array(39642);
		when "1001101011011011" => data_out <= rom_array(39643);
		when "1001101011011100" => data_out <= rom_array(39644);
		when "1001101011011101" => data_out <= rom_array(39645);
		when "1001101011011110" => data_out <= rom_array(39646);
		when "1001101011011111" => data_out <= rom_array(39647);
		when "1001101011100000" => data_out <= rom_array(39648);
		when "1001101011100001" => data_out <= rom_array(39649);
		when "1001101011100010" => data_out <= rom_array(39650);
		when "1001101011100011" => data_out <= rom_array(39651);
		when "1001101011100100" => data_out <= rom_array(39652);
		when "1001101011100101" => data_out <= rom_array(39653);
		when "1001101011100110" => data_out <= rom_array(39654);
		when "1001101011100111" => data_out <= rom_array(39655);
		when "1001101011101000" => data_out <= rom_array(39656);
		when "1001101011101001" => data_out <= rom_array(39657);
		when "1001101011101010" => data_out <= rom_array(39658);
		when "1001101011101011" => data_out <= rom_array(39659);
		when "1001101011101100" => data_out <= rom_array(39660);
		when "1001101011101101" => data_out <= rom_array(39661);
		when "1001101011101110" => data_out <= rom_array(39662);
		when "1001101011101111" => data_out <= rom_array(39663);
		when "1001101011110000" => data_out <= rom_array(39664);
		when "1001101011110001" => data_out <= rom_array(39665);
		when "1001101011110010" => data_out <= rom_array(39666);
		when "1001101011110011" => data_out <= rom_array(39667);
		when "1001101011110100" => data_out <= rom_array(39668);
		when "1001101011110101" => data_out <= rom_array(39669);
		when "1001101011110110" => data_out <= rom_array(39670);
		when "1001101011110111" => data_out <= rom_array(39671);
		when "1001101011111000" => data_out <= rom_array(39672);
		when "1001101011111001" => data_out <= rom_array(39673);
		when "1001101011111010" => data_out <= rom_array(39674);
		when "1001101011111011" => data_out <= rom_array(39675);
		when "1001101011111100" => data_out <= rom_array(39676);
		when "1001101011111101" => data_out <= rom_array(39677);
		when "1001101011111110" => data_out <= rom_array(39678);
		when "1001101011111111" => data_out <= rom_array(39679);
		when "1001101100000000" => data_out <= rom_array(39680);
		when "1001101100000001" => data_out <= rom_array(39681);
		when "1001101100000010" => data_out <= rom_array(39682);
		when "1001101100000011" => data_out <= rom_array(39683);
		when "1001101100000100" => data_out <= rom_array(39684);
		when "1001101100000101" => data_out <= rom_array(39685);
		when "1001101100000110" => data_out <= rom_array(39686);
		when "1001101100000111" => data_out <= rom_array(39687);
		when "1001101100001000" => data_out <= rom_array(39688);
		when "1001101100001001" => data_out <= rom_array(39689);
		when "1001101100001010" => data_out <= rom_array(39690);
		when "1001101100001011" => data_out <= rom_array(39691);
		when "1001101100001100" => data_out <= rom_array(39692);
		when "1001101100001101" => data_out <= rom_array(39693);
		when "1001101100001110" => data_out <= rom_array(39694);
		when "1001101100001111" => data_out <= rom_array(39695);
		when "1001101100010000" => data_out <= rom_array(39696);
		when "1001101100010001" => data_out <= rom_array(39697);
		when "1001101100010010" => data_out <= rom_array(39698);
		when "1001101100010011" => data_out <= rom_array(39699);
		when "1001101100010100" => data_out <= rom_array(39700);
		when "1001101100010101" => data_out <= rom_array(39701);
		when "1001101100010110" => data_out <= rom_array(39702);
		when "1001101100010111" => data_out <= rom_array(39703);
		when "1001101100011000" => data_out <= rom_array(39704);
		when "1001101100011001" => data_out <= rom_array(39705);
		when "1001101100011010" => data_out <= rom_array(39706);
		when "1001101100011011" => data_out <= rom_array(39707);
		when "1001101100011100" => data_out <= rom_array(39708);
		when "1001101100011101" => data_out <= rom_array(39709);
		when "1001101100011110" => data_out <= rom_array(39710);
		when "1001101100011111" => data_out <= rom_array(39711);
		when "1001101100100000" => data_out <= rom_array(39712);
		when "1001101100100001" => data_out <= rom_array(39713);
		when "1001101100100010" => data_out <= rom_array(39714);
		when "1001101100100011" => data_out <= rom_array(39715);
		when "1001101100100100" => data_out <= rom_array(39716);
		when "1001101100100101" => data_out <= rom_array(39717);
		when "1001101100100110" => data_out <= rom_array(39718);
		when "1001101100100111" => data_out <= rom_array(39719);
		when "1001101100101000" => data_out <= rom_array(39720);
		when "1001101100101001" => data_out <= rom_array(39721);
		when "1001101100101010" => data_out <= rom_array(39722);
		when "1001101100101011" => data_out <= rom_array(39723);
		when "1001101100101100" => data_out <= rom_array(39724);
		when "1001101100101101" => data_out <= rom_array(39725);
		when "1001101100101110" => data_out <= rom_array(39726);
		when "1001101100101111" => data_out <= rom_array(39727);
		when "1001101100110000" => data_out <= rom_array(39728);
		when "1001101100110001" => data_out <= rom_array(39729);
		when "1001101100110010" => data_out <= rom_array(39730);
		when "1001101100110011" => data_out <= rom_array(39731);
		when "1001101100110100" => data_out <= rom_array(39732);
		when "1001101100110101" => data_out <= rom_array(39733);
		when "1001101100110110" => data_out <= rom_array(39734);
		when "1001101100110111" => data_out <= rom_array(39735);
		when "1001101100111000" => data_out <= rom_array(39736);
		when "1001101100111001" => data_out <= rom_array(39737);
		when "1001101100111010" => data_out <= rom_array(39738);
		when "1001101100111011" => data_out <= rom_array(39739);
		when "1001101100111100" => data_out <= rom_array(39740);
		when "1001101100111101" => data_out <= rom_array(39741);
		when "1001101100111110" => data_out <= rom_array(39742);
		when "1001101100111111" => data_out <= rom_array(39743);
		when "1001101101000000" => data_out <= rom_array(39744);
		when "1001101101000001" => data_out <= rom_array(39745);
		when "1001101101000010" => data_out <= rom_array(39746);
		when "1001101101000011" => data_out <= rom_array(39747);
		when "1001101101000100" => data_out <= rom_array(39748);
		when "1001101101000101" => data_out <= rom_array(39749);
		when "1001101101000110" => data_out <= rom_array(39750);
		when "1001101101000111" => data_out <= rom_array(39751);
		when "1001101101001000" => data_out <= rom_array(39752);
		when "1001101101001001" => data_out <= rom_array(39753);
		when "1001101101001010" => data_out <= rom_array(39754);
		when "1001101101001011" => data_out <= rom_array(39755);
		when "1001101101001100" => data_out <= rom_array(39756);
		when "1001101101001101" => data_out <= rom_array(39757);
		when "1001101101001110" => data_out <= rom_array(39758);
		when "1001101101001111" => data_out <= rom_array(39759);
		when "1001101101010000" => data_out <= rom_array(39760);
		when "1001101101010001" => data_out <= rom_array(39761);
		when "1001101101010010" => data_out <= rom_array(39762);
		when "1001101101010011" => data_out <= rom_array(39763);
		when "1001101101010100" => data_out <= rom_array(39764);
		when "1001101101010101" => data_out <= rom_array(39765);
		when "1001101101010110" => data_out <= rom_array(39766);
		when "1001101101010111" => data_out <= rom_array(39767);
		when "1001101101011000" => data_out <= rom_array(39768);
		when "1001101101011001" => data_out <= rom_array(39769);
		when "1001101101011010" => data_out <= rom_array(39770);
		when "1001101101011011" => data_out <= rom_array(39771);
		when "1001101101011100" => data_out <= rom_array(39772);
		when "1001101101011101" => data_out <= rom_array(39773);
		when "1001101101011110" => data_out <= rom_array(39774);
		when "1001101101011111" => data_out <= rom_array(39775);
		when "1001101101100000" => data_out <= rom_array(39776);
		when "1001101101100001" => data_out <= rom_array(39777);
		when "1001101101100010" => data_out <= rom_array(39778);
		when "1001101101100011" => data_out <= rom_array(39779);
		when "1001101101100100" => data_out <= rom_array(39780);
		when "1001101101100101" => data_out <= rom_array(39781);
		when "1001101101100110" => data_out <= rom_array(39782);
		when "1001101101100111" => data_out <= rom_array(39783);
		when "1001101101101000" => data_out <= rom_array(39784);
		when "1001101101101001" => data_out <= rom_array(39785);
		when "1001101101101010" => data_out <= rom_array(39786);
		when "1001101101101011" => data_out <= rom_array(39787);
		when "1001101101101100" => data_out <= rom_array(39788);
		when "1001101101101101" => data_out <= rom_array(39789);
		when "1001101101101110" => data_out <= rom_array(39790);
		when "1001101101101111" => data_out <= rom_array(39791);
		when "1001101101110000" => data_out <= rom_array(39792);
		when "1001101101110001" => data_out <= rom_array(39793);
		when "1001101101110010" => data_out <= rom_array(39794);
		when "1001101101110011" => data_out <= rom_array(39795);
		when "1001101101110100" => data_out <= rom_array(39796);
		when "1001101101110101" => data_out <= rom_array(39797);
		when "1001101101110110" => data_out <= rom_array(39798);
		when "1001101101110111" => data_out <= rom_array(39799);
		when "1001101101111000" => data_out <= rom_array(39800);
		when "1001101101111001" => data_out <= rom_array(39801);
		when "1001101101111010" => data_out <= rom_array(39802);
		when "1001101101111011" => data_out <= rom_array(39803);
		when "1001101101111100" => data_out <= rom_array(39804);
		when "1001101101111101" => data_out <= rom_array(39805);
		when "1001101101111110" => data_out <= rom_array(39806);
		when "1001101101111111" => data_out <= rom_array(39807);
		when "1001101110000000" => data_out <= rom_array(39808);
		when "1001101110000001" => data_out <= rom_array(39809);
		when "1001101110000010" => data_out <= rom_array(39810);
		when "1001101110000011" => data_out <= rom_array(39811);
		when "1001101110000100" => data_out <= rom_array(39812);
		when "1001101110000101" => data_out <= rom_array(39813);
		when "1001101110000110" => data_out <= rom_array(39814);
		when "1001101110000111" => data_out <= rom_array(39815);
		when "1001101110001000" => data_out <= rom_array(39816);
		when "1001101110001001" => data_out <= rom_array(39817);
		when "1001101110001010" => data_out <= rom_array(39818);
		when "1001101110001011" => data_out <= rom_array(39819);
		when "1001101110001100" => data_out <= rom_array(39820);
		when "1001101110001101" => data_out <= rom_array(39821);
		when "1001101110001110" => data_out <= rom_array(39822);
		when "1001101110001111" => data_out <= rom_array(39823);
		when "1001101110010000" => data_out <= rom_array(39824);
		when "1001101110010001" => data_out <= rom_array(39825);
		when "1001101110010010" => data_out <= rom_array(39826);
		when "1001101110010011" => data_out <= rom_array(39827);
		when "1001101110010100" => data_out <= rom_array(39828);
		when "1001101110010101" => data_out <= rom_array(39829);
		when "1001101110010110" => data_out <= rom_array(39830);
		when "1001101110010111" => data_out <= rom_array(39831);
		when "1001101110011000" => data_out <= rom_array(39832);
		when "1001101110011001" => data_out <= rom_array(39833);
		when "1001101110011010" => data_out <= rom_array(39834);
		when "1001101110011011" => data_out <= rom_array(39835);
		when "1001101110011100" => data_out <= rom_array(39836);
		when "1001101110011101" => data_out <= rom_array(39837);
		when "1001101110011110" => data_out <= rom_array(39838);
		when "1001101110011111" => data_out <= rom_array(39839);
		when "1001101110100000" => data_out <= rom_array(39840);
		when "1001101110100001" => data_out <= rom_array(39841);
		when "1001101110100010" => data_out <= rom_array(39842);
		when "1001101110100011" => data_out <= rom_array(39843);
		when "1001101110100100" => data_out <= rom_array(39844);
		when "1001101110100101" => data_out <= rom_array(39845);
		when "1001101110100110" => data_out <= rom_array(39846);
		when "1001101110100111" => data_out <= rom_array(39847);
		when "1001101110101000" => data_out <= rom_array(39848);
		when "1001101110101001" => data_out <= rom_array(39849);
		when "1001101110101010" => data_out <= rom_array(39850);
		when "1001101110101011" => data_out <= rom_array(39851);
		when "1001101110101100" => data_out <= rom_array(39852);
		when "1001101110101101" => data_out <= rom_array(39853);
		when "1001101110101110" => data_out <= rom_array(39854);
		when "1001101110101111" => data_out <= rom_array(39855);
		when "1001101110110000" => data_out <= rom_array(39856);
		when "1001101110110001" => data_out <= rom_array(39857);
		when "1001101110110010" => data_out <= rom_array(39858);
		when "1001101110110011" => data_out <= rom_array(39859);
		when "1001101110110100" => data_out <= rom_array(39860);
		when "1001101110110101" => data_out <= rom_array(39861);
		when "1001101110110110" => data_out <= rom_array(39862);
		when "1001101110110111" => data_out <= rom_array(39863);
		when "1001101110111000" => data_out <= rom_array(39864);
		when "1001101110111001" => data_out <= rom_array(39865);
		when "1001101110111010" => data_out <= rom_array(39866);
		when "1001101110111011" => data_out <= rom_array(39867);
		when "1001101110111100" => data_out <= rom_array(39868);
		when "1001101110111101" => data_out <= rom_array(39869);
		when "1001101110111110" => data_out <= rom_array(39870);
		when "1001101110111111" => data_out <= rom_array(39871);
		when "1001101111000000" => data_out <= rom_array(39872);
		when "1001101111000001" => data_out <= rom_array(39873);
		when "1001101111000010" => data_out <= rom_array(39874);
		when "1001101111000011" => data_out <= rom_array(39875);
		when "1001101111000100" => data_out <= rom_array(39876);
		when "1001101111000101" => data_out <= rom_array(39877);
		when "1001101111000110" => data_out <= rom_array(39878);
		when "1001101111000111" => data_out <= rom_array(39879);
		when "1001101111001000" => data_out <= rom_array(39880);
		when "1001101111001001" => data_out <= rom_array(39881);
		when "1001101111001010" => data_out <= rom_array(39882);
		when "1001101111001011" => data_out <= rom_array(39883);
		when "1001101111001100" => data_out <= rom_array(39884);
		when "1001101111001101" => data_out <= rom_array(39885);
		when "1001101111001110" => data_out <= rom_array(39886);
		when "1001101111001111" => data_out <= rom_array(39887);
		when "1001101111010000" => data_out <= rom_array(39888);
		when "1001101111010001" => data_out <= rom_array(39889);
		when "1001101111010010" => data_out <= rom_array(39890);
		when "1001101111010011" => data_out <= rom_array(39891);
		when "1001101111010100" => data_out <= rom_array(39892);
		when "1001101111010101" => data_out <= rom_array(39893);
		when "1001101111010110" => data_out <= rom_array(39894);
		when "1001101111010111" => data_out <= rom_array(39895);
		when "1001101111011000" => data_out <= rom_array(39896);
		when "1001101111011001" => data_out <= rom_array(39897);
		when "1001101111011010" => data_out <= rom_array(39898);
		when "1001101111011011" => data_out <= rom_array(39899);
		when "1001101111011100" => data_out <= rom_array(39900);
		when "1001101111011101" => data_out <= rom_array(39901);
		when "1001101111011110" => data_out <= rom_array(39902);
		when "1001101111011111" => data_out <= rom_array(39903);
		when "1001101111100000" => data_out <= rom_array(39904);
		when "1001101111100001" => data_out <= rom_array(39905);
		when "1001101111100010" => data_out <= rom_array(39906);
		when "1001101111100011" => data_out <= rom_array(39907);
		when "1001101111100100" => data_out <= rom_array(39908);
		when "1001101111100101" => data_out <= rom_array(39909);
		when "1001101111100110" => data_out <= rom_array(39910);
		when "1001101111100111" => data_out <= rom_array(39911);
		when "1001101111101000" => data_out <= rom_array(39912);
		when "1001101111101001" => data_out <= rom_array(39913);
		when "1001101111101010" => data_out <= rom_array(39914);
		when "1001101111101011" => data_out <= rom_array(39915);
		when "1001101111101100" => data_out <= rom_array(39916);
		when "1001101111101101" => data_out <= rom_array(39917);
		when "1001101111101110" => data_out <= rom_array(39918);
		when "1001101111101111" => data_out <= rom_array(39919);
		when "1001101111110000" => data_out <= rom_array(39920);
		when "1001101111110001" => data_out <= rom_array(39921);
		when "1001101111110010" => data_out <= rom_array(39922);
		when "1001101111110011" => data_out <= rom_array(39923);
		when "1001101111110100" => data_out <= rom_array(39924);
		when "1001101111110101" => data_out <= rom_array(39925);
		when "1001101111110110" => data_out <= rom_array(39926);
		when "1001101111110111" => data_out <= rom_array(39927);
		when "1001101111111000" => data_out <= rom_array(39928);
		when "1001101111111001" => data_out <= rom_array(39929);
		when "1001101111111010" => data_out <= rom_array(39930);
		when "1001101111111011" => data_out <= rom_array(39931);
		when "1001101111111100" => data_out <= rom_array(39932);
		when "1001101111111101" => data_out <= rom_array(39933);
		when "1001101111111110" => data_out <= rom_array(39934);
		when "1001101111111111" => data_out <= rom_array(39935);
		when "1001110000000000" => data_out <= rom_array(39936);
		when "1001110000000001" => data_out <= rom_array(39937);
		when "1001110000000010" => data_out <= rom_array(39938);
		when "1001110000000011" => data_out <= rom_array(39939);
		when "1001110000000100" => data_out <= rom_array(39940);
		when "1001110000000101" => data_out <= rom_array(39941);
		when "1001110000000110" => data_out <= rom_array(39942);
		when "1001110000000111" => data_out <= rom_array(39943);
		when "1001110000001000" => data_out <= rom_array(39944);
		when "1001110000001001" => data_out <= rom_array(39945);
		when "1001110000001010" => data_out <= rom_array(39946);
		when "1001110000001011" => data_out <= rom_array(39947);
		when "1001110000001100" => data_out <= rom_array(39948);
		when "1001110000001101" => data_out <= rom_array(39949);
		when "1001110000001110" => data_out <= rom_array(39950);
		when "1001110000001111" => data_out <= rom_array(39951);
		when "1001110000010000" => data_out <= rom_array(39952);
		when "1001110000010001" => data_out <= rom_array(39953);
		when "1001110000010010" => data_out <= rom_array(39954);
		when "1001110000010011" => data_out <= rom_array(39955);
		when "1001110000010100" => data_out <= rom_array(39956);
		when "1001110000010101" => data_out <= rom_array(39957);
		when "1001110000010110" => data_out <= rom_array(39958);
		when "1001110000010111" => data_out <= rom_array(39959);
		when "1001110000011000" => data_out <= rom_array(39960);
		when "1001110000011001" => data_out <= rom_array(39961);
		when "1001110000011010" => data_out <= rom_array(39962);
		when "1001110000011011" => data_out <= rom_array(39963);
		when "1001110000011100" => data_out <= rom_array(39964);
		when "1001110000011101" => data_out <= rom_array(39965);
		when "1001110000011110" => data_out <= rom_array(39966);
		when "1001110000011111" => data_out <= rom_array(39967);
		when "1001110000100000" => data_out <= rom_array(39968);
		when "1001110000100001" => data_out <= rom_array(39969);
		when "1001110000100010" => data_out <= rom_array(39970);
		when "1001110000100011" => data_out <= rom_array(39971);
		when "1001110000100100" => data_out <= rom_array(39972);
		when "1001110000100101" => data_out <= rom_array(39973);
		when "1001110000100110" => data_out <= rom_array(39974);
		when "1001110000100111" => data_out <= rom_array(39975);
		when "1001110000101000" => data_out <= rom_array(39976);
		when "1001110000101001" => data_out <= rom_array(39977);
		when "1001110000101010" => data_out <= rom_array(39978);
		when "1001110000101011" => data_out <= rom_array(39979);
		when "1001110000101100" => data_out <= rom_array(39980);
		when "1001110000101101" => data_out <= rom_array(39981);
		when "1001110000101110" => data_out <= rom_array(39982);
		when "1001110000101111" => data_out <= rom_array(39983);
		when "1001110000110000" => data_out <= rom_array(39984);
		when "1001110000110001" => data_out <= rom_array(39985);
		when "1001110000110010" => data_out <= rom_array(39986);
		when "1001110000110011" => data_out <= rom_array(39987);
		when "1001110000110100" => data_out <= rom_array(39988);
		when "1001110000110101" => data_out <= rom_array(39989);
		when "1001110000110110" => data_out <= rom_array(39990);
		when "1001110000110111" => data_out <= rom_array(39991);
		when "1001110000111000" => data_out <= rom_array(39992);
		when "1001110000111001" => data_out <= rom_array(39993);
		when "1001110000111010" => data_out <= rom_array(39994);
		when "1001110000111011" => data_out <= rom_array(39995);
		when "1001110000111100" => data_out <= rom_array(39996);
		when "1001110000111101" => data_out <= rom_array(39997);
		when "1001110000111110" => data_out <= rom_array(39998);
		when "1001110000111111" => data_out <= rom_array(39999);
		when "1001110001000000" => data_out <= rom_array(40000);
		when "1001110001000001" => data_out <= rom_array(40001);
		when "1001110001000010" => data_out <= rom_array(40002);
		when "1001110001000011" => data_out <= rom_array(40003);
		when "1001110001000100" => data_out <= rom_array(40004);
		when "1001110001000101" => data_out <= rom_array(40005);
		when "1001110001000110" => data_out <= rom_array(40006);
		when "1001110001000111" => data_out <= rom_array(40007);
		when "1001110001001000" => data_out <= rom_array(40008);
		when "1001110001001001" => data_out <= rom_array(40009);
		when "1001110001001010" => data_out <= rom_array(40010);
		when "1001110001001011" => data_out <= rom_array(40011);
		when "1001110001001100" => data_out <= rom_array(40012);
		when "1001110001001101" => data_out <= rom_array(40013);
		when "1001110001001110" => data_out <= rom_array(40014);
		when "1001110001001111" => data_out <= rom_array(40015);
		when "1001110001010000" => data_out <= rom_array(40016);
		when "1001110001010001" => data_out <= rom_array(40017);
		when "1001110001010010" => data_out <= rom_array(40018);
		when "1001110001010011" => data_out <= rom_array(40019);
		when "1001110001010100" => data_out <= rom_array(40020);
		when "1001110001010101" => data_out <= rom_array(40021);
		when "1001110001010110" => data_out <= rom_array(40022);
		when "1001110001010111" => data_out <= rom_array(40023);
		when "1001110001011000" => data_out <= rom_array(40024);
		when "1001110001011001" => data_out <= rom_array(40025);
		when "1001110001011010" => data_out <= rom_array(40026);
		when "1001110001011011" => data_out <= rom_array(40027);
		when "1001110001011100" => data_out <= rom_array(40028);
		when "1001110001011101" => data_out <= rom_array(40029);
		when "1001110001011110" => data_out <= rom_array(40030);
		when "1001110001011111" => data_out <= rom_array(40031);
		when "1001110001100000" => data_out <= rom_array(40032);
		when "1001110001100001" => data_out <= rom_array(40033);
		when "1001110001100010" => data_out <= rom_array(40034);
		when "1001110001100011" => data_out <= rom_array(40035);
		when "1001110001100100" => data_out <= rom_array(40036);
		when "1001110001100101" => data_out <= rom_array(40037);
		when "1001110001100110" => data_out <= rom_array(40038);
		when "1001110001100111" => data_out <= rom_array(40039);
		when "1001110001101000" => data_out <= rom_array(40040);
		when "1001110001101001" => data_out <= rom_array(40041);
		when "1001110001101010" => data_out <= rom_array(40042);
		when "1001110001101011" => data_out <= rom_array(40043);
		when "1001110001101100" => data_out <= rom_array(40044);
		when "1001110001101101" => data_out <= rom_array(40045);
		when "1001110001101110" => data_out <= rom_array(40046);
		when "1001110001101111" => data_out <= rom_array(40047);
		when "1001110001110000" => data_out <= rom_array(40048);
		when "1001110001110001" => data_out <= rom_array(40049);
		when "1001110001110010" => data_out <= rom_array(40050);
		when "1001110001110011" => data_out <= rom_array(40051);
		when "1001110001110100" => data_out <= rom_array(40052);
		when "1001110001110101" => data_out <= rom_array(40053);
		when "1001110001110110" => data_out <= rom_array(40054);
		when "1001110001110111" => data_out <= rom_array(40055);
		when "1001110001111000" => data_out <= rom_array(40056);
		when "1001110001111001" => data_out <= rom_array(40057);
		when "1001110001111010" => data_out <= rom_array(40058);
		when "1001110001111011" => data_out <= rom_array(40059);
		when "1001110001111100" => data_out <= rom_array(40060);
		when "1001110001111101" => data_out <= rom_array(40061);
		when "1001110001111110" => data_out <= rom_array(40062);
		when "1001110001111111" => data_out <= rom_array(40063);
		when "1001110010000000" => data_out <= rom_array(40064);
		when "1001110010000001" => data_out <= rom_array(40065);
		when "1001110010000010" => data_out <= rom_array(40066);
		when "1001110010000011" => data_out <= rom_array(40067);
		when "1001110010000100" => data_out <= rom_array(40068);
		when "1001110010000101" => data_out <= rom_array(40069);
		when "1001110010000110" => data_out <= rom_array(40070);
		when "1001110010000111" => data_out <= rom_array(40071);
		when "1001110010001000" => data_out <= rom_array(40072);
		when "1001110010001001" => data_out <= rom_array(40073);
		when "1001110010001010" => data_out <= rom_array(40074);
		when "1001110010001011" => data_out <= rom_array(40075);
		when "1001110010001100" => data_out <= rom_array(40076);
		when "1001110010001101" => data_out <= rom_array(40077);
		when "1001110010001110" => data_out <= rom_array(40078);
		when "1001110010001111" => data_out <= rom_array(40079);
		when "1001110010010000" => data_out <= rom_array(40080);
		when "1001110010010001" => data_out <= rom_array(40081);
		when "1001110010010010" => data_out <= rom_array(40082);
		when "1001110010010011" => data_out <= rom_array(40083);
		when "1001110010010100" => data_out <= rom_array(40084);
		when "1001110010010101" => data_out <= rom_array(40085);
		when "1001110010010110" => data_out <= rom_array(40086);
		when "1001110010010111" => data_out <= rom_array(40087);
		when "1001110010011000" => data_out <= rom_array(40088);
		when "1001110010011001" => data_out <= rom_array(40089);
		when "1001110010011010" => data_out <= rom_array(40090);
		when "1001110010011011" => data_out <= rom_array(40091);
		when "1001110010011100" => data_out <= rom_array(40092);
		when "1001110010011101" => data_out <= rom_array(40093);
		when "1001110010011110" => data_out <= rom_array(40094);
		when "1001110010011111" => data_out <= rom_array(40095);
		when "1001110010100000" => data_out <= rom_array(40096);
		when "1001110010100001" => data_out <= rom_array(40097);
		when "1001110010100010" => data_out <= rom_array(40098);
		when "1001110010100011" => data_out <= rom_array(40099);
		when "1001110010100100" => data_out <= rom_array(40100);
		when "1001110010100101" => data_out <= rom_array(40101);
		when "1001110010100110" => data_out <= rom_array(40102);
		when "1001110010100111" => data_out <= rom_array(40103);
		when "1001110010101000" => data_out <= rom_array(40104);
		when "1001110010101001" => data_out <= rom_array(40105);
		when "1001110010101010" => data_out <= rom_array(40106);
		when "1001110010101011" => data_out <= rom_array(40107);
		when "1001110010101100" => data_out <= rom_array(40108);
		when "1001110010101101" => data_out <= rom_array(40109);
		when "1001110010101110" => data_out <= rom_array(40110);
		when "1001110010101111" => data_out <= rom_array(40111);
		when "1001110010110000" => data_out <= rom_array(40112);
		when "1001110010110001" => data_out <= rom_array(40113);
		when "1001110010110010" => data_out <= rom_array(40114);
		when "1001110010110011" => data_out <= rom_array(40115);
		when "1001110010110100" => data_out <= rom_array(40116);
		when "1001110010110101" => data_out <= rom_array(40117);
		when "1001110010110110" => data_out <= rom_array(40118);
		when "1001110010110111" => data_out <= rom_array(40119);
		when "1001110010111000" => data_out <= rom_array(40120);
		when "1001110010111001" => data_out <= rom_array(40121);
		when "1001110010111010" => data_out <= rom_array(40122);
		when "1001110010111011" => data_out <= rom_array(40123);
		when "1001110010111100" => data_out <= rom_array(40124);
		when "1001110010111101" => data_out <= rom_array(40125);
		when "1001110010111110" => data_out <= rom_array(40126);
		when "1001110010111111" => data_out <= rom_array(40127);
		when "1001110011000000" => data_out <= rom_array(40128);
		when "1001110011000001" => data_out <= rom_array(40129);
		when "1001110011000010" => data_out <= rom_array(40130);
		when "1001110011000011" => data_out <= rom_array(40131);
		when "1001110011000100" => data_out <= rom_array(40132);
		when "1001110011000101" => data_out <= rom_array(40133);
		when "1001110011000110" => data_out <= rom_array(40134);
		when "1001110011000111" => data_out <= rom_array(40135);
		when "1001110011001000" => data_out <= rom_array(40136);
		when "1001110011001001" => data_out <= rom_array(40137);
		when "1001110011001010" => data_out <= rom_array(40138);
		when "1001110011001011" => data_out <= rom_array(40139);
		when "1001110011001100" => data_out <= rom_array(40140);
		when "1001110011001101" => data_out <= rom_array(40141);
		when "1001110011001110" => data_out <= rom_array(40142);
		when "1001110011001111" => data_out <= rom_array(40143);
		when "1001110011010000" => data_out <= rom_array(40144);
		when "1001110011010001" => data_out <= rom_array(40145);
		when "1001110011010010" => data_out <= rom_array(40146);
		when "1001110011010011" => data_out <= rom_array(40147);
		when "1001110011010100" => data_out <= rom_array(40148);
		when "1001110011010101" => data_out <= rom_array(40149);
		when "1001110011010110" => data_out <= rom_array(40150);
		when "1001110011010111" => data_out <= rom_array(40151);
		when "1001110011011000" => data_out <= rom_array(40152);
		when "1001110011011001" => data_out <= rom_array(40153);
		when "1001110011011010" => data_out <= rom_array(40154);
		when "1001110011011011" => data_out <= rom_array(40155);
		when "1001110011011100" => data_out <= rom_array(40156);
		when "1001110011011101" => data_out <= rom_array(40157);
		when "1001110011011110" => data_out <= rom_array(40158);
		when "1001110011011111" => data_out <= rom_array(40159);
		when "1001110011100000" => data_out <= rom_array(40160);
		when "1001110011100001" => data_out <= rom_array(40161);
		when "1001110011100010" => data_out <= rom_array(40162);
		when "1001110011100011" => data_out <= rom_array(40163);
		when "1001110011100100" => data_out <= rom_array(40164);
		when "1001110011100101" => data_out <= rom_array(40165);
		when "1001110011100110" => data_out <= rom_array(40166);
		when "1001110011100111" => data_out <= rom_array(40167);
		when "1001110011101000" => data_out <= rom_array(40168);
		when "1001110011101001" => data_out <= rom_array(40169);
		when "1001110011101010" => data_out <= rom_array(40170);
		when "1001110011101011" => data_out <= rom_array(40171);
		when "1001110011101100" => data_out <= rom_array(40172);
		when "1001110011101101" => data_out <= rom_array(40173);
		when "1001110011101110" => data_out <= rom_array(40174);
		when "1001110011101111" => data_out <= rom_array(40175);
		when "1001110011110000" => data_out <= rom_array(40176);
		when "1001110011110001" => data_out <= rom_array(40177);
		when "1001110011110010" => data_out <= rom_array(40178);
		when "1001110011110011" => data_out <= rom_array(40179);
		when "1001110011110100" => data_out <= rom_array(40180);
		when "1001110011110101" => data_out <= rom_array(40181);
		when "1001110011110110" => data_out <= rom_array(40182);
		when "1001110011110111" => data_out <= rom_array(40183);
		when "1001110011111000" => data_out <= rom_array(40184);
		when "1001110011111001" => data_out <= rom_array(40185);
		when "1001110011111010" => data_out <= rom_array(40186);
		when "1001110011111011" => data_out <= rom_array(40187);
		when "1001110011111100" => data_out <= rom_array(40188);
		when "1001110011111101" => data_out <= rom_array(40189);
		when "1001110011111110" => data_out <= rom_array(40190);
		when "1001110011111111" => data_out <= rom_array(40191);
		when "1001110100000000" => data_out <= rom_array(40192);
		when "1001110100000001" => data_out <= rom_array(40193);
		when "1001110100000010" => data_out <= rom_array(40194);
		when "1001110100000011" => data_out <= rom_array(40195);
		when "1001110100000100" => data_out <= rom_array(40196);
		when "1001110100000101" => data_out <= rom_array(40197);
		when "1001110100000110" => data_out <= rom_array(40198);
		when "1001110100000111" => data_out <= rom_array(40199);
		when "1001110100001000" => data_out <= rom_array(40200);
		when "1001110100001001" => data_out <= rom_array(40201);
		when "1001110100001010" => data_out <= rom_array(40202);
		when "1001110100001011" => data_out <= rom_array(40203);
		when "1001110100001100" => data_out <= rom_array(40204);
		when "1001110100001101" => data_out <= rom_array(40205);
		when "1001110100001110" => data_out <= rom_array(40206);
		when "1001110100001111" => data_out <= rom_array(40207);
		when "1001110100010000" => data_out <= rom_array(40208);
		when "1001110100010001" => data_out <= rom_array(40209);
		when "1001110100010010" => data_out <= rom_array(40210);
		when "1001110100010011" => data_out <= rom_array(40211);
		when "1001110100010100" => data_out <= rom_array(40212);
		when "1001110100010101" => data_out <= rom_array(40213);
		when "1001110100010110" => data_out <= rom_array(40214);
		when "1001110100010111" => data_out <= rom_array(40215);
		when "1001110100011000" => data_out <= rom_array(40216);
		when "1001110100011001" => data_out <= rom_array(40217);
		when "1001110100011010" => data_out <= rom_array(40218);
		when "1001110100011011" => data_out <= rom_array(40219);
		when "1001110100011100" => data_out <= rom_array(40220);
		when "1001110100011101" => data_out <= rom_array(40221);
		when "1001110100011110" => data_out <= rom_array(40222);
		when "1001110100011111" => data_out <= rom_array(40223);
		when "1001110100100000" => data_out <= rom_array(40224);
		when "1001110100100001" => data_out <= rom_array(40225);
		when "1001110100100010" => data_out <= rom_array(40226);
		when "1001110100100011" => data_out <= rom_array(40227);
		when "1001110100100100" => data_out <= rom_array(40228);
		when "1001110100100101" => data_out <= rom_array(40229);
		when "1001110100100110" => data_out <= rom_array(40230);
		when "1001110100100111" => data_out <= rom_array(40231);
		when "1001110100101000" => data_out <= rom_array(40232);
		when "1001110100101001" => data_out <= rom_array(40233);
		when "1001110100101010" => data_out <= rom_array(40234);
		when "1001110100101011" => data_out <= rom_array(40235);
		when "1001110100101100" => data_out <= rom_array(40236);
		when "1001110100101101" => data_out <= rom_array(40237);
		when "1001110100101110" => data_out <= rom_array(40238);
		when "1001110100101111" => data_out <= rom_array(40239);
		when "1001110100110000" => data_out <= rom_array(40240);
		when "1001110100110001" => data_out <= rom_array(40241);
		when "1001110100110010" => data_out <= rom_array(40242);
		when "1001110100110011" => data_out <= rom_array(40243);
		when "1001110100110100" => data_out <= rom_array(40244);
		when "1001110100110101" => data_out <= rom_array(40245);
		when "1001110100110110" => data_out <= rom_array(40246);
		when "1001110100110111" => data_out <= rom_array(40247);
		when "1001110100111000" => data_out <= rom_array(40248);
		when "1001110100111001" => data_out <= rom_array(40249);
		when "1001110100111010" => data_out <= rom_array(40250);
		when "1001110100111011" => data_out <= rom_array(40251);
		when "1001110100111100" => data_out <= rom_array(40252);
		when "1001110100111101" => data_out <= rom_array(40253);
		when "1001110100111110" => data_out <= rom_array(40254);
		when "1001110100111111" => data_out <= rom_array(40255);
		when "1001110101000000" => data_out <= rom_array(40256);
		when "1001110101000001" => data_out <= rom_array(40257);
		when "1001110101000010" => data_out <= rom_array(40258);
		when "1001110101000011" => data_out <= rom_array(40259);
		when "1001110101000100" => data_out <= rom_array(40260);
		when "1001110101000101" => data_out <= rom_array(40261);
		when "1001110101000110" => data_out <= rom_array(40262);
		when "1001110101000111" => data_out <= rom_array(40263);
		when "1001110101001000" => data_out <= rom_array(40264);
		when "1001110101001001" => data_out <= rom_array(40265);
		when "1001110101001010" => data_out <= rom_array(40266);
		when "1001110101001011" => data_out <= rom_array(40267);
		when "1001110101001100" => data_out <= rom_array(40268);
		when "1001110101001101" => data_out <= rom_array(40269);
		when "1001110101001110" => data_out <= rom_array(40270);
		when "1001110101001111" => data_out <= rom_array(40271);
		when "1001110101010000" => data_out <= rom_array(40272);
		when "1001110101010001" => data_out <= rom_array(40273);
		when "1001110101010010" => data_out <= rom_array(40274);
		when "1001110101010011" => data_out <= rom_array(40275);
		when "1001110101010100" => data_out <= rom_array(40276);
		when "1001110101010101" => data_out <= rom_array(40277);
		when "1001110101010110" => data_out <= rom_array(40278);
		when "1001110101010111" => data_out <= rom_array(40279);
		when "1001110101011000" => data_out <= rom_array(40280);
		when "1001110101011001" => data_out <= rom_array(40281);
		when "1001110101011010" => data_out <= rom_array(40282);
		when "1001110101011011" => data_out <= rom_array(40283);
		when "1001110101011100" => data_out <= rom_array(40284);
		when "1001110101011101" => data_out <= rom_array(40285);
		when "1001110101011110" => data_out <= rom_array(40286);
		when "1001110101011111" => data_out <= rom_array(40287);
		when "1001110101100000" => data_out <= rom_array(40288);
		when "1001110101100001" => data_out <= rom_array(40289);
		when "1001110101100010" => data_out <= rom_array(40290);
		when "1001110101100011" => data_out <= rom_array(40291);
		when "1001110101100100" => data_out <= rom_array(40292);
		when "1001110101100101" => data_out <= rom_array(40293);
		when "1001110101100110" => data_out <= rom_array(40294);
		when "1001110101100111" => data_out <= rom_array(40295);
		when "1001110101101000" => data_out <= rom_array(40296);
		when "1001110101101001" => data_out <= rom_array(40297);
		when "1001110101101010" => data_out <= rom_array(40298);
		when "1001110101101011" => data_out <= rom_array(40299);
		when "1001110101101100" => data_out <= rom_array(40300);
		when "1001110101101101" => data_out <= rom_array(40301);
		when "1001110101101110" => data_out <= rom_array(40302);
		when "1001110101101111" => data_out <= rom_array(40303);
		when "1001110101110000" => data_out <= rom_array(40304);
		when "1001110101110001" => data_out <= rom_array(40305);
		when "1001110101110010" => data_out <= rom_array(40306);
		when "1001110101110011" => data_out <= rom_array(40307);
		when "1001110101110100" => data_out <= rom_array(40308);
		when "1001110101110101" => data_out <= rom_array(40309);
		when "1001110101110110" => data_out <= rom_array(40310);
		when "1001110101110111" => data_out <= rom_array(40311);
		when "1001110101111000" => data_out <= rom_array(40312);
		when "1001110101111001" => data_out <= rom_array(40313);
		when "1001110101111010" => data_out <= rom_array(40314);
		when "1001110101111011" => data_out <= rom_array(40315);
		when "1001110101111100" => data_out <= rom_array(40316);
		when "1001110101111101" => data_out <= rom_array(40317);
		when "1001110101111110" => data_out <= rom_array(40318);
		when "1001110101111111" => data_out <= rom_array(40319);
		when "1001110110000000" => data_out <= rom_array(40320);
		when "1001110110000001" => data_out <= rom_array(40321);
		when "1001110110000010" => data_out <= rom_array(40322);
		when "1001110110000011" => data_out <= rom_array(40323);
		when "1001110110000100" => data_out <= rom_array(40324);
		when "1001110110000101" => data_out <= rom_array(40325);
		when "1001110110000110" => data_out <= rom_array(40326);
		when "1001110110000111" => data_out <= rom_array(40327);
		when "1001110110001000" => data_out <= rom_array(40328);
		when "1001110110001001" => data_out <= rom_array(40329);
		when "1001110110001010" => data_out <= rom_array(40330);
		when "1001110110001011" => data_out <= rom_array(40331);
		when "1001110110001100" => data_out <= rom_array(40332);
		when "1001110110001101" => data_out <= rom_array(40333);
		when "1001110110001110" => data_out <= rom_array(40334);
		when "1001110110001111" => data_out <= rom_array(40335);
		when "1001110110010000" => data_out <= rom_array(40336);
		when "1001110110010001" => data_out <= rom_array(40337);
		when "1001110110010010" => data_out <= rom_array(40338);
		when "1001110110010011" => data_out <= rom_array(40339);
		when "1001110110010100" => data_out <= rom_array(40340);
		when "1001110110010101" => data_out <= rom_array(40341);
		when "1001110110010110" => data_out <= rom_array(40342);
		when "1001110110010111" => data_out <= rom_array(40343);
		when "1001110110011000" => data_out <= rom_array(40344);
		when "1001110110011001" => data_out <= rom_array(40345);
		when "1001110110011010" => data_out <= rom_array(40346);
		when "1001110110011011" => data_out <= rom_array(40347);
		when "1001110110011100" => data_out <= rom_array(40348);
		when "1001110110011101" => data_out <= rom_array(40349);
		when "1001110110011110" => data_out <= rom_array(40350);
		when "1001110110011111" => data_out <= rom_array(40351);
		when "1001110110100000" => data_out <= rom_array(40352);
		when "1001110110100001" => data_out <= rom_array(40353);
		when "1001110110100010" => data_out <= rom_array(40354);
		when "1001110110100011" => data_out <= rom_array(40355);
		when "1001110110100100" => data_out <= rom_array(40356);
		when "1001110110100101" => data_out <= rom_array(40357);
		when "1001110110100110" => data_out <= rom_array(40358);
		when "1001110110100111" => data_out <= rom_array(40359);
		when "1001110110101000" => data_out <= rom_array(40360);
		when "1001110110101001" => data_out <= rom_array(40361);
		when "1001110110101010" => data_out <= rom_array(40362);
		when "1001110110101011" => data_out <= rom_array(40363);
		when "1001110110101100" => data_out <= rom_array(40364);
		when "1001110110101101" => data_out <= rom_array(40365);
		when "1001110110101110" => data_out <= rom_array(40366);
		when "1001110110101111" => data_out <= rom_array(40367);
		when "1001110110110000" => data_out <= rom_array(40368);
		when "1001110110110001" => data_out <= rom_array(40369);
		when "1001110110110010" => data_out <= rom_array(40370);
		when "1001110110110011" => data_out <= rom_array(40371);
		when "1001110110110100" => data_out <= rom_array(40372);
		when "1001110110110101" => data_out <= rom_array(40373);
		when "1001110110110110" => data_out <= rom_array(40374);
		when "1001110110110111" => data_out <= rom_array(40375);
		when "1001110110111000" => data_out <= rom_array(40376);
		when "1001110110111001" => data_out <= rom_array(40377);
		when "1001110110111010" => data_out <= rom_array(40378);
		when "1001110110111011" => data_out <= rom_array(40379);
		when "1001110110111100" => data_out <= rom_array(40380);
		when "1001110110111101" => data_out <= rom_array(40381);
		when "1001110110111110" => data_out <= rom_array(40382);
		when "1001110110111111" => data_out <= rom_array(40383);
		when "1001110111000000" => data_out <= rom_array(40384);
		when "1001110111000001" => data_out <= rom_array(40385);
		when "1001110111000010" => data_out <= rom_array(40386);
		when "1001110111000011" => data_out <= rom_array(40387);
		when "1001110111000100" => data_out <= rom_array(40388);
		when "1001110111000101" => data_out <= rom_array(40389);
		when "1001110111000110" => data_out <= rom_array(40390);
		when "1001110111000111" => data_out <= rom_array(40391);
		when "1001110111001000" => data_out <= rom_array(40392);
		when "1001110111001001" => data_out <= rom_array(40393);
		when "1001110111001010" => data_out <= rom_array(40394);
		when "1001110111001011" => data_out <= rom_array(40395);
		when "1001110111001100" => data_out <= rom_array(40396);
		when "1001110111001101" => data_out <= rom_array(40397);
		when "1001110111001110" => data_out <= rom_array(40398);
		when "1001110111001111" => data_out <= rom_array(40399);
		when "1001110111010000" => data_out <= rom_array(40400);
		when "1001110111010001" => data_out <= rom_array(40401);
		when "1001110111010010" => data_out <= rom_array(40402);
		when "1001110111010011" => data_out <= rom_array(40403);
		when "1001110111010100" => data_out <= rom_array(40404);
		when "1001110111010101" => data_out <= rom_array(40405);
		when "1001110111010110" => data_out <= rom_array(40406);
		when "1001110111010111" => data_out <= rom_array(40407);
		when "1001110111011000" => data_out <= rom_array(40408);
		when "1001110111011001" => data_out <= rom_array(40409);
		when "1001110111011010" => data_out <= rom_array(40410);
		when "1001110111011011" => data_out <= rom_array(40411);
		when "1001110111011100" => data_out <= rom_array(40412);
		when "1001110111011101" => data_out <= rom_array(40413);
		when "1001110111011110" => data_out <= rom_array(40414);
		when "1001110111011111" => data_out <= rom_array(40415);
		when "1001110111100000" => data_out <= rom_array(40416);
		when "1001110111100001" => data_out <= rom_array(40417);
		when "1001110111100010" => data_out <= rom_array(40418);
		when "1001110111100011" => data_out <= rom_array(40419);
		when "1001110111100100" => data_out <= rom_array(40420);
		when "1001110111100101" => data_out <= rom_array(40421);
		when "1001110111100110" => data_out <= rom_array(40422);
		when "1001110111100111" => data_out <= rom_array(40423);
		when "1001110111101000" => data_out <= rom_array(40424);
		when "1001110111101001" => data_out <= rom_array(40425);
		when "1001110111101010" => data_out <= rom_array(40426);
		when "1001110111101011" => data_out <= rom_array(40427);
		when "1001110111101100" => data_out <= rom_array(40428);
		when "1001110111101101" => data_out <= rom_array(40429);
		when "1001110111101110" => data_out <= rom_array(40430);
		when "1001110111101111" => data_out <= rom_array(40431);
		when "1001110111110000" => data_out <= rom_array(40432);
		when "1001110111110001" => data_out <= rom_array(40433);
		when "1001110111110010" => data_out <= rom_array(40434);
		when "1001110111110011" => data_out <= rom_array(40435);
		when "1001110111110100" => data_out <= rom_array(40436);
		when "1001110111110101" => data_out <= rom_array(40437);
		when "1001110111110110" => data_out <= rom_array(40438);
		when "1001110111110111" => data_out <= rom_array(40439);
		when "1001110111111000" => data_out <= rom_array(40440);
		when "1001110111111001" => data_out <= rom_array(40441);
		when "1001110111111010" => data_out <= rom_array(40442);
		when "1001110111111011" => data_out <= rom_array(40443);
		when "1001110111111100" => data_out <= rom_array(40444);
		when "1001110111111101" => data_out <= rom_array(40445);
		when "1001110111111110" => data_out <= rom_array(40446);
		when "1001110111111111" => data_out <= rom_array(40447);
		when "1001111000000000" => data_out <= rom_array(40448);
		when "1001111000000001" => data_out <= rom_array(40449);
		when "1001111000000010" => data_out <= rom_array(40450);
		when "1001111000000011" => data_out <= rom_array(40451);
		when "1001111000000100" => data_out <= rom_array(40452);
		when "1001111000000101" => data_out <= rom_array(40453);
		when "1001111000000110" => data_out <= rom_array(40454);
		when "1001111000000111" => data_out <= rom_array(40455);
		when "1001111000001000" => data_out <= rom_array(40456);
		when "1001111000001001" => data_out <= rom_array(40457);
		when "1001111000001010" => data_out <= rom_array(40458);
		when "1001111000001011" => data_out <= rom_array(40459);
		when "1001111000001100" => data_out <= rom_array(40460);
		when "1001111000001101" => data_out <= rom_array(40461);
		when "1001111000001110" => data_out <= rom_array(40462);
		when "1001111000001111" => data_out <= rom_array(40463);
		when "1001111000010000" => data_out <= rom_array(40464);
		when "1001111000010001" => data_out <= rom_array(40465);
		when "1001111000010010" => data_out <= rom_array(40466);
		when "1001111000010011" => data_out <= rom_array(40467);
		when "1001111000010100" => data_out <= rom_array(40468);
		when "1001111000010101" => data_out <= rom_array(40469);
		when "1001111000010110" => data_out <= rom_array(40470);
		when "1001111000010111" => data_out <= rom_array(40471);
		when "1001111000011000" => data_out <= rom_array(40472);
		when "1001111000011001" => data_out <= rom_array(40473);
		when "1001111000011010" => data_out <= rom_array(40474);
		when "1001111000011011" => data_out <= rom_array(40475);
		when "1001111000011100" => data_out <= rom_array(40476);
		when "1001111000011101" => data_out <= rom_array(40477);
		when "1001111000011110" => data_out <= rom_array(40478);
		when "1001111000011111" => data_out <= rom_array(40479);
		when "1001111000100000" => data_out <= rom_array(40480);
		when "1001111000100001" => data_out <= rom_array(40481);
		when "1001111000100010" => data_out <= rom_array(40482);
		when "1001111000100011" => data_out <= rom_array(40483);
		when "1001111000100100" => data_out <= rom_array(40484);
		when "1001111000100101" => data_out <= rom_array(40485);
		when "1001111000100110" => data_out <= rom_array(40486);
		when "1001111000100111" => data_out <= rom_array(40487);
		when "1001111000101000" => data_out <= rom_array(40488);
		when "1001111000101001" => data_out <= rom_array(40489);
		when "1001111000101010" => data_out <= rom_array(40490);
		when "1001111000101011" => data_out <= rom_array(40491);
		when "1001111000101100" => data_out <= rom_array(40492);
		when "1001111000101101" => data_out <= rom_array(40493);
		when "1001111000101110" => data_out <= rom_array(40494);
		when "1001111000101111" => data_out <= rom_array(40495);
		when "1001111000110000" => data_out <= rom_array(40496);
		when "1001111000110001" => data_out <= rom_array(40497);
		when "1001111000110010" => data_out <= rom_array(40498);
		when "1001111000110011" => data_out <= rom_array(40499);
		when "1001111000110100" => data_out <= rom_array(40500);
		when "1001111000110101" => data_out <= rom_array(40501);
		when "1001111000110110" => data_out <= rom_array(40502);
		when "1001111000110111" => data_out <= rom_array(40503);
		when "1001111000111000" => data_out <= rom_array(40504);
		when "1001111000111001" => data_out <= rom_array(40505);
		when "1001111000111010" => data_out <= rom_array(40506);
		when "1001111000111011" => data_out <= rom_array(40507);
		when "1001111000111100" => data_out <= rom_array(40508);
		when "1001111000111101" => data_out <= rom_array(40509);
		when "1001111000111110" => data_out <= rom_array(40510);
		when "1001111000111111" => data_out <= rom_array(40511);
		when "1001111001000000" => data_out <= rom_array(40512);
		when "1001111001000001" => data_out <= rom_array(40513);
		when "1001111001000010" => data_out <= rom_array(40514);
		when "1001111001000011" => data_out <= rom_array(40515);
		when "1001111001000100" => data_out <= rom_array(40516);
		when "1001111001000101" => data_out <= rom_array(40517);
		when "1001111001000110" => data_out <= rom_array(40518);
		when "1001111001000111" => data_out <= rom_array(40519);
		when "1001111001001000" => data_out <= rom_array(40520);
		when "1001111001001001" => data_out <= rom_array(40521);
		when "1001111001001010" => data_out <= rom_array(40522);
		when "1001111001001011" => data_out <= rom_array(40523);
		when "1001111001001100" => data_out <= rom_array(40524);
		when "1001111001001101" => data_out <= rom_array(40525);
		when "1001111001001110" => data_out <= rom_array(40526);
		when "1001111001001111" => data_out <= rom_array(40527);
		when "1001111001010000" => data_out <= rom_array(40528);
		when "1001111001010001" => data_out <= rom_array(40529);
		when "1001111001010010" => data_out <= rom_array(40530);
		when "1001111001010011" => data_out <= rom_array(40531);
		when "1001111001010100" => data_out <= rom_array(40532);
		when "1001111001010101" => data_out <= rom_array(40533);
		when "1001111001010110" => data_out <= rom_array(40534);
		when "1001111001010111" => data_out <= rom_array(40535);
		when "1001111001011000" => data_out <= rom_array(40536);
		when "1001111001011001" => data_out <= rom_array(40537);
		when "1001111001011010" => data_out <= rom_array(40538);
		when "1001111001011011" => data_out <= rom_array(40539);
		when "1001111001011100" => data_out <= rom_array(40540);
		when "1001111001011101" => data_out <= rom_array(40541);
		when "1001111001011110" => data_out <= rom_array(40542);
		when "1001111001011111" => data_out <= rom_array(40543);
		when "1001111001100000" => data_out <= rom_array(40544);
		when "1001111001100001" => data_out <= rom_array(40545);
		when "1001111001100010" => data_out <= rom_array(40546);
		when "1001111001100011" => data_out <= rom_array(40547);
		when "1001111001100100" => data_out <= rom_array(40548);
		when "1001111001100101" => data_out <= rom_array(40549);
		when "1001111001100110" => data_out <= rom_array(40550);
		when "1001111001100111" => data_out <= rom_array(40551);
		when "1001111001101000" => data_out <= rom_array(40552);
		when "1001111001101001" => data_out <= rom_array(40553);
		when "1001111001101010" => data_out <= rom_array(40554);
		when "1001111001101011" => data_out <= rom_array(40555);
		when "1001111001101100" => data_out <= rom_array(40556);
		when "1001111001101101" => data_out <= rom_array(40557);
		when "1001111001101110" => data_out <= rom_array(40558);
		when "1001111001101111" => data_out <= rom_array(40559);
		when "1001111001110000" => data_out <= rom_array(40560);
		when "1001111001110001" => data_out <= rom_array(40561);
		when "1001111001110010" => data_out <= rom_array(40562);
		when "1001111001110011" => data_out <= rom_array(40563);
		when "1001111001110100" => data_out <= rom_array(40564);
		when "1001111001110101" => data_out <= rom_array(40565);
		when "1001111001110110" => data_out <= rom_array(40566);
		when "1001111001110111" => data_out <= rom_array(40567);
		when "1001111001111000" => data_out <= rom_array(40568);
		when "1001111001111001" => data_out <= rom_array(40569);
		when "1001111001111010" => data_out <= rom_array(40570);
		when "1001111001111011" => data_out <= rom_array(40571);
		when "1001111001111100" => data_out <= rom_array(40572);
		when "1001111001111101" => data_out <= rom_array(40573);
		when "1001111001111110" => data_out <= rom_array(40574);
		when "1001111001111111" => data_out <= rom_array(40575);
		when "1001111010000000" => data_out <= rom_array(40576);
		when "1001111010000001" => data_out <= rom_array(40577);
		when "1001111010000010" => data_out <= rom_array(40578);
		when "1001111010000011" => data_out <= rom_array(40579);
		when "1001111010000100" => data_out <= rom_array(40580);
		when "1001111010000101" => data_out <= rom_array(40581);
		when "1001111010000110" => data_out <= rom_array(40582);
		when "1001111010000111" => data_out <= rom_array(40583);
		when "1001111010001000" => data_out <= rom_array(40584);
		when "1001111010001001" => data_out <= rom_array(40585);
		when "1001111010001010" => data_out <= rom_array(40586);
		when "1001111010001011" => data_out <= rom_array(40587);
		when "1001111010001100" => data_out <= rom_array(40588);
		when "1001111010001101" => data_out <= rom_array(40589);
		when "1001111010001110" => data_out <= rom_array(40590);
		when "1001111010001111" => data_out <= rom_array(40591);
		when "1001111010010000" => data_out <= rom_array(40592);
		when "1001111010010001" => data_out <= rom_array(40593);
		when "1001111010010010" => data_out <= rom_array(40594);
		when "1001111010010011" => data_out <= rom_array(40595);
		when "1001111010010100" => data_out <= rom_array(40596);
		when "1001111010010101" => data_out <= rom_array(40597);
		when "1001111010010110" => data_out <= rom_array(40598);
		when "1001111010010111" => data_out <= rom_array(40599);
		when "1001111010011000" => data_out <= rom_array(40600);
		when "1001111010011001" => data_out <= rom_array(40601);
		when "1001111010011010" => data_out <= rom_array(40602);
		when "1001111010011011" => data_out <= rom_array(40603);
		when "1001111010011100" => data_out <= rom_array(40604);
		when "1001111010011101" => data_out <= rom_array(40605);
		when "1001111010011110" => data_out <= rom_array(40606);
		when "1001111010011111" => data_out <= rom_array(40607);
		when "1001111010100000" => data_out <= rom_array(40608);
		when "1001111010100001" => data_out <= rom_array(40609);
		when "1001111010100010" => data_out <= rom_array(40610);
		when "1001111010100011" => data_out <= rom_array(40611);
		when "1001111010100100" => data_out <= rom_array(40612);
		when "1001111010100101" => data_out <= rom_array(40613);
		when "1001111010100110" => data_out <= rom_array(40614);
		when "1001111010100111" => data_out <= rom_array(40615);
		when "1001111010101000" => data_out <= rom_array(40616);
		when "1001111010101001" => data_out <= rom_array(40617);
		when "1001111010101010" => data_out <= rom_array(40618);
		when "1001111010101011" => data_out <= rom_array(40619);
		when "1001111010101100" => data_out <= rom_array(40620);
		when "1001111010101101" => data_out <= rom_array(40621);
		when "1001111010101110" => data_out <= rom_array(40622);
		when "1001111010101111" => data_out <= rom_array(40623);
		when "1001111010110000" => data_out <= rom_array(40624);
		when "1001111010110001" => data_out <= rom_array(40625);
		when "1001111010110010" => data_out <= rom_array(40626);
		when "1001111010110011" => data_out <= rom_array(40627);
		when "1001111010110100" => data_out <= rom_array(40628);
		when "1001111010110101" => data_out <= rom_array(40629);
		when "1001111010110110" => data_out <= rom_array(40630);
		when "1001111010110111" => data_out <= rom_array(40631);
		when "1001111010111000" => data_out <= rom_array(40632);
		when "1001111010111001" => data_out <= rom_array(40633);
		when "1001111010111010" => data_out <= rom_array(40634);
		when "1001111010111011" => data_out <= rom_array(40635);
		when "1001111010111100" => data_out <= rom_array(40636);
		when "1001111010111101" => data_out <= rom_array(40637);
		when "1001111010111110" => data_out <= rom_array(40638);
		when "1001111010111111" => data_out <= rom_array(40639);
		when "1001111011000000" => data_out <= rom_array(40640);
		when "1001111011000001" => data_out <= rom_array(40641);
		when "1001111011000010" => data_out <= rom_array(40642);
		when "1001111011000011" => data_out <= rom_array(40643);
		when "1001111011000100" => data_out <= rom_array(40644);
		when "1001111011000101" => data_out <= rom_array(40645);
		when "1001111011000110" => data_out <= rom_array(40646);
		when "1001111011000111" => data_out <= rom_array(40647);
		when "1001111011001000" => data_out <= rom_array(40648);
		when "1001111011001001" => data_out <= rom_array(40649);
		when "1001111011001010" => data_out <= rom_array(40650);
		when "1001111011001011" => data_out <= rom_array(40651);
		when "1001111011001100" => data_out <= rom_array(40652);
		when "1001111011001101" => data_out <= rom_array(40653);
		when "1001111011001110" => data_out <= rom_array(40654);
		when "1001111011001111" => data_out <= rom_array(40655);
		when "1001111011010000" => data_out <= rom_array(40656);
		when "1001111011010001" => data_out <= rom_array(40657);
		when "1001111011010010" => data_out <= rom_array(40658);
		when "1001111011010011" => data_out <= rom_array(40659);
		when "1001111011010100" => data_out <= rom_array(40660);
		when "1001111011010101" => data_out <= rom_array(40661);
		when "1001111011010110" => data_out <= rom_array(40662);
		when "1001111011010111" => data_out <= rom_array(40663);
		when "1001111011011000" => data_out <= rom_array(40664);
		when "1001111011011001" => data_out <= rom_array(40665);
		when "1001111011011010" => data_out <= rom_array(40666);
		when "1001111011011011" => data_out <= rom_array(40667);
		when "1001111011011100" => data_out <= rom_array(40668);
		when "1001111011011101" => data_out <= rom_array(40669);
		when "1001111011011110" => data_out <= rom_array(40670);
		when "1001111011011111" => data_out <= rom_array(40671);
		when "1001111011100000" => data_out <= rom_array(40672);
		when "1001111011100001" => data_out <= rom_array(40673);
		when "1001111011100010" => data_out <= rom_array(40674);
		when "1001111011100011" => data_out <= rom_array(40675);
		when "1001111011100100" => data_out <= rom_array(40676);
		when "1001111011100101" => data_out <= rom_array(40677);
		when "1001111011100110" => data_out <= rom_array(40678);
		when "1001111011100111" => data_out <= rom_array(40679);
		when "1001111011101000" => data_out <= rom_array(40680);
		when "1001111011101001" => data_out <= rom_array(40681);
		when "1001111011101010" => data_out <= rom_array(40682);
		when "1001111011101011" => data_out <= rom_array(40683);
		when "1001111011101100" => data_out <= rom_array(40684);
		when "1001111011101101" => data_out <= rom_array(40685);
		when "1001111011101110" => data_out <= rom_array(40686);
		when "1001111011101111" => data_out <= rom_array(40687);
		when "1001111011110000" => data_out <= rom_array(40688);
		when "1001111011110001" => data_out <= rom_array(40689);
		when "1001111011110010" => data_out <= rom_array(40690);
		when "1001111011110011" => data_out <= rom_array(40691);
		when "1001111011110100" => data_out <= rom_array(40692);
		when "1001111011110101" => data_out <= rom_array(40693);
		when "1001111011110110" => data_out <= rom_array(40694);
		when "1001111011110111" => data_out <= rom_array(40695);
		when "1001111011111000" => data_out <= rom_array(40696);
		when "1001111011111001" => data_out <= rom_array(40697);
		when "1001111011111010" => data_out <= rom_array(40698);
		when "1001111011111011" => data_out <= rom_array(40699);
		when "1001111011111100" => data_out <= rom_array(40700);
		when "1001111011111101" => data_out <= rom_array(40701);
		when "1001111011111110" => data_out <= rom_array(40702);
		when "1001111011111111" => data_out <= rom_array(40703);
		when "1001111100000000" => data_out <= rom_array(40704);
		when "1001111100000001" => data_out <= rom_array(40705);
		when "1001111100000010" => data_out <= rom_array(40706);
		when "1001111100000011" => data_out <= rom_array(40707);
		when "1001111100000100" => data_out <= rom_array(40708);
		when "1001111100000101" => data_out <= rom_array(40709);
		when "1001111100000110" => data_out <= rom_array(40710);
		when "1001111100000111" => data_out <= rom_array(40711);
		when "1001111100001000" => data_out <= rom_array(40712);
		when "1001111100001001" => data_out <= rom_array(40713);
		when "1001111100001010" => data_out <= rom_array(40714);
		when "1001111100001011" => data_out <= rom_array(40715);
		when "1001111100001100" => data_out <= rom_array(40716);
		when "1001111100001101" => data_out <= rom_array(40717);
		when "1001111100001110" => data_out <= rom_array(40718);
		when "1001111100001111" => data_out <= rom_array(40719);
		when "1001111100010000" => data_out <= rom_array(40720);
		when "1001111100010001" => data_out <= rom_array(40721);
		when "1001111100010010" => data_out <= rom_array(40722);
		when "1001111100010011" => data_out <= rom_array(40723);
		when "1001111100010100" => data_out <= rom_array(40724);
		when "1001111100010101" => data_out <= rom_array(40725);
		when "1001111100010110" => data_out <= rom_array(40726);
		when "1001111100010111" => data_out <= rom_array(40727);
		when "1001111100011000" => data_out <= rom_array(40728);
		when "1001111100011001" => data_out <= rom_array(40729);
		when "1001111100011010" => data_out <= rom_array(40730);
		when "1001111100011011" => data_out <= rom_array(40731);
		when "1001111100011100" => data_out <= rom_array(40732);
		when "1001111100011101" => data_out <= rom_array(40733);
		when "1001111100011110" => data_out <= rom_array(40734);
		when "1001111100011111" => data_out <= rom_array(40735);
		when "1001111100100000" => data_out <= rom_array(40736);
		when "1001111100100001" => data_out <= rom_array(40737);
		when "1001111100100010" => data_out <= rom_array(40738);
		when "1001111100100011" => data_out <= rom_array(40739);
		when "1001111100100100" => data_out <= rom_array(40740);
		when "1001111100100101" => data_out <= rom_array(40741);
		when "1001111100100110" => data_out <= rom_array(40742);
		when "1001111100100111" => data_out <= rom_array(40743);
		when "1001111100101000" => data_out <= rom_array(40744);
		when "1001111100101001" => data_out <= rom_array(40745);
		when "1001111100101010" => data_out <= rom_array(40746);
		when "1001111100101011" => data_out <= rom_array(40747);
		when "1001111100101100" => data_out <= rom_array(40748);
		when "1001111100101101" => data_out <= rom_array(40749);
		when "1001111100101110" => data_out <= rom_array(40750);
		when "1001111100101111" => data_out <= rom_array(40751);
		when "1001111100110000" => data_out <= rom_array(40752);
		when "1001111100110001" => data_out <= rom_array(40753);
		when "1001111100110010" => data_out <= rom_array(40754);
		when "1001111100110011" => data_out <= rom_array(40755);
		when "1001111100110100" => data_out <= rom_array(40756);
		when "1001111100110101" => data_out <= rom_array(40757);
		when "1001111100110110" => data_out <= rom_array(40758);
		when "1001111100110111" => data_out <= rom_array(40759);
		when "1001111100111000" => data_out <= rom_array(40760);
		when "1001111100111001" => data_out <= rom_array(40761);
		when "1001111100111010" => data_out <= rom_array(40762);
		when "1001111100111011" => data_out <= rom_array(40763);
		when "1001111100111100" => data_out <= rom_array(40764);
		when "1001111100111101" => data_out <= rom_array(40765);
		when "1001111100111110" => data_out <= rom_array(40766);
		when "1001111100111111" => data_out <= rom_array(40767);
		when "1001111101000000" => data_out <= rom_array(40768);
		when "1001111101000001" => data_out <= rom_array(40769);
		when "1001111101000010" => data_out <= rom_array(40770);
		when "1001111101000011" => data_out <= rom_array(40771);
		when "1001111101000100" => data_out <= rom_array(40772);
		when "1001111101000101" => data_out <= rom_array(40773);
		when "1001111101000110" => data_out <= rom_array(40774);
		when "1001111101000111" => data_out <= rom_array(40775);
		when "1001111101001000" => data_out <= rom_array(40776);
		when "1001111101001001" => data_out <= rom_array(40777);
		when "1001111101001010" => data_out <= rom_array(40778);
		when "1001111101001011" => data_out <= rom_array(40779);
		when "1001111101001100" => data_out <= rom_array(40780);
		when "1001111101001101" => data_out <= rom_array(40781);
		when "1001111101001110" => data_out <= rom_array(40782);
		when "1001111101001111" => data_out <= rom_array(40783);
		when "1001111101010000" => data_out <= rom_array(40784);
		when "1001111101010001" => data_out <= rom_array(40785);
		when "1001111101010010" => data_out <= rom_array(40786);
		when "1001111101010011" => data_out <= rom_array(40787);
		when "1001111101010100" => data_out <= rom_array(40788);
		when "1001111101010101" => data_out <= rom_array(40789);
		when "1001111101010110" => data_out <= rom_array(40790);
		when "1001111101010111" => data_out <= rom_array(40791);
		when "1001111101011000" => data_out <= rom_array(40792);
		when "1001111101011001" => data_out <= rom_array(40793);
		when "1001111101011010" => data_out <= rom_array(40794);
		when "1001111101011011" => data_out <= rom_array(40795);
		when "1001111101011100" => data_out <= rom_array(40796);
		when "1001111101011101" => data_out <= rom_array(40797);
		when "1001111101011110" => data_out <= rom_array(40798);
		when "1001111101011111" => data_out <= rom_array(40799);
		when "1001111101100000" => data_out <= rom_array(40800);
		when "1001111101100001" => data_out <= rom_array(40801);
		when "1001111101100010" => data_out <= rom_array(40802);
		when "1001111101100011" => data_out <= rom_array(40803);
		when "1001111101100100" => data_out <= rom_array(40804);
		when "1001111101100101" => data_out <= rom_array(40805);
		when "1001111101100110" => data_out <= rom_array(40806);
		when "1001111101100111" => data_out <= rom_array(40807);
		when "1001111101101000" => data_out <= rom_array(40808);
		when "1001111101101001" => data_out <= rom_array(40809);
		when "1001111101101010" => data_out <= rom_array(40810);
		when "1001111101101011" => data_out <= rom_array(40811);
		when "1001111101101100" => data_out <= rom_array(40812);
		when "1001111101101101" => data_out <= rom_array(40813);
		when "1001111101101110" => data_out <= rom_array(40814);
		when "1001111101101111" => data_out <= rom_array(40815);
		when "1001111101110000" => data_out <= rom_array(40816);
		when "1001111101110001" => data_out <= rom_array(40817);
		when "1001111101110010" => data_out <= rom_array(40818);
		when "1001111101110011" => data_out <= rom_array(40819);
		when "1001111101110100" => data_out <= rom_array(40820);
		when "1001111101110101" => data_out <= rom_array(40821);
		when "1001111101110110" => data_out <= rom_array(40822);
		when "1001111101110111" => data_out <= rom_array(40823);
		when "1001111101111000" => data_out <= rom_array(40824);
		when "1001111101111001" => data_out <= rom_array(40825);
		when "1001111101111010" => data_out <= rom_array(40826);
		when "1001111101111011" => data_out <= rom_array(40827);
		when "1001111101111100" => data_out <= rom_array(40828);
		when "1001111101111101" => data_out <= rom_array(40829);
		when "1001111101111110" => data_out <= rom_array(40830);
		when "1001111101111111" => data_out <= rom_array(40831);
		when "1001111110000000" => data_out <= rom_array(40832);
		when "1001111110000001" => data_out <= rom_array(40833);
		when "1001111110000010" => data_out <= rom_array(40834);
		when "1001111110000011" => data_out <= rom_array(40835);
		when "1001111110000100" => data_out <= rom_array(40836);
		when "1001111110000101" => data_out <= rom_array(40837);
		when "1001111110000110" => data_out <= rom_array(40838);
		when "1001111110000111" => data_out <= rom_array(40839);
		when "1001111110001000" => data_out <= rom_array(40840);
		when "1001111110001001" => data_out <= rom_array(40841);
		when "1001111110001010" => data_out <= rom_array(40842);
		when "1001111110001011" => data_out <= rom_array(40843);
		when "1001111110001100" => data_out <= rom_array(40844);
		when "1001111110001101" => data_out <= rom_array(40845);
		when "1001111110001110" => data_out <= rom_array(40846);
		when "1001111110001111" => data_out <= rom_array(40847);
		when "1001111110010000" => data_out <= rom_array(40848);
		when "1001111110010001" => data_out <= rom_array(40849);
		when "1001111110010010" => data_out <= rom_array(40850);
		when "1001111110010011" => data_out <= rom_array(40851);
		when "1001111110010100" => data_out <= rom_array(40852);
		when "1001111110010101" => data_out <= rom_array(40853);
		when "1001111110010110" => data_out <= rom_array(40854);
		when "1001111110010111" => data_out <= rom_array(40855);
		when "1001111110011000" => data_out <= rom_array(40856);
		when "1001111110011001" => data_out <= rom_array(40857);
		when "1001111110011010" => data_out <= rom_array(40858);
		when "1001111110011011" => data_out <= rom_array(40859);
		when "1001111110011100" => data_out <= rom_array(40860);
		when "1001111110011101" => data_out <= rom_array(40861);
		when "1001111110011110" => data_out <= rom_array(40862);
		when "1001111110011111" => data_out <= rom_array(40863);
		when "1001111110100000" => data_out <= rom_array(40864);
		when "1001111110100001" => data_out <= rom_array(40865);
		when "1001111110100010" => data_out <= rom_array(40866);
		when "1001111110100011" => data_out <= rom_array(40867);
		when "1001111110100100" => data_out <= rom_array(40868);
		when "1001111110100101" => data_out <= rom_array(40869);
		when "1001111110100110" => data_out <= rom_array(40870);
		when "1001111110100111" => data_out <= rom_array(40871);
		when "1001111110101000" => data_out <= rom_array(40872);
		when "1001111110101001" => data_out <= rom_array(40873);
		when "1001111110101010" => data_out <= rom_array(40874);
		when "1001111110101011" => data_out <= rom_array(40875);
		when "1001111110101100" => data_out <= rom_array(40876);
		when "1001111110101101" => data_out <= rom_array(40877);
		when "1001111110101110" => data_out <= rom_array(40878);
		when "1001111110101111" => data_out <= rom_array(40879);
		when "1001111110110000" => data_out <= rom_array(40880);
		when "1001111110110001" => data_out <= rom_array(40881);
		when "1001111110110010" => data_out <= rom_array(40882);
		when "1001111110110011" => data_out <= rom_array(40883);
		when "1001111110110100" => data_out <= rom_array(40884);
		when "1001111110110101" => data_out <= rom_array(40885);
		when "1001111110110110" => data_out <= rom_array(40886);
		when "1001111110110111" => data_out <= rom_array(40887);
		when "1001111110111000" => data_out <= rom_array(40888);
		when "1001111110111001" => data_out <= rom_array(40889);
		when "1001111110111010" => data_out <= rom_array(40890);
		when "1001111110111011" => data_out <= rom_array(40891);
		when "1001111110111100" => data_out <= rom_array(40892);
		when "1001111110111101" => data_out <= rom_array(40893);
		when "1001111110111110" => data_out <= rom_array(40894);
		when "1001111110111111" => data_out <= rom_array(40895);
		when "1001111111000000" => data_out <= rom_array(40896);
		when "1001111111000001" => data_out <= rom_array(40897);
		when "1001111111000010" => data_out <= rom_array(40898);
		when "1001111111000011" => data_out <= rom_array(40899);
		when "1001111111000100" => data_out <= rom_array(40900);
		when "1001111111000101" => data_out <= rom_array(40901);
		when "1001111111000110" => data_out <= rom_array(40902);
		when "1001111111000111" => data_out <= rom_array(40903);
		when "1001111111001000" => data_out <= rom_array(40904);
		when "1001111111001001" => data_out <= rom_array(40905);
		when "1001111111001010" => data_out <= rom_array(40906);
		when "1001111111001011" => data_out <= rom_array(40907);
		when "1001111111001100" => data_out <= rom_array(40908);
		when "1001111111001101" => data_out <= rom_array(40909);
		when "1001111111001110" => data_out <= rom_array(40910);
		when "1001111111001111" => data_out <= rom_array(40911);
		when "1001111111010000" => data_out <= rom_array(40912);
		when "1001111111010001" => data_out <= rom_array(40913);
		when "1001111111010010" => data_out <= rom_array(40914);
		when "1001111111010011" => data_out <= rom_array(40915);
		when "1001111111010100" => data_out <= rom_array(40916);
		when "1001111111010101" => data_out <= rom_array(40917);
		when "1001111111010110" => data_out <= rom_array(40918);
		when "1001111111010111" => data_out <= rom_array(40919);
		when "1001111111011000" => data_out <= rom_array(40920);
		when "1001111111011001" => data_out <= rom_array(40921);
		when "1001111111011010" => data_out <= rom_array(40922);
		when "1001111111011011" => data_out <= rom_array(40923);
		when "1001111111011100" => data_out <= rom_array(40924);
		when "1001111111011101" => data_out <= rom_array(40925);
		when "1001111111011110" => data_out <= rom_array(40926);
		when "1001111111011111" => data_out <= rom_array(40927);
		when "1001111111100000" => data_out <= rom_array(40928);
		when "1001111111100001" => data_out <= rom_array(40929);
		when "1001111111100010" => data_out <= rom_array(40930);
		when "1001111111100011" => data_out <= rom_array(40931);
		when "1001111111100100" => data_out <= rom_array(40932);
		when "1001111111100101" => data_out <= rom_array(40933);
		when "1001111111100110" => data_out <= rom_array(40934);
		when "1001111111100111" => data_out <= rom_array(40935);
		when "1001111111101000" => data_out <= rom_array(40936);
		when "1001111111101001" => data_out <= rom_array(40937);
		when "1001111111101010" => data_out <= rom_array(40938);
		when "1001111111101011" => data_out <= rom_array(40939);
		when "1001111111101100" => data_out <= rom_array(40940);
		when "1001111111101101" => data_out <= rom_array(40941);
		when "1001111111101110" => data_out <= rom_array(40942);
		when "1001111111101111" => data_out <= rom_array(40943);
		when "1001111111110000" => data_out <= rom_array(40944);
		when "1001111111110001" => data_out <= rom_array(40945);
		when "1001111111110010" => data_out <= rom_array(40946);
		when "1001111111110011" => data_out <= rom_array(40947);
		when "1001111111110100" => data_out <= rom_array(40948);
		when "1001111111110101" => data_out <= rom_array(40949);
		when "1001111111110110" => data_out <= rom_array(40950);
		when "1001111111110111" => data_out <= rom_array(40951);
		when "1001111111111000" => data_out <= rom_array(40952);
		when "1001111111111001" => data_out <= rom_array(40953);
		when "1001111111111010" => data_out <= rom_array(40954);
		when "1001111111111011" => data_out <= rom_array(40955);
		when "1001111111111100" => data_out <= rom_array(40956);
		when "1001111111111101" => data_out <= rom_array(40957);
		when "1001111111111110" => data_out <= rom_array(40958);
		when "1001111111111111" => data_out <= rom_array(40959);
		when "1010000000000000" => data_out <= rom_array(40960);
		when "1010000000000001" => data_out <= rom_array(40961);
		when "1010000000000010" => data_out <= rom_array(40962);
		when "1010000000000011" => data_out <= rom_array(40963);
		when "1010000000000100" => data_out <= rom_array(40964);
		when "1010000000000101" => data_out <= rom_array(40965);
		when "1010000000000110" => data_out <= rom_array(40966);
		when "1010000000000111" => data_out <= rom_array(40967);
		when "1010000000001000" => data_out <= rom_array(40968);
		when "1010000000001001" => data_out <= rom_array(40969);
		when "1010000000001010" => data_out <= rom_array(40970);
		when "1010000000001011" => data_out <= rom_array(40971);
		when "1010000000001100" => data_out <= rom_array(40972);
		when "1010000000001101" => data_out <= rom_array(40973);
		when "1010000000001110" => data_out <= rom_array(40974);
		when "1010000000001111" => data_out <= rom_array(40975);
		when "1010000000010000" => data_out <= rom_array(40976);
		when "1010000000010001" => data_out <= rom_array(40977);
		when "1010000000010010" => data_out <= rom_array(40978);
		when "1010000000010011" => data_out <= rom_array(40979);
		when "1010000000010100" => data_out <= rom_array(40980);
		when "1010000000010101" => data_out <= rom_array(40981);
		when "1010000000010110" => data_out <= rom_array(40982);
		when "1010000000010111" => data_out <= rom_array(40983);
		when "1010000000011000" => data_out <= rom_array(40984);
		when "1010000000011001" => data_out <= rom_array(40985);
		when "1010000000011010" => data_out <= rom_array(40986);
		when "1010000000011011" => data_out <= rom_array(40987);
		when "1010000000011100" => data_out <= rom_array(40988);
		when "1010000000011101" => data_out <= rom_array(40989);
		when "1010000000011110" => data_out <= rom_array(40990);
		when "1010000000011111" => data_out <= rom_array(40991);
		when "1010000000100000" => data_out <= rom_array(40992);
		when "1010000000100001" => data_out <= rom_array(40993);
		when "1010000000100010" => data_out <= rom_array(40994);
		when "1010000000100011" => data_out <= rom_array(40995);
		when "1010000000100100" => data_out <= rom_array(40996);
		when "1010000000100101" => data_out <= rom_array(40997);
		when "1010000000100110" => data_out <= rom_array(40998);
		when "1010000000100111" => data_out <= rom_array(40999);
		when "1010000000101000" => data_out <= rom_array(41000);
		when "1010000000101001" => data_out <= rom_array(41001);
		when "1010000000101010" => data_out <= rom_array(41002);
		when "1010000000101011" => data_out <= rom_array(41003);
		when "1010000000101100" => data_out <= rom_array(41004);
		when "1010000000101101" => data_out <= rom_array(41005);
		when "1010000000101110" => data_out <= rom_array(41006);
		when "1010000000101111" => data_out <= rom_array(41007);
		when "1010000000110000" => data_out <= rom_array(41008);
		when "1010000000110001" => data_out <= rom_array(41009);
		when "1010000000110010" => data_out <= rom_array(41010);
		when "1010000000110011" => data_out <= rom_array(41011);
		when "1010000000110100" => data_out <= rom_array(41012);
		when "1010000000110101" => data_out <= rom_array(41013);
		when "1010000000110110" => data_out <= rom_array(41014);
		when "1010000000110111" => data_out <= rom_array(41015);
		when "1010000000111000" => data_out <= rom_array(41016);
		when "1010000000111001" => data_out <= rom_array(41017);
		when "1010000000111010" => data_out <= rom_array(41018);
		when "1010000000111011" => data_out <= rom_array(41019);
		when "1010000000111100" => data_out <= rom_array(41020);
		when "1010000000111101" => data_out <= rom_array(41021);
		when "1010000000111110" => data_out <= rom_array(41022);
		when "1010000000111111" => data_out <= rom_array(41023);
		when "1010000001000000" => data_out <= rom_array(41024);
		when "1010000001000001" => data_out <= rom_array(41025);
		when "1010000001000010" => data_out <= rom_array(41026);
		when "1010000001000011" => data_out <= rom_array(41027);
		when "1010000001000100" => data_out <= rom_array(41028);
		when "1010000001000101" => data_out <= rom_array(41029);
		when "1010000001000110" => data_out <= rom_array(41030);
		when "1010000001000111" => data_out <= rom_array(41031);
		when "1010000001001000" => data_out <= rom_array(41032);
		when "1010000001001001" => data_out <= rom_array(41033);
		when "1010000001001010" => data_out <= rom_array(41034);
		when "1010000001001011" => data_out <= rom_array(41035);
		when "1010000001001100" => data_out <= rom_array(41036);
		when "1010000001001101" => data_out <= rom_array(41037);
		when "1010000001001110" => data_out <= rom_array(41038);
		when "1010000001001111" => data_out <= rom_array(41039);
		when "1010000001010000" => data_out <= rom_array(41040);
		when "1010000001010001" => data_out <= rom_array(41041);
		when "1010000001010010" => data_out <= rom_array(41042);
		when "1010000001010011" => data_out <= rom_array(41043);
		when "1010000001010100" => data_out <= rom_array(41044);
		when "1010000001010101" => data_out <= rom_array(41045);
		when "1010000001010110" => data_out <= rom_array(41046);
		when "1010000001010111" => data_out <= rom_array(41047);
		when "1010000001011000" => data_out <= rom_array(41048);
		when "1010000001011001" => data_out <= rom_array(41049);
		when "1010000001011010" => data_out <= rom_array(41050);
		when "1010000001011011" => data_out <= rom_array(41051);
		when "1010000001011100" => data_out <= rom_array(41052);
		when "1010000001011101" => data_out <= rom_array(41053);
		when "1010000001011110" => data_out <= rom_array(41054);
		when "1010000001011111" => data_out <= rom_array(41055);
		when "1010000001100000" => data_out <= rom_array(41056);
		when "1010000001100001" => data_out <= rom_array(41057);
		when "1010000001100010" => data_out <= rom_array(41058);
		when "1010000001100011" => data_out <= rom_array(41059);
		when "1010000001100100" => data_out <= rom_array(41060);
		when "1010000001100101" => data_out <= rom_array(41061);
		when "1010000001100110" => data_out <= rom_array(41062);
		when "1010000001100111" => data_out <= rom_array(41063);
		when "1010000001101000" => data_out <= rom_array(41064);
		when "1010000001101001" => data_out <= rom_array(41065);
		when "1010000001101010" => data_out <= rom_array(41066);
		when "1010000001101011" => data_out <= rom_array(41067);
		when "1010000001101100" => data_out <= rom_array(41068);
		when "1010000001101101" => data_out <= rom_array(41069);
		when "1010000001101110" => data_out <= rom_array(41070);
		when "1010000001101111" => data_out <= rom_array(41071);
		when "1010000001110000" => data_out <= rom_array(41072);
		when "1010000001110001" => data_out <= rom_array(41073);
		when "1010000001110010" => data_out <= rom_array(41074);
		when "1010000001110011" => data_out <= rom_array(41075);
		when "1010000001110100" => data_out <= rom_array(41076);
		when "1010000001110101" => data_out <= rom_array(41077);
		when "1010000001110110" => data_out <= rom_array(41078);
		when "1010000001110111" => data_out <= rom_array(41079);
		when "1010000001111000" => data_out <= rom_array(41080);
		when "1010000001111001" => data_out <= rom_array(41081);
		when "1010000001111010" => data_out <= rom_array(41082);
		when "1010000001111011" => data_out <= rom_array(41083);
		when "1010000001111100" => data_out <= rom_array(41084);
		when "1010000001111101" => data_out <= rom_array(41085);
		when "1010000001111110" => data_out <= rom_array(41086);
		when "1010000001111111" => data_out <= rom_array(41087);
		when "1010000010000000" => data_out <= rom_array(41088);
		when "1010000010000001" => data_out <= rom_array(41089);
		when "1010000010000010" => data_out <= rom_array(41090);
		when "1010000010000011" => data_out <= rom_array(41091);
		when "1010000010000100" => data_out <= rom_array(41092);
		when "1010000010000101" => data_out <= rom_array(41093);
		when "1010000010000110" => data_out <= rom_array(41094);
		when "1010000010000111" => data_out <= rom_array(41095);
		when "1010000010001000" => data_out <= rom_array(41096);
		when "1010000010001001" => data_out <= rom_array(41097);
		when "1010000010001010" => data_out <= rom_array(41098);
		when "1010000010001011" => data_out <= rom_array(41099);
		when "1010000010001100" => data_out <= rom_array(41100);
		when "1010000010001101" => data_out <= rom_array(41101);
		when "1010000010001110" => data_out <= rom_array(41102);
		when "1010000010001111" => data_out <= rom_array(41103);
		when "1010000010010000" => data_out <= rom_array(41104);
		when "1010000010010001" => data_out <= rom_array(41105);
		when "1010000010010010" => data_out <= rom_array(41106);
		when "1010000010010011" => data_out <= rom_array(41107);
		when "1010000010010100" => data_out <= rom_array(41108);
		when "1010000010010101" => data_out <= rom_array(41109);
		when "1010000010010110" => data_out <= rom_array(41110);
		when "1010000010010111" => data_out <= rom_array(41111);
		when "1010000010011000" => data_out <= rom_array(41112);
		when "1010000010011001" => data_out <= rom_array(41113);
		when "1010000010011010" => data_out <= rom_array(41114);
		when "1010000010011011" => data_out <= rom_array(41115);
		when "1010000010011100" => data_out <= rom_array(41116);
		when "1010000010011101" => data_out <= rom_array(41117);
		when "1010000010011110" => data_out <= rom_array(41118);
		when "1010000010011111" => data_out <= rom_array(41119);
		when "1010000010100000" => data_out <= rom_array(41120);
		when "1010000010100001" => data_out <= rom_array(41121);
		when "1010000010100010" => data_out <= rom_array(41122);
		when "1010000010100011" => data_out <= rom_array(41123);
		when "1010000010100100" => data_out <= rom_array(41124);
		when "1010000010100101" => data_out <= rom_array(41125);
		when "1010000010100110" => data_out <= rom_array(41126);
		when "1010000010100111" => data_out <= rom_array(41127);
		when "1010000010101000" => data_out <= rom_array(41128);
		when "1010000010101001" => data_out <= rom_array(41129);
		when "1010000010101010" => data_out <= rom_array(41130);
		when "1010000010101011" => data_out <= rom_array(41131);
		when "1010000010101100" => data_out <= rom_array(41132);
		when "1010000010101101" => data_out <= rom_array(41133);
		when "1010000010101110" => data_out <= rom_array(41134);
		when "1010000010101111" => data_out <= rom_array(41135);
		when "1010000010110000" => data_out <= rom_array(41136);
		when "1010000010110001" => data_out <= rom_array(41137);
		when "1010000010110010" => data_out <= rom_array(41138);
		when "1010000010110011" => data_out <= rom_array(41139);
		when "1010000010110100" => data_out <= rom_array(41140);
		when "1010000010110101" => data_out <= rom_array(41141);
		when "1010000010110110" => data_out <= rom_array(41142);
		when "1010000010110111" => data_out <= rom_array(41143);
		when "1010000010111000" => data_out <= rom_array(41144);
		when "1010000010111001" => data_out <= rom_array(41145);
		when "1010000010111010" => data_out <= rom_array(41146);
		when "1010000010111011" => data_out <= rom_array(41147);
		when "1010000010111100" => data_out <= rom_array(41148);
		when "1010000010111101" => data_out <= rom_array(41149);
		when "1010000010111110" => data_out <= rom_array(41150);
		when "1010000010111111" => data_out <= rom_array(41151);
		when "1010000011000000" => data_out <= rom_array(41152);
		when "1010000011000001" => data_out <= rom_array(41153);
		when "1010000011000010" => data_out <= rom_array(41154);
		when "1010000011000011" => data_out <= rom_array(41155);
		when "1010000011000100" => data_out <= rom_array(41156);
		when "1010000011000101" => data_out <= rom_array(41157);
		when "1010000011000110" => data_out <= rom_array(41158);
		when "1010000011000111" => data_out <= rom_array(41159);
		when "1010000011001000" => data_out <= rom_array(41160);
		when "1010000011001001" => data_out <= rom_array(41161);
		when "1010000011001010" => data_out <= rom_array(41162);
		when "1010000011001011" => data_out <= rom_array(41163);
		when "1010000011001100" => data_out <= rom_array(41164);
		when "1010000011001101" => data_out <= rom_array(41165);
		when "1010000011001110" => data_out <= rom_array(41166);
		when "1010000011001111" => data_out <= rom_array(41167);
		when "1010000011010000" => data_out <= rom_array(41168);
		when "1010000011010001" => data_out <= rom_array(41169);
		when "1010000011010010" => data_out <= rom_array(41170);
		when "1010000011010011" => data_out <= rom_array(41171);
		when "1010000011010100" => data_out <= rom_array(41172);
		when "1010000011010101" => data_out <= rom_array(41173);
		when "1010000011010110" => data_out <= rom_array(41174);
		when "1010000011010111" => data_out <= rom_array(41175);
		when "1010000011011000" => data_out <= rom_array(41176);
		when "1010000011011001" => data_out <= rom_array(41177);
		when "1010000011011010" => data_out <= rom_array(41178);
		when "1010000011011011" => data_out <= rom_array(41179);
		when "1010000011011100" => data_out <= rom_array(41180);
		when "1010000011011101" => data_out <= rom_array(41181);
		when "1010000011011110" => data_out <= rom_array(41182);
		when "1010000011011111" => data_out <= rom_array(41183);
		when "1010000011100000" => data_out <= rom_array(41184);
		when "1010000011100001" => data_out <= rom_array(41185);
		when "1010000011100010" => data_out <= rom_array(41186);
		when "1010000011100011" => data_out <= rom_array(41187);
		when "1010000011100100" => data_out <= rom_array(41188);
		when "1010000011100101" => data_out <= rom_array(41189);
		when "1010000011100110" => data_out <= rom_array(41190);
		when "1010000011100111" => data_out <= rom_array(41191);
		when "1010000011101000" => data_out <= rom_array(41192);
		when "1010000011101001" => data_out <= rom_array(41193);
		when "1010000011101010" => data_out <= rom_array(41194);
		when "1010000011101011" => data_out <= rom_array(41195);
		when "1010000011101100" => data_out <= rom_array(41196);
		when "1010000011101101" => data_out <= rom_array(41197);
		when "1010000011101110" => data_out <= rom_array(41198);
		when "1010000011101111" => data_out <= rom_array(41199);
		when "1010000011110000" => data_out <= rom_array(41200);
		when "1010000011110001" => data_out <= rom_array(41201);
		when "1010000011110010" => data_out <= rom_array(41202);
		when "1010000011110011" => data_out <= rom_array(41203);
		when "1010000011110100" => data_out <= rom_array(41204);
		when "1010000011110101" => data_out <= rom_array(41205);
		when "1010000011110110" => data_out <= rom_array(41206);
		when "1010000011110111" => data_out <= rom_array(41207);
		when "1010000011111000" => data_out <= rom_array(41208);
		when "1010000011111001" => data_out <= rom_array(41209);
		when "1010000011111010" => data_out <= rom_array(41210);
		when "1010000011111011" => data_out <= rom_array(41211);
		when "1010000011111100" => data_out <= rom_array(41212);
		when "1010000011111101" => data_out <= rom_array(41213);
		when "1010000011111110" => data_out <= rom_array(41214);
		when "1010000011111111" => data_out <= rom_array(41215);
		when "1010000100000000" => data_out <= rom_array(41216);
		when "1010000100000001" => data_out <= rom_array(41217);
		when "1010000100000010" => data_out <= rom_array(41218);
		when "1010000100000011" => data_out <= rom_array(41219);
		when "1010000100000100" => data_out <= rom_array(41220);
		when "1010000100000101" => data_out <= rom_array(41221);
		when "1010000100000110" => data_out <= rom_array(41222);
		when "1010000100000111" => data_out <= rom_array(41223);
		when "1010000100001000" => data_out <= rom_array(41224);
		when "1010000100001001" => data_out <= rom_array(41225);
		when "1010000100001010" => data_out <= rom_array(41226);
		when "1010000100001011" => data_out <= rom_array(41227);
		when "1010000100001100" => data_out <= rom_array(41228);
		when "1010000100001101" => data_out <= rom_array(41229);
		when "1010000100001110" => data_out <= rom_array(41230);
		when "1010000100001111" => data_out <= rom_array(41231);
		when "1010000100010000" => data_out <= rom_array(41232);
		when "1010000100010001" => data_out <= rom_array(41233);
		when "1010000100010010" => data_out <= rom_array(41234);
		when "1010000100010011" => data_out <= rom_array(41235);
		when "1010000100010100" => data_out <= rom_array(41236);
		when "1010000100010101" => data_out <= rom_array(41237);
		when "1010000100010110" => data_out <= rom_array(41238);
		when "1010000100010111" => data_out <= rom_array(41239);
		when "1010000100011000" => data_out <= rom_array(41240);
		when "1010000100011001" => data_out <= rom_array(41241);
		when "1010000100011010" => data_out <= rom_array(41242);
		when "1010000100011011" => data_out <= rom_array(41243);
		when "1010000100011100" => data_out <= rom_array(41244);
		when "1010000100011101" => data_out <= rom_array(41245);
		when "1010000100011110" => data_out <= rom_array(41246);
		when "1010000100011111" => data_out <= rom_array(41247);
		when "1010000100100000" => data_out <= rom_array(41248);
		when "1010000100100001" => data_out <= rom_array(41249);
		when "1010000100100010" => data_out <= rom_array(41250);
		when "1010000100100011" => data_out <= rom_array(41251);
		when "1010000100100100" => data_out <= rom_array(41252);
		when "1010000100100101" => data_out <= rom_array(41253);
		when "1010000100100110" => data_out <= rom_array(41254);
		when "1010000100100111" => data_out <= rom_array(41255);
		when "1010000100101000" => data_out <= rom_array(41256);
		when "1010000100101001" => data_out <= rom_array(41257);
		when "1010000100101010" => data_out <= rom_array(41258);
		when "1010000100101011" => data_out <= rom_array(41259);
		when "1010000100101100" => data_out <= rom_array(41260);
		when "1010000100101101" => data_out <= rom_array(41261);
		when "1010000100101110" => data_out <= rom_array(41262);
		when "1010000100101111" => data_out <= rom_array(41263);
		when "1010000100110000" => data_out <= rom_array(41264);
		when "1010000100110001" => data_out <= rom_array(41265);
		when "1010000100110010" => data_out <= rom_array(41266);
		when "1010000100110011" => data_out <= rom_array(41267);
		when "1010000100110100" => data_out <= rom_array(41268);
		when "1010000100110101" => data_out <= rom_array(41269);
		when "1010000100110110" => data_out <= rom_array(41270);
		when "1010000100110111" => data_out <= rom_array(41271);
		when "1010000100111000" => data_out <= rom_array(41272);
		when "1010000100111001" => data_out <= rom_array(41273);
		when "1010000100111010" => data_out <= rom_array(41274);
		when "1010000100111011" => data_out <= rom_array(41275);
		when "1010000100111100" => data_out <= rom_array(41276);
		when "1010000100111101" => data_out <= rom_array(41277);
		when "1010000100111110" => data_out <= rom_array(41278);
		when "1010000100111111" => data_out <= rom_array(41279);
		when "1010000101000000" => data_out <= rom_array(41280);
		when "1010000101000001" => data_out <= rom_array(41281);
		when "1010000101000010" => data_out <= rom_array(41282);
		when "1010000101000011" => data_out <= rom_array(41283);
		when "1010000101000100" => data_out <= rom_array(41284);
		when "1010000101000101" => data_out <= rom_array(41285);
		when "1010000101000110" => data_out <= rom_array(41286);
		when "1010000101000111" => data_out <= rom_array(41287);
		when "1010000101001000" => data_out <= rom_array(41288);
		when "1010000101001001" => data_out <= rom_array(41289);
		when "1010000101001010" => data_out <= rom_array(41290);
		when "1010000101001011" => data_out <= rom_array(41291);
		when "1010000101001100" => data_out <= rom_array(41292);
		when "1010000101001101" => data_out <= rom_array(41293);
		when "1010000101001110" => data_out <= rom_array(41294);
		when "1010000101001111" => data_out <= rom_array(41295);
		when "1010000101010000" => data_out <= rom_array(41296);
		when "1010000101010001" => data_out <= rom_array(41297);
		when "1010000101010010" => data_out <= rom_array(41298);
		when "1010000101010011" => data_out <= rom_array(41299);
		when "1010000101010100" => data_out <= rom_array(41300);
		when "1010000101010101" => data_out <= rom_array(41301);
		when "1010000101010110" => data_out <= rom_array(41302);
		when "1010000101010111" => data_out <= rom_array(41303);
		when "1010000101011000" => data_out <= rom_array(41304);
		when "1010000101011001" => data_out <= rom_array(41305);
		when "1010000101011010" => data_out <= rom_array(41306);
		when "1010000101011011" => data_out <= rom_array(41307);
		when "1010000101011100" => data_out <= rom_array(41308);
		when "1010000101011101" => data_out <= rom_array(41309);
		when "1010000101011110" => data_out <= rom_array(41310);
		when "1010000101011111" => data_out <= rom_array(41311);
		when "1010000101100000" => data_out <= rom_array(41312);
		when "1010000101100001" => data_out <= rom_array(41313);
		when "1010000101100010" => data_out <= rom_array(41314);
		when "1010000101100011" => data_out <= rom_array(41315);
		when "1010000101100100" => data_out <= rom_array(41316);
		when "1010000101100101" => data_out <= rom_array(41317);
		when "1010000101100110" => data_out <= rom_array(41318);
		when "1010000101100111" => data_out <= rom_array(41319);
		when "1010000101101000" => data_out <= rom_array(41320);
		when "1010000101101001" => data_out <= rom_array(41321);
		when "1010000101101010" => data_out <= rom_array(41322);
		when "1010000101101011" => data_out <= rom_array(41323);
		when "1010000101101100" => data_out <= rom_array(41324);
		when "1010000101101101" => data_out <= rom_array(41325);
		when "1010000101101110" => data_out <= rom_array(41326);
		when "1010000101101111" => data_out <= rom_array(41327);
		when "1010000101110000" => data_out <= rom_array(41328);
		when "1010000101110001" => data_out <= rom_array(41329);
		when "1010000101110010" => data_out <= rom_array(41330);
		when "1010000101110011" => data_out <= rom_array(41331);
		when "1010000101110100" => data_out <= rom_array(41332);
		when "1010000101110101" => data_out <= rom_array(41333);
		when "1010000101110110" => data_out <= rom_array(41334);
		when "1010000101110111" => data_out <= rom_array(41335);
		when "1010000101111000" => data_out <= rom_array(41336);
		when "1010000101111001" => data_out <= rom_array(41337);
		when "1010000101111010" => data_out <= rom_array(41338);
		when "1010000101111011" => data_out <= rom_array(41339);
		when "1010000101111100" => data_out <= rom_array(41340);
		when "1010000101111101" => data_out <= rom_array(41341);
		when "1010000101111110" => data_out <= rom_array(41342);
		when "1010000101111111" => data_out <= rom_array(41343);
		when "1010000110000000" => data_out <= rom_array(41344);
		when "1010000110000001" => data_out <= rom_array(41345);
		when "1010000110000010" => data_out <= rom_array(41346);
		when "1010000110000011" => data_out <= rom_array(41347);
		when "1010000110000100" => data_out <= rom_array(41348);
		when "1010000110000101" => data_out <= rom_array(41349);
		when "1010000110000110" => data_out <= rom_array(41350);
		when "1010000110000111" => data_out <= rom_array(41351);
		when "1010000110001000" => data_out <= rom_array(41352);
		when "1010000110001001" => data_out <= rom_array(41353);
		when "1010000110001010" => data_out <= rom_array(41354);
		when "1010000110001011" => data_out <= rom_array(41355);
		when "1010000110001100" => data_out <= rom_array(41356);
		when "1010000110001101" => data_out <= rom_array(41357);
		when "1010000110001110" => data_out <= rom_array(41358);
		when "1010000110001111" => data_out <= rom_array(41359);
		when "1010000110010000" => data_out <= rom_array(41360);
		when "1010000110010001" => data_out <= rom_array(41361);
		when "1010000110010010" => data_out <= rom_array(41362);
		when "1010000110010011" => data_out <= rom_array(41363);
		when "1010000110010100" => data_out <= rom_array(41364);
		when "1010000110010101" => data_out <= rom_array(41365);
		when "1010000110010110" => data_out <= rom_array(41366);
		when "1010000110010111" => data_out <= rom_array(41367);
		when "1010000110011000" => data_out <= rom_array(41368);
		when "1010000110011001" => data_out <= rom_array(41369);
		when "1010000110011010" => data_out <= rom_array(41370);
		when "1010000110011011" => data_out <= rom_array(41371);
		when "1010000110011100" => data_out <= rom_array(41372);
		when "1010000110011101" => data_out <= rom_array(41373);
		when "1010000110011110" => data_out <= rom_array(41374);
		when "1010000110011111" => data_out <= rom_array(41375);
		when "1010000110100000" => data_out <= rom_array(41376);
		when "1010000110100001" => data_out <= rom_array(41377);
		when "1010000110100010" => data_out <= rom_array(41378);
		when "1010000110100011" => data_out <= rom_array(41379);
		when "1010000110100100" => data_out <= rom_array(41380);
		when "1010000110100101" => data_out <= rom_array(41381);
		when "1010000110100110" => data_out <= rom_array(41382);
		when "1010000110100111" => data_out <= rom_array(41383);
		when "1010000110101000" => data_out <= rom_array(41384);
		when "1010000110101001" => data_out <= rom_array(41385);
		when "1010000110101010" => data_out <= rom_array(41386);
		when "1010000110101011" => data_out <= rom_array(41387);
		when "1010000110101100" => data_out <= rom_array(41388);
		when "1010000110101101" => data_out <= rom_array(41389);
		when "1010000110101110" => data_out <= rom_array(41390);
		when "1010000110101111" => data_out <= rom_array(41391);
		when "1010000110110000" => data_out <= rom_array(41392);
		when "1010000110110001" => data_out <= rom_array(41393);
		when "1010000110110010" => data_out <= rom_array(41394);
		when "1010000110110011" => data_out <= rom_array(41395);
		when "1010000110110100" => data_out <= rom_array(41396);
		when "1010000110110101" => data_out <= rom_array(41397);
		when "1010000110110110" => data_out <= rom_array(41398);
		when "1010000110110111" => data_out <= rom_array(41399);
		when "1010000110111000" => data_out <= rom_array(41400);
		when "1010000110111001" => data_out <= rom_array(41401);
		when "1010000110111010" => data_out <= rom_array(41402);
		when "1010000110111011" => data_out <= rom_array(41403);
		when "1010000110111100" => data_out <= rom_array(41404);
		when "1010000110111101" => data_out <= rom_array(41405);
		when "1010000110111110" => data_out <= rom_array(41406);
		when "1010000110111111" => data_out <= rom_array(41407);
		when "1010000111000000" => data_out <= rom_array(41408);
		when "1010000111000001" => data_out <= rom_array(41409);
		when "1010000111000010" => data_out <= rom_array(41410);
		when "1010000111000011" => data_out <= rom_array(41411);
		when "1010000111000100" => data_out <= rom_array(41412);
		when "1010000111000101" => data_out <= rom_array(41413);
		when "1010000111000110" => data_out <= rom_array(41414);
		when "1010000111000111" => data_out <= rom_array(41415);
		when "1010000111001000" => data_out <= rom_array(41416);
		when "1010000111001001" => data_out <= rom_array(41417);
		when "1010000111001010" => data_out <= rom_array(41418);
		when "1010000111001011" => data_out <= rom_array(41419);
		when "1010000111001100" => data_out <= rom_array(41420);
		when "1010000111001101" => data_out <= rom_array(41421);
		when "1010000111001110" => data_out <= rom_array(41422);
		when "1010000111001111" => data_out <= rom_array(41423);
		when "1010000111010000" => data_out <= rom_array(41424);
		when "1010000111010001" => data_out <= rom_array(41425);
		when "1010000111010010" => data_out <= rom_array(41426);
		when "1010000111010011" => data_out <= rom_array(41427);
		when "1010000111010100" => data_out <= rom_array(41428);
		when "1010000111010101" => data_out <= rom_array(41429);
		when "1010000111010110" => data_out <= rom_array(41430);
		when "1010000111010111" => data_out <= rom_array(41431);
		when "1010000111011000" => data_out <= rom_array(41432);
		when "1010000111011001" => data_out <= rom_array(41433);
		when "1010000111011010" => data_out <= rom_array(41434);
		when "1010000111011011" => data_out <= rom_array(41435);
		when "1010000111011100" => data_out <= rom_array(41436);
		when "1010000111011101" => data_out <= rom_array(41437);
		when "1010000111011110" => data_out <= rom_array(41438);
		when "1010000111011111" => data_out <= rom_array(41439);
		when "1010000111100000" => data_out <= rom_array(41440);
		when "1010000111100001" => data_out <= rom_array(41441);
		when "1010000111100010" => data_out <= rom_array(41442);
		when "1010000111100011" => data_out <= rom_array(41443);
		when "1010000111100100" => data_out <= rom_array(41444);
		when "1010000111100101" => data_out <= rom_array(41445);
		when "1010000111100110" => data_out <= rom_array(41446);
		when "1010000111100111" => data_out <= rom_array(41447);
		when "1010000111101000" => data_out <= rom_array(41448);
		when "1010000111101001" => data_out <= rom_array(41449);
		when "1010000111101010" => data_out <= rom_array(41450);
		when "1010000111101011" => data_out <= rom_array(41451);
		when "1010000111101100" => data_out <= rom_array(41452);
		when "1010000111101101" => data_out <= rom_array(41453);
		when "1010000111101110" => data_out <= rom_array(41454);
		when "1010000111101111" => data_out <= rom_array(41455);
		when "1010000111110000" => data_out <= rom_array(41456);
		when "1010000111110001" => data_out <= rom_array(41457);
		when "1010000111110010" => data_out <= rom_array(41458);
		when "1010000111110011" => data_out <= rom_array(41459);
		when "1010000111110100" => data_out <= rom_array(41460);
		when "1010000111110101" => data_out <= rom_array(41461);
		when "1010000111110110" => data_out <= rom_array(41462);
		when "1010000111110111" => data_out <= rom_array(41463);
		when "1010000111111000" => data_out <= rom_array(41464);
		when "1010000111111001" => data_out <= rom_array(41465);
		when "1010000111111010" => data_out <= rom_array(41466);
		when "1010000111111011" => data_out <= rom_array(41467);
		when "1010000111111100" => data_out <= rom_array(41468);
		when "1010000111111101" => data_out <= rom_array(41469);
		when "1010000111111110" => data_out <= rom_array(41470);
		when "1010000111111111" => data_out <= rom_array(41471);
		when "1010001000000000" => data_out <= rom_array(41472);
		when "1010001000000001" => data_out <= rom_array(41473);
		when "1010001000000010" => data_out <= rom_array(41474);
		when "1010001000000011" => data_out <= rom_array(41475);
		when "1010001000000100" => data_out <= rom_array(41476);
		when "1010001000000101" => data_out <= rom_array(41477);
		when "1010001000000110" => data_out <= rom_array(41478);
		when "1010001000000111" => data_out <= rom_array(41479);
		when "1010001000001000" => data_out <= rom_array(41480);
		when "1010001000001001" => data_out <= rom_array(41481);
		when "1010001000001010" => data_out <= rom_array(41482);
		when "1010001000001011" => data_out <= rom_array(41483);
		when "1010001000001100" => data_out <= rom_array(41484);
		when "1010001000001101" => data_out <= rom_array(41485);
		when "1010001000001110" => data_out <= rom_array(41486);
		when "1010001000001111" => data_out <= rom_array(41487);
		when "1010001000010000" => data_out <= rom_array(41488);
		when "1010001000010001" => data_out <= rom_array(41489);
		when "1010001000010010" => data_out <= rom_array(41490);
		when "1010001000010011" => data_out <= rom_array(41491);
		when "1010001000010100" => data_out <= rom_array(41492);
		when "1010001000010101" => data_out <= rom_array(41493);
		when "1010001000010110" => data_out <= rom_array(41494);
		when "1010001000010111" => data_out <= rom_array(41495);
		when "1010001000011000" => data_out <= rom_array(41496);
		when "1010001000011001" => data_out <= rom_array(41497);
		when "1010001000011010" => data_out <= rom_array(41498);
		when "1010001000011011" => data_out <= rom_array(41499);
		when "1010001000011100" => data_out <= rom_array(41500);
		when "1010001000011101" => data_out <= rom_array(41501);
		when "1010001000011110" => data_out <= rom_array(41502);
		when "1010001000011111" => data_out <= rom_array(41503);
		when "1010001000100000" => data_out <= rom_array(41504);
		when "1010001000100001" => data_out <= rom_array(41505);
		when "1010001000100010" => data_out <= rom_array(41506);
		when "1010001000100011" => data_out <= rom_array(41507);
		when "1010001000100100" => data_out <= rom_array(41508);
		when "1010001000100101" => data_out <= rom_array(41509);
		when "1010001000100110" => data_out <= rom_array(41510);
		when "1010001000100111" => data_out <= rom_array(41511);
		when "1010001000101000" => data_out <= rom_array(41512);
		when "1010001000101001" => data_out <= rom_array(41513);
		when "1010001000101010" => data_out <= rom_array(41514);
		when "1010001000101011" => data_out <= rom_array(41515);
		when "1010001000101100" => data_out <= rom_array(41516);
		when "1010001000101101" => data_out <= rom_array(41517);
		when "1010001000101110" => data_out <= rom_array(41518);
		when "1010001000101111" => data_out <= rom_array(41519);
		when "1010001000110000" => data_out <= rom_array(41520);
		when "1010001000110001" => data_out <= rom_array(41521);
		when "1010001000110010" => data_out <= rom_array(41522);
		when "1010001000110011" => data_out <= rom_array(41523);
		when "1010001000110100" => data_out <= rom_array(41524);
		when "1010001000110101" => data_out <= rom_array(41525);
		when "1010001000110110" => data_out <= rom_array(41526);
		when "1010001000110111" => data_out <= rom_array(41527);
		when "1010001000111000" => data_out <= rom_array(41528);
		when "1010001000111001" => data_out <= rom_array(41529);
		when "1010001000111010" => data_out <= rom_array(41530);
		when "1010001000111011" => data_out <= rom_array(41531);
		when "1010001000111100" => data_out <= rom_array(41532);
		when "1010001000111101" => data_out <= rom_array(41533);
		when "1010001000111110" => data_out <= rom_array(41534);
		when "1010001000111111" => data_out <= rom_array(41535);
		when "1010001001000000" => data_out <= rom_array(41536);
		when "1010001001000001" => data_out <= rom_array(41537);
		when "1010001001000010" => data_out <= rom_array(41538);
		when "1010001001000011" => data_out <= rom_array(41539);
		when "1010001001000100" => data_out <= rom_array(41540);
		when "1010001001000101" => data_out <= rom_array(41541);
		when "1010001001000110" => data_out <= rom_array(41542);
		when "1010001001000111" => data_out <= rom_array(41543);
		when "1010001001001000" => data_out <= rom_array(41544);
		when "1010001001001001" => data_out <= rom_array(41545);
		when "1010001001001010" => data_out <= rom_array(41546);
		when "1010001001001011" => data_out <= rom_array(41547);
		when "1010001001001100" => data_out <= rom_array(41548);
		when "1010001001001101" => data_out <= rom_array(41549);
		when "1010001001001110" => data_out <= rom_array(41550);
		when "1010001001001111" => data_out <= rom_array(41551);
		when "1010001001010000" => data_out <= rom_array(41552);
		when "1010001001010001" => data_out <= rom_array(41553);
		when "1010001001010010" => data_out <= rom_array(41554);
		when "1010001001010011" => data_out <= rom_array(41555);
		when "1010001001010100" => data_out <= rom_array(41556);
		when "1010001001010101" => data_out <= rom_array(41557);
		when "1010001001010110" => data_out <= rom_array(41558);
		when "1010001001010111" => data_out <= rom_array(41559);
		when "1010001001011000" => data_out <= rom_array(41560);
		when "1010001001011001" => data_out <= rom_array(41561);
		when "1010001001011010" => data_out <= rom_array(41562);
		when "1010001001011011" => data_out <= rom_array(41563);
		when "1010001001011100" => data_out <= rom_array(41564);
		when "1010001001011101" => data_out <= rom_array(41565);
		when "1010001001011110" => data_out <= rom_array(41566);
		when "1010001001011111" => data_out <= rom_array(41567);
		when "1010001001100000" => data_out <= rom_array(41568);
		when "1010001001100001" => data_out <= rom_array(41569);
		when "1010001001100010" => data_out <= rom_array(41570);
		when "1010001001100011" => data_out <= rom_array(41571);
		when "1010001001100100" => data_out <= rom_array(41572);
		when "1010001001100101" => data_out <= rom_array(41573);
		when "1010001001100110" => data_out <= rom_array(41574);
		when "1010001001100111" => data_out <= rom_array(41575);
		when "1010001001101000" => data_out <= rom_array(41576);
		when "1010001001101001" => data_out <= rom_array(41577);
		when "1010001001101010" => data_out <= rom_array(41578);
		when "1010001001101011" => data_out <= rom_array(41579);
		when "1010001001101100" => data_out <= rom_array(41580);
		when "1010001001101101" => data_out <= rom_array(41581);
		when "1010001001101110" => data_out <= rom_array(41582);
		when "1010001001101111" => data_out <= rom_array(41583);
		when "1010001001110000" => data_out <= rom_array(41584);
		when "1010001001110001" => data_out <= rom_array(41585);
		when "1010001001110010" => data_out <= rom_array(41586);
		when "1010001001110011" => data_out <= rom_array(41587);
		when "1010001001110100" => data_out <= rom_array(41588);
		when "1010001001110101" => data_out <= rom_array(41589);
		when "1010001001110110" => data_out <= rom_array(41590);
		when "1010001001110111" => data_out <= rom_array(41591);
		when "1010001001111000" => data_out <= rom_array(41592);
		when "1010001001111001" => data_out <= rom_array(41593);
		when "1010001001111010" => data_out <= rom_array(41594);
		when "1010001001111011" => data_out <= rom_array(41595);
		when "1010001001111100" => data_out <= rom_array(41596);
		when "1010001001111101" => data_out <= rom_array(41597);
		when "1010001001111110" => data_out <= rom_array(41598);
		when "1010001001111111" => data_out <= rom_array(41599);
		when "1010001010000000" => data_out <= rom_array(41600);
		when "1010001010000001" => data_out <= rom_array(41601);
		when "1010001010000010" => data_out <= rom_array(41602);
		when "1010001010000011" => data_out <= rom_array(41603);
		when "1010001010000100" => data_out <= rom_array(41604);
		when "1010001010000101" => data_out <= rom_array(41605);
		when "1010001010000110" => data_out <= rom_array(41606);
		when "1010001010000111" => data_out <= rom_array(41607);
		when "1010001010001000" => data_out <= rom_array(41608);
		when "1010001010001001" => data_out <= rom_array(41609);
		when "1010001010001010" => data_out <= rom_array(41610);
		when "1010001010001011" => data_out <= rom_array(41611);
		when "1010001010001100" => data_out <= rom_array(41612);
		when "1010001010001101" => data_out <= rom_array(41613);
		when "1010001010001110" => data_out <= rom_array(41614);
		when "1010001010001111" => data_out <= rom_array(41615);
		when "1010001010010000" => data_out <= rom_array(41616);
		when "1010001010010001" => data_out <= rom_array(41617);
		when "1010001010010010" => data_out <= rom_array(41618);
		when "1010001010010011" => data_out <= rom_array(41619);
		when "1010001010010100" => data_out <= rom_array(41620);
		when "1010001010010101" => data_out <= rom_array(41621);
		when "1010001010010110" => data_out <= rom_array(41622);
		when "1010001010010111" => data_out <= rom_array(41623);
		when "1010001010011000" => data_out <= rom_array(41624);
		when "1010001010011001" => data_out <= rom_array(41625);
		when "1010001010011010" => data_out <= rom_array(41626);
		when "1010001010011011" => data_out <= rom_array(41627);
		when "1010001010011100" => data_out <= rom_array(41628);
		when "1010001010011101" => data_out <= rom_array(41629);
		when "1010001010011110" => data_out <= rom_array(41630);
		when "1010001010011111" => data_out <= rom_array(41631);
		when "1010001010100000" => data_out <= rom_array(41632);
		when "1010001010100001" => data_out <= rom_array(41633);
		when "1010001010100010" => data_out <= rom_array(41634);
		when "1010001010100011" => data_out <= rom_array(41635);
		when "1010001010100100" => data_out <= rom_array(41636);
		when "1010001010100101" => data_out <= rom_array(41637);
		when "1010001010100110" => data_out <= rom_array(41638);
		when "1010001010100111" => data_out <= rom_array(41639);
		when "1010001010101000" => data_out <= rom_array(41640);
		when "1010001010101001" => data_out <= rom_array(41641);
		when "1010001010101010" => data_out <= rom_array(41642);
		when "1010001010101011" => data_out <= rom_array(41643);
		when "1010001010101100" => data_out <= rom_array(41644);
		when "1010001010101101" => data_out <= rom_array(41645);
		when "1010001010101110" => data_out <= rom_array(41646);
		when "1010001010101111" => data_out <= rom_array(41647);
		when "1010001010110000" => data_out <= rom_array(41648);
		when "1010001010110001" => data_out <= rom_array(41649);
		when "1010001010110010" => data_out <= rom_array(41650);
		when "1010001010110011" => data_out <= rom_array(41651);
		when "1010001010110100" => data_out <= rom_array(41652);
		when "1010001010110101" => data_out <= rom_array(41653);
		when "1010001010110110" => data_out <= rom_array(41654);
		when "1010001010110111" => data_out <= rom_array(41655);
		when "1010001010111000" => data_out <= rom_array(41656);
		when "1010001010111001" => data_out <= rom_array(41657);
		when "1010001010111010" => data_out <= rom_array(41658);
		when "1010001010111011" => data_out <= rom_array(41659);
		when "1010001010111100" => data_out <= rom_array(41660);
		when "1010001010111101" => data_out <= rom_array(41661);
		when "1010001010111110" => data_out <= rom_array(41662);
		when "1010001010111111" => data_out <= rom_array(41663);
		when "1010001011000000" => data_out <= rom_array(41664);
		when "1010001011000001" => data_out <= rom_array(41665);
		when "1010001011000010" => data_out <= rom_array(41666);
		when "1010001011000011" => data_out <= rom_array(41667);
		when "1010001011000100" => data_out <= rom_array(41668);
		when "1010001011000101" => data_out <= rom_array(41669);
		when "1010001011000110" => data_out <= rom_array(41670);
		when "1010001011000111" => data_out <= rom_array(41671);
		when "1010001011001000" => data_out <= rom_array(41672);
		when "1010001011001001" => data_out <= rom_array(41673);
		when "1010001011001010" => data_out <= rom_array(41674);
		when "1010001011001011" => data_out <= rom_array(41675);
		when "1010001011001100" => data_out <= rom_array(41676);
		when "1010001011001101" => data_out <= rom_array(41677);
		when "1010001011001110" => data_out <= rom_array(41678);
		when "1010001011001111" => data_out <= rom_array(41679);
		when "1010001011010000" => data_out <= rom_array(41680);
		when "1010001011010001" => data_out <= rom_array(41681);
		when "1010001011010010" => data_out <= rom_array(41682);
		when "1010001011010011" => data_out <= rom_array(41683);
		when "1010001011010100" => data_out <= rom_array(41684);
		when "1010001011010101" => data_out <= rom_array(41685);
		when "1010001011010110" => data_out <= rom_array(41686);
		when "1010001011010111" => data_out <= rom_array(41687);
		when "1010001011011000" => data_out <= rom_array(41688);
		when "1010001011011001" => data_out <= rom_array(41689);
		when "1010001011011010" => data_out <= rom_array(41690);
		when "1010001011011011" => data_out <= rom_array(41691);
		when "1010001011011100" => data_out <= rom_array(41692);
		when "1010001011011101" => data_out <= rom_array(41693);
		when "1010001011011110" => data_out <= rom_array(41694);
		when "1010001011011111" => data_out <= rom_array(41695);
		when "1010001011100000" => data_out <= rom_array(41696);
		when "1010001011100001" => data_out <= rom_array(41697);
		when "1010001011100010" => data_out <= rom_array(41698);
		when "1010001011100011" => data_out <= rom_array(41699);
		when "1010001011100100" => data_out <= rom_array(41700);
		when "1010001011100101" => data_out <= rom_array(41701);
		when "1010001011100110" => data_out <= rom_array(41702);
		when "1010001011100111" => data_out <= rom_array(41703);
		when "1010001011101000" => data_out <= rom_array(41704);
		when "1010001011101001" => data_out <= rom_array(41705);
		when "1010001011101010" => data_out <= rom_array(41706);
		when "1010001011101011" => data_out <= rom_array(41707);
		when "1010001011101100" => data_out <= rom_array(41708);
		when "1010001011101101" => data_out <= rom_array(41709);
		when "1010001011101110" => data_out <= rom_array(41710);
		when "1010001011101111" => data_out <= rom_array(41711);
		when "1010001011110000" => data_out <= rom_array(41712);
		when "1010001011110001" => data_out <= rom_array(41713);
		when "1010001011110010" => data_out <= rom_array(41714);
		when "1010001011110011" => data_out <= rom_array(41715);
		when "1010001011110100" => data_out <= rom_array(41716);
		when "1010001011110101" => data_out <= rom_array(41717);
		when "1010001011110110" => data_out <= rom_array(41718);
		when "1010001011110111" => data_out <= rom_array(41719);
		when "1010001011111000" => data_out <= rom_array(41720);
		when "1010001011111001" => data_out <= rom_array(41721);
		when "1010001011111010" => data_out <= rom_array(41722);
		when "1010001011111011" => data_out <= rom_array(41723);
		when "1010001011111100" => data_out <= rom_array(41724);
		when "1010001011111101" => data_out <= rom_array(41725);
		when "1010001011111110" => data_out <= rom_array(41726);
		when "1010001011111111" => data_out <= rom_array(41727);
		when "1010001100000000" => data_out <= rom_array(41728);
		when "1010001100000001" => data_out <= rom_array(41729);
		when "1010001100000010" => data_out <= rom_array(41730);
		when "1010001100000011" => data_out <= rom_array(41731);
		when "1010001100000100" => data_out <= rom_array(41732);
		when "1010001100000101" => data_out <= rom_array(41733);
		when "1010001100000110" => data_out <= rom_array(41734);
		when "1010001100000111" => data_out <= rom_array(41735);
		when "1010001100001000" => data_out <= rom_array(41736);
		when "1010001100001001" => data_out <= rom_array(41737);
		when "1010001100001010" => data_out <= rom_array(41738);
		when "1010001100001011" => data_out <= rom_array(41739);
		when "1010001100001100" => data_out <= rom_array(41740);
		when "1010001100001101" => data_out <= rom_array(41741);
		when "1010001100001110" => data_out <= rom_array(41742);
		when "1010001100001111" => data_out <= rom_array(41743);
		when "1010001100010000" => data_out <= rom_array(41744);
		when "1010001100010001" => data_out <= rom_array(41745);
		when "1010001100010010" => data_out <= rom_array(41746);
		when "1010001100010011" => data_out <= rom_array(41747);
		when "1010001100010100" => data_out <= rom_array(41748);
		when "1010001100010101" => data_out <= rom_array(41749);
		when "1010001100010110" => data_out <= rom_array(41750);
		when "1010001100010111" => data_out <= rom_array(41751);
		when "1010001100011000" => data_out <= rom_array(41752);
		when "1010001100011001" => data_out <= rom_array(41753);
		when "1010001100011010" => data_out <= rom_array(41754);
		when "1010001100011011" => data_out <= rom_array(41755);
		when "1010001100011100" => data_out <= rom_array(41756);
		when "1010001100011101" => data_out <= rom_array(41757);
		when "1010001100011110" => data_out <= rom_array(41758);
		when "1010001100011111" => data_out <= rom_array(41759);
		when "1010001100100000" => data_out <= rom_array(41760);
		when "1010001100100001" => data_out <= rom_array(41761);
		when "1010001100100010" => data_out <= rom_array(41762);
		when "1010001100100011" => data_out <= rom_array(41763);
		when "1010001100100100" => data_out <= rom_array(41764);
		when "1010001100100101" => data_out <= rom_array(41765);
		when "1010001100100110" => data_out <= rom_array(41766);
		when "1010001100100111" => data_out <= rom_array(41767);
		when "1010001100101000" => data_out <= rom_array(41768);
		when "1010001100101001" => data_out <= rom_array(41769);
		when "1010001100101010" => data_out <= rom_array(41770);
		when "1010001100101011" => data_out <= rom_array(41771);
		when "1010001100101100" => data_out <= rom_array(41772);
		when "1010001100101101" => data_out <= rom_array(41773);
		when "1010001100101110" => data_out <= rom_array(41774);
		when "1010001100101111" => data_out <= rom_array(41775);
		when "1010001100110000" => data_out <= rom_array(41776);
		when "1010001100110001" => data_out <= rom_array(41777);
		when "1010001100110010" => data_out <= rom_array(41778);
		when "1010001100110011" => data_out <= rom_array(41779);
		when "1010001100110100" => data_out <= rom_array(41780);
		when "1010001100110101" => data_out <= rom_array(41781);
		when "1010001100110110" => data_out <= rom_array(41782);
		when "1010001100110111" => data_out <= rom_array(41783);
		when "1010001100111000" => data_out <= rom_array(41784);
		when "1010001100111001" => data_out <= rom_array(41785);
		when "1010001100111010" => data_out <= rom_array(41786);
		when "1010001100111011" => data_out <= rom_array(41787);
		when "1010001100111100" => data_out <= rom_array(41788);
		when "1010001100111101" => data_out <= rom_array(41789);
		when "1010001100111110" => data_out <= rom_array(41790);
		when "1010001100111111" => data_out <= rom_array(41791);
		when "1010001101000000" => data_out <= rom_array(41792);
		when "1010001101000001" => data_out <= rom_array(41793);
		when "1010001101000010" => data_out <= rom_array(41794);
		when "1010001101000011" => data_out <= rom_array(41795);
		when "1010001101000100" => data_out <= rom_array(41796);
		when "1010001101000101" => data_out <= rom_array(41797);
		when "1010001101000110" => data_out <= rom_array(41798);
		when "1010001101000111" => data_out <= rom_array(41799);
		when "1010001101001000" => data_out <= rom_array(41800);
		when "1010001101001001" => data_out <= rom_array(41801);
		when "1010001101001010" => data_out <= rom_array(41802);
		when "1010001101001011" => data_out <= rom_array(41803);
		when "1010001101001100" => data_out <= rom_array(41804);
		when "1010001101001101" => data_out <= rom_array(41805);
		when "1010001101001110" => data_out <= rom_array(41806);
		when "1010001101001111" => data_out <= rom_array(41807);
		when "1010001101010000" => data_out <= rom_array(41808);
		when "1010001101010001" => data_out <= rom_array(41809);
		when "1010001101010010" => data_out <= rom_array(41810);
		when "1010001101010011" => data_out <= rom_array(41811);
		when "1010001101010100" => data_out <= rom_array(41812);
		when "1010001101010101" => data_out <= rom_array(41813);
		when "1010001101010110" => data_out <= rom_array(41814);
		when "1010001101010111" => data_out <= rom_array(41815);
		when "1010001101011000" => data_out <= rom_array(41816);
		when "1010001101011001" => data_out <= rom_array(41817);
		when "1010001101011010" => data_out <= rom_array(41818);
		when "1010001101011011" => data_out <= rom_array(41819);
		when "1010001101011100" => data_out <= rom_array(41820);
		when "1010001101011101" => data_out <= rom_array(41821);
		when "1010001101011110" => data_out <= rom_array(41822);
		when "1010001101011111" => data_out <= rom_array(41823);
		when "1010001101100000" => data_out <= rom_array(41824);
		when "1010001101100001" => data_out <= rom_array(41825);
		when "1010001101100010" => data_out <= rom_array(41826);
		when "1010001101100011" => data_out <= rom_array(41827);
		when "1010001101100100" => data_out <= rom_array(41828);
		when "1010001101100101" => data_out <= rom_array(41829);
		when "1010001101100110" => data_out <= rom_array(41830);
		when "1010001101100111" => data_out <= rom_array(41831);
		when "1010001101101000" => data_out <= rom_array(41832);
		when "1010001101101001" => data_out <= rom_array(41833);
		when "1010001101101010" => data_out <= rom_array(41834);
		when "1010001101101011" => data_out <= rom_array(41835);
		when "1010001101101100" => data_out <= rom_array(41836);
		when "1010001101101101" => data_out <= rom_array(41837);
		when "1010001101101110" => data_out <= rom_array(41838);
		when "1010001101101111" => data_out <= rom_array(41839);
		when "1010001101110000" => data_out <= rom_array(41840);
		when "1010001101110001" => data_out <= rom_array(41841);
		when "1010001101110010" => data_out <= rom_array(41842);
		when "1010001101110011" => data_out <= rom_array(41843);
		when "1010001101110100" => data_out <= rom_array(41844);
		when "1010001101110101" => data_out <= rom_array(41845);
		when "1010001101110110" => data_out <= rom_array(41846);
		when "1010001101110111" => data_out <= rom_array(41847);
		when "1010001101111000" => data_out <= rom_array(41848);
		when "1010001101111001" => data_out <= rom_array(41849);
		when "1010001101111010" => data_out <= rom_array(41850);
		when "1010001101111011" => data_out <= rom_array(41851);
		when "1010001101111100" => data_out <= rom_array(41852);
		when "1010001101111101" => data_out <= rom_array(41853);
		when "1010001101111110" => data_out <= rom_array(41854);
		when "1010001101111111" => data_out <= rom_array(41855);
		when "1010001110000000" => data_out <= rom_array(41856);
		when "1010001110000001" => data_out <= rom_array(41857);
		when "1010001110000010" => data_out <= rom_array(41858);
		when "1010001110000011" => data_out <= rom_array(41859);
		when "1010001110000100" => data_out <= rom_array(41860);
		when "1010001110000101" => data_out <= rom_array(41861);
		when "1010001110000110" => data_out <= rom_array(41862);
		when "1010001110000111" => data_out <= rom_array(41863);
		when "1010001110001000" => data_out <= rom_array(41864);
		when "1010001110001001" => data_out <= rom_array(41865);
		when "1010001110001010" => data_out <= rom_array(41866);
		when "1010001110001011" => data_out <= rom_array(41867);
		when "1010001110001100" => data_out <= rom_array(41868);
		when "1010001110001101" => data_out <= rom_array(41869);
		when "1010001110001110" => data_out <= rom_array(41870);
		when "1010001110001111" => data_out <= rom_array(41871);
		when "1010001110010000" => data_out <= rom_array(41872);
		when "1010001110010001" => data_out <= rom_array(41873);
		when "1010001110010010" => data_out <= rom_array(41874);
		when "1010001110010011" => data_out <= rom_array(41875);
		when "1010001110010100" => data_out <= rom_array(41876);
		when "1010001110010101" => data_out <= rom_array(41877);
		when "1010001110010110" => data_out <= rom_array(41878);
		when "1010001110010111" => data_out <= rom_array(41879);
		when "1010001110011000" => data_out <= rom_array(41880);
		when "1010001110011001" => data_out <= rom_array(41881);
		when "1010001110011010" => data_out <= rom_array(41882);
		when "1010001110011011" => data_out <= rom_array(41883);
		when "1010001110011100" => data_out <= rom_array(41884);
		when "1010001110011101" => data_out <= rom_array(41885);
		when "1010001110011110" => data_out <= rom_array(41886);
		when "1010001110011111" => data_out <= rom_array(41887);
		when "1010001110100000" => data_out <= rom_array(41888);
		when "1010001110100001" => data_out <= rom_array(41889);
		when "1010001110100010" => data_out <= rom_array(41890);
		when "1010001110100011" => data_out <= rom_array(41891);
		when "1010001110100100" => data_out <= rom_array(41892);
		when "1010001110100101" => data_out <= rom_array(41893);
		when "1010001110100110" => data_out <= rom_array(41894);
		when "1010001110100111" => data_out <= rom_array(41895);
		when "1010001110101000" => data_out <= rom_array(41896);
		when "1010001110101001" => data_out <= rom_array(41897);
		when "1010001110101010" => data_out <= rom_array(41898);
		when "1010001110101011" => data_out <= rom_array(41899);
		when "1010001110101100" => data_out <= rom_array(41900);
		when "1010001110101101" => data_out <= rom_array(41901);
		when "1010001110101110" => data_out <= rom_array(41902);
		when "1010001110101111" => data_out <= rom_array(41903);
		when "1010001110110000" => data_out <= rom_array(41904);
		when "1010001110110001" => data_out <= rom_array(41905);
		when "1010001110110010" => data_out <= rom_array(41906);
		when "1010001110110011" => data_out <= rom_array(41907);
		when "1010001110110100" => data_out <= rom_array(41908);
		when "1010001110110101" => data_out <= rom_array(41909);
		when "1010001110110110" => data_out <= rom_array(41910);
		when "1010001110110111" => data_out <= rom_array(41911);
		when "1010001110111000" => data_out <= rom_array(41912);
		when "1010001110111001" => data_out <= rom_array(41913);
		when "1010001110111010" => data_out <= rom_array(41914);
		when "1010001110111011" => data_out <= rom_array(41915);
		when "1010001110111100" => data_out <= rom_array(41916);
		when "1010001110111101" => data_out <= rom_array(41917);
		when "1010001110111110" => data_out <= rom_array(41918);
		when "1010001110111111" => data_out <= rom_array(41919);
		when "1010001111000000" => data_out <= rom_array(41920);
		when "1010001111000001" => data_out <= rom_array(41921);
		when "1010001111000010" => data_out <= rom_array(41922);
		when "1010001111000011" => data_out <= rom_array(41923);
		when "1010001111000100" => data_out <= rom_array(41924);
		when "1010001111000101" => data_out <= rom_array(41925);
		when "1010001111000110" => data_out <= rom_array(41926);
		when "1010001111000111" => data_out <= rom_array(41927);
		when "1010001111001000" => data_out <= rom_array(41928);
		when "1010001111001001" => data_out <= rom_array(41929);
		when "1010001111001010" => data_out <= rom_array(41930);
		when "1010001111001011" => data_out <= rom_array(41931);
		when "1010001111001100" => data_out <= rom_array(41932);
		when "1010001111001101" => data_out <= rom_array(41933);
		when "1010001111001110" => data_out <= rom_array(41934);
		when "1010001111001111" => data_out <= rom_array(41935);
		when "1010001111010000" => data_out <= rom_array(41936);
		when "1010001111010001" => data_out <= rom_array(41937);
		when "1010001111010010" => data_out <= rom_array(41938);
		when "1010001111010011" => data_out <= rom_array(41939);
		when "1010001111010100" => data_out <= rom_array(41940);
		when "1010001111010101" => data_out <= rom_array(41941);
		when "1010001111010110" => data_out <= rom_array(41942);
		when "1010001111010111" => data_out <= rom_array(41943);
		when "1010001111011000" => data_out <= rom_array(41944);
		when "1010001111011001" => data_out <= rom_array(41945);
		when "1010001111011010" => data_out <= rom_array(41946);
		when "1010001111011011" => data_out <= rom_array(41947);
		when "1010001111011100" => data_out <= rom_array(41948);
		when "1010001111011101" => data_out <= rom_array(41949);
		when "1010001111011110" => data_out <= rom_array(41950);
		when "1010001111011111" => data_out <= rom_array(41951);
		when "1010001111100000" => data_out <= rom_array(41952);
		when "1010001111100001" => data_out <= rom_array(41953);
		when "1010001111100010" => data_out <= rom_array(41954);
		when "1010001111100011" => data_out <= rom_array(41955);
		when "1010001111100100" => data_out <= rom_array(41956);
		when "1010001111100101" => data_out <= rom_array(41957);
		when "1010001111100110" => data_out <= rom_array(41958);
		when "1010001111100111" => data_out <= rom_array(41959);
		when "1010001111101000" => data_out <= rom_array(41960);
		when "1010001111101001" => data_out <= rom_array(41961);
		when "1010001111101010" => data_out <= rom_array(41962);
		when "1010001111101011" => data_out <= rom_array(41963);
		when "1010001111101100" => data_out <= rom_array(41964);
		when "1010001111101101" => data_out <= rom_array(41965);
		when "1010001111101110" => data_out <= rom_array(41966);
		when "1010001111101111" => data_out <= rom_array(41967);
		when "1010001111110000" => data_out <= rom_array(41968);
		when "1010001111110001" => data_out <= rom_array(41969);
		when "1010001111110010" => data_out <= rom_array(41970);
		when "1010001111110011" => data_out <= rom_array(41971);
		when "1010001111110100" => data_out <= rom_array(41972);
		when "1010001111110101" => data_out <= rom_array(41973);
		when "1010001111110110" => data_out <= rom_array(41974);
		when "1010001111110111" => data_out <= rom_array(41975);
		when "1010001111111000" => data_out <= rom_array(41976);
		when "1010001111111001" => data_out <= rom_array(41977);
		when "1010001111111010" => data_out <= rom_array(41978);
		when "1010001111111011" => data_out <= rom_array(41979);
		when "1010001111111100" => data_out <= rom_array(41980);
		when "1010001111111101" => data_out <= rom_array(41981);
		when "1010001111111110" => data_out <= rom_array(41982);
		when "1010001111111111" => data_out <= rom_array(41983);
		when "1010010000000000" => data_out <= rom_array(41984);
		when "1010010000000001" => data_out <= rom_array(41985);
		when "1010010000000010" => data_out <= rom_array(41986);
		when "1010010000000011" => data_out <= rom_array(41987);
		when "1010010000000100" => data_out <= rom_array(41988);
		when "1010010000000101" => data_out <= rom_array(41989);
		when "1010010000000110" => data_out <= rom_array(41990);
		when "1010010000000111" => data_out <= rom_array(41991);
		when "1010010000001000" => data_out <= rom_array(41992);
		when "1010010000001001" => data_out <= rom_array(41993);
		when "1010010000001010" => data_out <= rom_array(41994);
		when "1010010000001011" => data_out <= rom_array(41995);
		when "1010010000001100" => data_out <= rom_array(41996);
		when "1010010000001101" => data_out <= rom_array(41997);
		when "1010010000001110" => data_out <= rom_array(41998);
		when "1010010000001111" => data_out <= rom_array(41999);
		when "1010010000010000" => data_out <= rom_array(42000);
		when "1010010000010001" => data_out <= rom_array(42001);
		when "1010010000010010" => data_out <= rom_array(42002);
		when "1010010000010011" => data_out <= rom_array(42003);
		when "1010010000010100" => data_out <= rom_array(42004);
		when "1010010000010101" => data_out <= rom_array(42005);
		when "1010010000010110" => data_out <= rom_array(42006);
		when "1010010000010111" => data_out <= rom_array(42007);
		when "1010010000011000" => data_out <= rom_array(42008);
		when "1010010000011001" => data_out <= rom_array(42009);
		when "1010010000011010" => data_out <= rom_array(42010);
		when "1010010000011011" => data_out <= rom_array(42011);
		when "1010010000011100" => data_out <= rom_array(42012);
		when "1010010000011101" => data_out <= rom_array(42013);
		when "1010010000011110" => data_out <= rom_array(42014);
		when "1010010000011111" => data_out <= rom_array(42015);
		when "1010010000100000" => data_out <= rom_array(42016);
		when "1010010000100001" => data_out <= rom_array(42017);
		when "1010010000100010" => data_out <= rom_array(42018);
		when "1010010000100011" => data_out <= rom_array(42019);
		when "1010010000100100" => data_out <= rom_array(42020);
		when "1010010000100101" => data_out <= rom_array(42021);
		when "1010010000100110" => data_out <= rom_array(42022);
		when "1010010000100111" => data_out <= rom_array(42023);
		when "1010010000101000" => data_out <= rom_array(42024);
		when "1010010000101001" => data_out <= rom_array(42025);
		when "1010010000101010" => data_out <= rom_array(42026);
		when "1010010000101011" => data_out <= rom_array(42027);
		when "1010010000101100" => data_out <= rom_array(42028);
		when "1010010000101101" => data_out <= rom_array(42029);
		when "1010010000101110" => data_out <= rom_array(42030);
		when "1010010000101111" => data_out <= rom_array(42031);
		when "1010010000110000" => data_out <= rom_array(42032);
		when "1010010000110001" => data_out <= rom_array(42033);
		when "1010010000110010" => data_out <= rom_array(42034);
		when "1010010000110011" => data_out <= rom_array(42035);
		when "1010010000110100" => data_out <= rom_array(42036);
		when "1010010000110101" => data_out <= rom_array(42037);
		when "1010010000110110" => data_out <= rom_array(42038);
		when "1010010000110111" => data_out <= rom_array(42039);
		when "1010010000111000" => data_out <= rom_array(42040);
		when "1010010000111001" => data_out <= rom_array(42041);
		when "1010010000111010" => data_out <= rom_array(42042);
		when "1010010000111011" => data_out <= rom_array(42043);
		when "1010010000111100" => data_out <= rom_array(42044);
		when "1010010000111101" => data_out <= rom_array(42045);
		when "1010010000111110" => data_out <= rom_array(42046);
		when "1010010000111111" => data_out <= rom_array(42047);
		when "1010010001000000" => data_out <= rom_array(42048);
		when "1010010001000001" => data_out <= rom_array(42049);
		when "1010010001000010" => data_out <= rom_array(42050);
		when "1010010001000011" => data_out <= rom_array(42051);
		when "1010010001000100" => data_out <= rom_array(42052);
		when "1010010001000101" => data_out <= rom_array(42053);
		when "1010010001000110" => data_out <= rom_array(42054);
		when "1010010001000111" => data_out <= rom_array(42055);
		when "1010010001001000" => data_out <= rom_array(42056);
		when "1010010001001001" => data_out <= rom_array(42057);
		when "1010010001001010" => data_out <= rom_array(42058);
		when "1010010001001011" => data_out <= rom_array(42059);
		when "1010010001001100" => data_out <= rom_array(42060);
		when "1010010001001101" => data_out <= rom_array(42061);
		when "1010010001001110" => data_out <= rom_array(42062);
		when "1010010001001111" => data_out <= rom_array(42063);
		when "1010010001010000" => data_out <= rom_array(42064);
		when "1010010001010001" => data_out <= rom_array(42065);
		when "1010010001010010" => data_out <= rom_array(42066);
		when "1010010001010011" => data_out <= rom_array(42067);
		when "1010010001010100" => data_out <= rom_array(42068);
		when "1010010001010101" => data_out <= rom_array(42069);
		when "1010010001010110" => data_out <= rom_array(42070);
		when "1010010001010111" => data_out <= rom_array(42071);
		when "1010010001011000" => data_out <= rom_array(42072);
		when "1010010001011001" => data_out <= rom_array(42073);
		when "1010010001011010" => data_out <= rom_array(42074);
		when "1010010001011011" => data_out <= rom_array(42075);
		when "1010010001011100" => data_out <= rom_array(42076);
		when "1010010001011101" => data_out <= rom_array(42077);
		when "1010010001011110" => data_out <= rom_array(42078);
		when "1010010001011111" => data_out <= rom_array(42079);
		when "1010010001100000" => data_out <= rom_array(42080);
		when "1010010001100001" => data_out <= rom_array(42081);
		when "1010010001100010" => data_out <= rom_array(42082);
		when "1010010001100011" => data_out <= rom_array(42083);
		when "1010010001100100" => data_out <= rom_array(42084);
		when "1010010001100101" => data_out <= rom_array(42085);
		when "1010010001100110" => data_out <= rom_array(42086);
		when "1010010001100111" => data_out <= rom_array(42087);
		when "1010010001101000" => data_out <= rom_array(42088);
		when "1010010001101001" => data_out <= rom_array(42089);
		when "1010010001101010" => data_out <= rom_array(42090);
		when "1010010001101011" => data_out <= rom_array(42091);
		when "1010010001101100" => data_out <= rom_array(42092);
		when "1010010001101101" => data_out <= rom_array(42093);
		when "1010010001101110" => data_out <= rom_array(42094);
		when "1010010001101111" => data_out <= rom_array(42095);
		when "1010010001110000" => data_out <= rom_array(42096);
		when "1010010001110001" => data_out <= rom_array(42097);
		when "1010010001110010" => data_out <= rom_array(42098);
		when "1010010001110011" => data_out <= rom_array(42099);
		when "1010010001110100" => data_out <= rom_array(42100);
		when "1010010001110101" => data_out <= rom_array(42101);
		when "1010010001110110" => data_out <= rom_array(42102);
		when "1010010001110111" => data_out <= rom_array(42103);
		when "1010010001111000" => data_out <= rom_array(42104);
		when "1010010001111001" => data_out <= rom_array(42105);
		when "1010010001111010" => data_out <= rom_array(42106);
		when "1010010001111011" => data_out <= rom_array(42107);
		when "1010010001111100" => data_out <= rom_array(42108);
		when "1010010001111101" => data_out <= rom_array(42109);
		when "1010010001111110" => data_out <= rom_array(42110);
		when "1010010001111111" => data_out <= rom_array(42111);
		when "1010010010000000" => data_out <= rom_array(42112);
		when "1010010010000001" => data_out <= rom_array(42113);
		when "1010010010000010" => data_out <= rom_array(42114);
		when "1010010010000011" => data_out <= rom_array(42115);
		when "1010010010000100" => data_out <= rom_array(42116);
		when "1010010010000101" => data_out <= rom_array(42117);
		when "1010010010000110" => data_out <= rom_array(42118);
		when "1010010010000111" => data_out <= rom_array(42119);
		when "1010010010001000" => data_out <= rom_array(42120);
		when "1010010010001001" => data_out <= rom_array(42121);
		when "1010010010001010" => data_out <= rom_array(42122);
		when "1010010010001011" => data_out <= rom_array(42123);
		when "1010010010001100" => data_out <= rom_array(42124);
		when "1010010010001101" => data_out <= rom_array(42125);
		when "1010010010001110" => data_out <= rom_array(42126);
		when "1010010010001111" => data_out <= rom_array(42127);
		when "1010010010010000" => data_out <= rom_array(42128);
		when "1010010010010001" => data_out <= rom_array(42129);
		when "1010010010010010" => data_out <= rom_array(42130);
		when "1010010010010011" => data_out <= rom_array(42131);
		when "1010010010010100" => data_out <= rom_array(42132);
		when "1010010010010101" => data_out <= rom_array(42133);
		when "1010010010010110" => data_out <= rom_array(42134);
		when "1010010010010111" => data_out <= rom_array(42135);
		when "1010010010011000" => data_out <= rom_array(42136);
		when "1010010010011001" => data_out <= rom_array(42137);
		when "1010010010011010" => data_out <= rom_array(42138);
		when "1010010010011011" => data_out <= rom_array(42139);
		when "1010010010011100" => data_out <= rom_array(42140);
		when "1010010010011101" => data_out <= rom_array(42141);
		when "1010010010011110" => data_out <= rom_array(42142);
		when "1010010010011111" => data_out <= rom_array(42143);
		when "1010010010100000" => data_out <= rom_array(42144);
		when "1010010010100001" => data_out <= rom_array(42145);
		when "1010010010100010" => data_out <= rom_array(42146);
		when "1010010010100011" => data_out <= rom_array(42147);
		when "1010010010100100" => data_out <= rom_array(42148);
		when "1010010010100101" => data_out <= rom_array(42149);
		when "1010010010100110" => data_out <= rom_array(42150);
		when "1010010010100111" => data_out <= rom_array(42151);
		when "1010010010101000" => data_out <= rom_array(42152);
		when "1010010010101001" => data_out <= rom_array(42153);
		when "1010010010101010" => data_out <= rom_array(42154);
		when "1010010010101011" => data_out <= rom_array(42155);
		when "1010010010101100" => data_out <= rom_array(42156);
		when "1010010010101101" => data_out <= rom_array(42157);
		when "1010010010101110" => data_out <= rom_array(42158);
		when "1010010010101111" => data_out <= rom_array(42159);
		when "1010010010110000" => data_out <= rom_array(42160);
		when "1010010010110001" => data_out <= rom_array(42161);
		when "1010010010110010" => data_out <= rom_array(42162);
		when "1010010010110011" => data_out <= rom_array(42163);
		when "1010010010110100" => data_out <= rom_array(42164);
		when "1010010010110101" => data_out <= rom_array(42165);
		when "1010010010110110" => data_out <= rom_array(42166);
		when "1010010010110111" => data_out <= rom_array(42167);
		when "1010010010111000" => data_out <= rom_array(42168);
		when "1010010010111001" => data_out <= rom_array(42169);
		when "1010010010111010" => data_out <= rom_array(42170);
		when "1010010010111011" => data_out <= rom_array(42171);
		when "1010010010111100" => data_out <= rom_array(42172);
		when "1010010010111101" => data_out <= rom_array(42173);
		when "1010010010111110" => data_out <= rom_array(42174);
		when "1010010010111111" => data_out <= rom_array(42175);
		when "1010010011000000" => data_out <= rom_array(42176);
		when "1010010011000001" => data_out <= rom_array(42177);
		when "1010010011000010" => data_out <= rom_array(42178);
		when "1010010011000011" => data_out <= rom_array(42179);
		when "1010010011000100" => data_out <= rom_array(42180);
		when "1010010011000101" => data_out <= rom_array(42181);
		when "1010010011000110" => data_out <= rom_array(42182);
		when "1010010011000111" => data_out <= rom_array(42183);
		when "1010010011001000" => data_out <= rom_array(42184);
		when "1010010011001001" => data_out <= rom_array(42185);
		when "1010010011001010" => data_out <= rom_array(42186);
		when "1010010011001011" => data_out <= rom_array(42187);
		when "1010010011001100" => data_out <= rom_array(42188);
		when "1010010011001101" => data_out <= rom_array(42189);
		when "1010010011001110" => data_out <= rom_array(42190);
		when "1010010011001111" => data_out <= rom_array(42191);
		when "1010010011010000" => data_out <= rom_array(42192);
		when "1010010011010001" => data_out <= rom_array(42193);
		when "1010010011010010" => data_out <= rom_array(42194);
		when "1010010011010011" => data_out <= rom_array(42195);
		when "1010010011010100" => data_out <= rom_array(42196);
		when "1010010011010101" => data_out <= rom_array(42197);
		when "1010010011010110" => data_out <= rom_array(42198);
		when "1010010011010111" => data_out <= rom_array(42199);
		when "1010010011011000" => data_out <= rom_array(42200);
		when "1010010011011001" => data_out <= rom_array(42201);
		when "1010010011011010" => data_out <= rom_array(42202);
		when "1010010011011011" => data_out <= rom_array(42203);
		when "1010010011011100" => data_out <= rom_array(42204);
		when "1010010011011101" => data_out <= rom_array(42205);
		when "1010010011011110" => data_out <= rom_array(42206);
		when "1010010011011111" => data_out <= rom_array(42207);
		when "1010010011100000" => data_out <= rom_array(42208);
		when "1010010011100001" => data_out <= rom_array(42209);
		when "1010010011100010" => data_out <= rom_array(42210);
		when "1010010011100011" => data_out <= rom_array(42211);
		when "1010010011100100" => data_out <= rom_array(42212);
		when "1010010011100101" => data_out <= rom_array(42213);
		when "1010010011100110" => data_out <= rom_array(42214);
		when "1010010011100111" => data_out <= rom_array(42215);
		when "1010010011101000" => data_out <= rom_array(42216);
		when "1010010011101001" => data_out <= rom_array(42217);
		when "1010010011101010" => data_out <= rom_array(42218);
		when "1010010011101011" => data_out <= rom_array(42219);
		when "1010010011101100" => data_out <= rom_array(42220);
		when "1010010011101101" => data_out <= rom_array(42221);
		when "1010010011101110" => data_out <= rom_array(42222);
		when "1010010011101111" => data_out <= rom_array(42223);
		when "1010010011110000" => data_out <= rom_array(42224);
		when "1010010011110001" => data_out <= rom_array(42225);
		when "1010010011110010" => data_out <= rom_array(42226);
		when "1010010011110011" => data_out <= rom_array(42227);
		when "1010010011110100" => data_out <= rom_array(42228);
		when "1010010011110101" => data_out <= rom_array(42229);
		when "1010010011110110" => data_out <= rom_array(42230);
		when "1010010011110111" => data_out <= rom_array(42231);
		when "1010010011111000" => data_out <= rom_array(42232);
		when "1010010011111001" => data_out <= rom_array(42233);
		when "1010010011111010" => data_out <= rom_array(42234);
		when "1010010011111011" => data_out <= rom_array(42235);
		when "1010010011111100" => data_out <= rom_array(42236);
		when "1010010011111101" => data_out <= rom_array(42237);
		when "1010010011111110" => data_out <= rom_array(42238);
		when "1010010011111111" => data_out <= rom_array(42239);
		when "1010010100000000" => data_out <= rom_array(42240);
		when "1010010100000001" => data_out <= rom_array(42241);
		when "1010010100000010" => data_out <= rom_array(42242);
		when "1010010100000011" => data_out <= rom_array(42243);
		when "1010010100000100" => data_out <= rom_array(42244);
		when "1010010100000101" => data_out <= rom_array(42245);
		when "1010010100000110" => data_out <= rom_array(42246);
		when "1010010100000111" => data_out <= rom_array(42247);
		when "1010010100001000" => data_out <= rom_array(42248);
		when "1010010100001001" => data_out <= rom_array(42249);
		when "1010010100001010" => data_out <= rom_array(42250);
		when "1010010100001011" => data_out <= rom_array(42251);
		when "1010010100001100" => data_out <= rom_array(42252);
		when "1010010100001101" => data_out <= rom_array(42253);
		when "1010010100001110" => data_out <= rom_array(42254);
		when "1010010100001111" => data_out <= rom_array(42255);
		when "1010010100010000" => data_out <= rom_array(42256);
		when "1010010100010001" => data_out <= rom_array(42257);
		when "1010010100010010" => data_out <= rom_array(42258);
		when "1010010100010011" => data_out <= rom_array(42259);
		when "1010010100010100" => data_out <= rom_array(42260);
		when "1010010100010101" => data_out <= rom_array(42261);
		when "1010010100010110" => data_out <= rom_array(42262);
		when "1010010100010111" => data_out <= rom_array(42263);
		when "1010010100011000" => data_out <= rom_array(42264);
		when "1010010100011001" => data_out <= rom_array(42265);
		when "1010010100011010" => data_out <= rom_array(42266);
		when "1010010100011011" => data_out <= rom_array(42267);
		when "1010010100011100" => data_out <= rom_array(42268);
		when "1010010100011101" => data_out <= rom_array(42269);
		when "1010010100011110" => data_out <= rom_array(42270);
		when "1010010100011111" => data_out <= rom_array(42271);
		when "1010010100100000" => data_out <= rom_array(42272);
		when "1010010100100001" => data_out <= rom_array(42273);
		when "1010010100100010" => data_out <= rom_array(42274);
		when "1010010100100011" => data_out <= rom_array(42275);
		when "1010010100100100" => data_out <= rom_array(42276);
		when "1010010100100101" => data_out <= rom_array(42277);
		when "1010010100100110" => data_out <= rom_array(42278);
		when "1010010100100111" => data_out <= rom_array(42279);
		when "1010010100101000" => data_out <= rom_array(42280);
		when "1010010100101001" => data_out <= rom_array(42281);
		when "1010010100101010" => data_out <= rom_array(42282);
		when "1010010100101011" => data_out <= rom_array(42283);
		when "1010010100101100" => data_out <= rom_array(42284);
		when "1010010100101101" => data_out <= rom_array(42285);
		when "1010010100101110" => data_out <= rom_array(42286);
		when "1010010100101111" => data_out <= rom_array(42287);
		when "1010010100110000" => data_out <= rom_array(42288);
		when "1010010100110001" => data_out <= rom_array(42289);
		when "1010010100110010" => data_out <= rom_array(42290);
		when "1010010100110011" => data_out <= rom_array(42291);
		when "1010010100110100" => data_out <= rom_array(42292);
		when "1010010100110101" => data_out <= rom_array(42293);
		when "1010010100110110" => data_out <= rom_array(42294);
		when "1010010100110111" => data_out <= rom_array(42295);
		when "1010010100111000" => data_out <= rom_array(42296);
		when "1010010100111001" => data_out <= rom_array(42297);
		when "1010010100111010" => data_out <= rom_array(42298);
		when "1010010100111011" => data_out <= rom_array(42299);
		when "1010010100111100" => data_out <= rom_array(42300);
		when "1010010100111101" => data_out <= rom_array(42301);
		when "1010010100111110" => data_out <= rom_array(42302);
		when "1010010100111111" => data_out <= rom_array(42303);
		when "1010010101000000" => data_out <= rom_array(42304);
		when "1010010101000001" => data_out <= rom_array(42305);
		when "1010010101000010" => data_out <= rom_array(42306);
		when "1010010101000011" => data_out <= rom_array(42307);
		when "1010010101000100" => data_out <= rom_array(42308);
		when "1010010101000101" => data_out <= rom_array(42309);
		when "1010010101000110" => data_out <= rom_array(42310);
		when "1010010101000111" => data_out <= rom_array(42311);
		when "1010010101001000" => data_out <= rom_array(42312);
		when "1010010101001001" => data_out <= rom_array(42313);
		when "1010010101001010" => data_out <= rom_array(42314);
		when "1010010101001011" => data_out <= rom_array(42315);
		when "1010010101001100" => data_out <= rom_array(42316);
		when "1010010101001101" => data_out <= rom_array(42317);
		when "1010010101001110" => data_out <= rom_array(42318);
		when "1010010101001111" => data_out <= rom_array(42319);
		when "1010010101010000" => data_out <= rom_array(42320);
		when "1010010101010001" => data_out <= rom_array(42321);
		when "1010010101010010" => data_out <= rom_array(42322);
		when "1010010101010011" => data_out <= rom_array(42323);
		when "1010010101010100" => data_out <= rom_array(42324);
		when "1010010101010101" => data_out <= rom_array(42325);
		when "1010010101010110" => data_out <= rom_array(42326);
		when "1010010101010111" => data_out <= rom_array(42327);
		when "1010010101011000" => data_out <= rom_array(42328);
		when "1010010101011001" => data_out <= rom_array(42329);
		when "1010010101011010" => data_out <= rom_array(42330);
		when "1010010101011011" => data_out <= rom_array(42331);
		when "1010010101011100" => data_out <= rom_array(42332);
		when "1010010101011101" => data_out <= rom_array(42333);
		when "1010010101011110" => data_out <= rom_array(42334);
		when "1010010101011111" => data_out <= rom_array(42335);
		when "1010010101100000" => data_out <= rom_array(42336);
		when "1010010101100001" => data_out <= rom_array(42337);
		when "1010010101100010" => data_out <= rom_array(42338);
		when "1010010101100011" => data_out <= rom_array(42339);
		when "1010010101100100" => data_out <= rom_array(42340);
		when "1010010101100101" => data_out <= rom_array(42341);
		when "1010010101100110" => data_out <= rom_array(42342);
		when "1010010101100111" => data_out <= rom_array(42343);
		when "1010010101101000" => data_out <= rom_array(42344);
		when "1010010101101001" => data_out <= rom_array(42345);
		when "1010010101101010" => data_out <= rom_array(42346);
		when "1010010101101011" => data_out <= rom_array(42347);
		when "1010010101101100" => data_out <= rom_array(42348);
		when "1010010101101101" => data_out <= rom_array(42349);
		when "1010010101101110" => data_out <= rom_array(42350);
		when "1010010101101111" => data_out <= rom_array(42351);
		when "1010010101110000" => data_out <= rom_array(42352);
		when "1010010101110001" => data_out <= rom_array(42353);
		when "1010010101110010" => data_out <= rom_array(42354);
		when "1010010101110011" => data_out <= rom_array(42355);
		when "1010010101110100" => data_out <= rom_array(42356);
		when "1010010101110101" => data_out <= rom_array(42357);
		when "1010010101110110" => data_out <= rom_array(42358);
		when "1010010101110111" => data_out <= rom_array(42359);
		when "1010010101111000" => data_out <= rom_array(42360);
		when "1010010101111001" => data_out <= rom_array(42361);
		when "1010010101111010" => data_out <= rom_array(42362);
		when "1010010101111011" => data_out <= rom_array(42363);
		when "1010010101111100" => data_out <= rom_array(42364);
		when "1010010101111101" => data_out <= rom_array(42365);
		when "1010010101111110" => data_out <= rom_array(42366);
		when "1010010101111111" => data_out <= rom_array(42367);
		when "1010010110000000" => data_out <= rom_array(42368);
		when "1010010110000001" => data_out <= rom_array(42369);
		when "1010010110000010" => data_out <= rom_array(42370);
		when "1010010110000011" => data_out <= rom_array(42371);
		when "1010010110000100" => data_out <= rom_array(42372);
		when "1010010110000101" => data_out <= rom_array(42373);
		when "1010010110000110" => data_out <= rom_array(42374);
		when "1010010110000111" => data_out <= rom_array(42375);
		when "1010010110001000" => data_out <= rom_array(42376);
		when "1010010110001001" => data_out <= rom_array(42377);
		when "1010010110001010" => data_out <= rom_array(42378);
		when "1010010110001011" => data_out <= rom_array(42379);
		when "1010010110001100" => data_out <= rom_array(42380);
		when "1010010110001101" => data_out <= rom_array(42381);
		when "1010010110001110" => data_out <= rom_array(42382);
		when "1010010110001111" => data_out <= rom_array(42383);
		when "1010010110010000" => data_out <= rom_array(42384);
		when "1010010110010001" => data_out <= rom_array(42385);
		when "1010010110010010" => data_out <= rom_array(42386);
		when "1010010110010011" => data_out <= rom_array(42387);
		when "1010010110010100" => data_out <= rom_array(42388);
		when "1010010110010101" => data_out <= rom_array(42389);
		when "1010010110010110" => data_out <= rom_array(42390);
		when "1010010110010111" => data_out <= rom_array(42391);
		when "1010010110011000" => data_out <= rom_array(42392);
		when "1010010110011001" => data_out <= rom_array(42393);
		when "1010010110011010" => data_out <= rom_array(42394);
		when "1010010110011011" => data_out <= rom_array(42395);
		when "1010010110011100" => data_out <= rom_array(42396);
		when "1010010110011101" => data_out <= rom_array(42397);
		when "1010010110011110" => data_out <= rom_array(42398);
		when "1010010110011111" => data_out <= rom_array(42399);
		when "1010010110100000" => data_out <= rom_array(42400);
		when "1010010110100001" => data_out <= rom_array(42401);
		when "1010010110100010" => data_out <= rom_array(42402);
		when "1010010110100011" => data_out <= rom_array(42403);
		when "1010010110100100" => data_out <= rom_array(42404);
		when "1010010110100101" => data_out <= rom_array(42405);
		when "1010010110100110" => data_out <= rom_array(42406);
		when "1010010110100111" => data_out <= rom_array(42407);
		when "1010010110101000" => data_out <= rom_array(42408);
		when "1010010110101001" => data_out <= rom_array(42409);
		when "1010010110101010" => data_out <= rom_array(42410);
		when "1010010110101011" => data_out <= rom_array(42411);
		when "1010010110101100" => data_out <= rom_array(42412);
		when "1010010110101101" => data_out <= rom_array(42413);
		when "1010010110101110" => data_out <= rom_array(42414);
		when "1010010110101111" => data_out <= rom_array(42415);
		when "1010010110110000" => data_out <= rom_array(42416);
		when "1010010110110001" => data_out <= rom_array(42417);
		when "1010010110110010" => data_out <= rom_array(42418);
		when "1010010110110011" => data_out <= rom_array(42419);
		when "1010010110110100" => data_out <= rom_array(42420);
		when "1010010110110101" => data_out <= rom_array(42421);
		when "1010010110110110" => data_out <= rom_array(42422);
		when "1010010110110111" => data_out <= rom_array(42423);
		when "1010010110111000" => data_out <= rom_array(42424);
		when "1010010110111001" => data_out <= rom_array(42425);
		when "1010010110111010" => data_out <= rom_array(42426);
		when "1010010110111011" => data_out <= rom_array(42427);
		when "1010010110111100" => data_out <= rom_array(42428);
		when "1010010110111101" => data_out <= rom_array(42429);
		when "1010010110111110" => data_out <= rom_array(42430);
		when "1010010110111111" => data_out <= rom_array(42431);
		when "1010010111000000" => data_out <= rom_array(42432);
		when "1010010111000001" => data_out <= rom_array(42433);
		when "1010010111000010" => data_out <= rom_array(42434);
		when "1010010111000011" => data_out <= rom_array(42435);
		when "1010010111000100" => data_out <= rom_array(42436);
		when "1010010111000101" => data_out <= rom_array(42437);
		when "1010010111000110" => data_out <= rom_array(42438);
		when "1010010111000111" => data_out <= rom_array(42439);
		when "1010010111001000" => data_out <= rom_array(42440);
		when "1010010111001001" => data_out <= rom_array(42441);
		when "1010010111001010" => data_out <= rom_array(42442);
		when "1010010111001011" => data_out <= rom_array(42443);
		when "1010010111001100" => data_out <= rom_array(42444);
		when "1010010111001101" => data_out <= rom_array(42445);
		when "1010010111001110" => data_out <= rom_array(42446);
		when "1010010111001111" => data_out <= rom_array(42447);
		when "1010010111010000" => data_out <= rom_array(42448);
		when "1010010111010001" => data_out <= rom_array(42449);
		when "1010010111010010" => data_out <= rom_array(42450);
		when "1010010111010011" => data_out <= rom_array(42451);
		when "1010010111010100" => data_out <= rom_array(42452);
		when "1010010111010101" => data_out <= rom_array(42453);
		when "1010010111010110" => data_out <= rom_array(42454);
		when "1010010111010111" => data_out <= rom_array(42455);
		when "1010010111011000" => data_out <= rom_array(42456);
		when "1010010111011001" => data_out <= rom_array(42457);
		when "1010010111011010" => data_out <= rom_array(42458);
		when "1010010111011011" => data_out <= rom_array(42459);
		when "1010010111011100" => data_out <= rom_array(42460);
		when "1010010111011101" => data_out <= rom_array(42461);
		when "1010010111011110" => data_out <= rom_array(42462);
		when "1010010111011111" => data_out <= rom_array(42463);
		when "1010010111100000" => data_out <= rom_array(42464);
		when "1010010111100001" => data_out <= rom_array(42465);
		when "1010010111100010" => data_out <= rom_array(42466);
		when "1010010111100011" => data_out <= rom_array(42467);
		when "1010010111100100" => data_out <= rom_array(42468);
		when "1010010111100101" => data_out <= rom_array(42469);
		when "1010010111100110" => data_out <= rom_array(42470);
		when "1010010111100111" => data_out <= rom_array(42471);
		when "1010010111101000" => data_out <= rom_array(42472);
		when "1010010111101001" => data_out <= rom_array(42473);
		when "1010010111101010" => data_out <= rom_array(42474);
		when "1010010111101011" => data_out <= rom_array(42475);
		when "1010010111101100" => data_out <= rom_array(42476);
		when "1010010111101101" => data_out <= rom_array(42477);
		when "1010010111101110" => data_out <= rom_array(42478);
		when "1010010111101111" => data_out <= rom_array(42479);
		when "1010010111110000" => data_out <= rom_array(42480);
		when "1010010111110001" => data_out <= rom_array(42481);
		when "1010010111110010" => data_out <= rom_array(42482);
		when "1010010111110011" => data_out <= rom_array(42483);
		when "1010010111110100" => data_out <= rom_array(42484);
		when "1010010111110101" => data_out <= rom_array(42485);
		when "1010010111110110" => data_out <= rom_array(42486);
		when "1010010111110111" => data_out <= rom_array(42487);
		when "1010010111111000" => data_out <= rom_array(42488);
		when "1010010111111001" => data_out <= rom_array(42489);
		when "1010010111111010" => data_out <= rom_array(42490);
		when "1010010111111011" => data_out <= rom_array(42491);
		when "1010010111111100" => data_out <= rom_array(42492);
		when "1010010111111101" => data_out <= rom_array(42493);
		when "1010010111111110" => data_out <= rom_array(42494);
		when "1010010111111111" => data_out <= rom_array(42495);
		when "1010011000000000" => data_out <= rom_array(42496);
		when "1010011000000001" => data_out <= rom_array(42497);
		when "1010011000000010" => data_out <= rom_array(42498);
		when "1010011000000011" => data_out <= rom_array(42499);
		when "1010011000000100" => data_out <= rom_array(42500);
		when "1010011000000101" => data_out <= rom_array(42501);
		when "1010011000000110" => data_out <= rom_array(42502);
		when "1010011000000111" => data_out <= rom_array(42503);
		when "1010011000001000" => data_out <= rom_array(42504);
		when "1010011000001001" => data_out <= rom_array(42505);
		when "1010011000001010" => data_out <= rom_array(42506);
		when "1010011000001011" => data_out <= rom_array(42507);
		when "1010011000001100" => data_out <= rom_array(42508);
		when "1010011000001101" => data_out <= rom_array(42509);
		when "1010011000001110" => data_out <= rom_array(42510);
		when "1010011000001111" => data_out <= rom_array(42511);
		when "1010011000010000" => data_out <= rom_array(42512);
		when "1010011000010001" => data_out <= rom_array(42513);
		when "1010011000010010" => data_out <= rom_array(42514);
		when "1010011000010011" => data_out <= rom_array(42515);
		when "1010011000010100" => data_out <= rom_array(42516);
		when "1010011000010101" => data_out <= rom_array(42517);
		when "1010011000010110" => data_out <= rom_array(42518);
		when "1010011000010111" => data_out <= rom_array(42519);
		when "1010011000011000" => data_out <= rom_array(42520);
		when "1010011000011001" => data_out <= rom_array(42521);
		when "1010011000011010" => data_out <= rom_array(42522);
		when "1010011000011011" => data_out <= rom_array(42523);
		when "1010011000011100" => data_out <= rom_array(42524);
		when "1010011000011101" => data_out <= rom_array(42525);
		when "1010011000011110" => data_out <= rom_array(42526);
		when "1010011000011111" => data_out <= rom_array(42527);
		when "1010011000100000" => data_out <= rom_array(42528);
		when "1010011000100001" => data_out <= rom_array(42529);
		when "1010011000100010" => data_out <= rom_array(42530);
		when "1010011000100011" => data_out <= rom_array(42531);
		when "1010011000100100" => data_out <= rom_array(42532);
		when "1010011000100101" => data_out <= rom_array(42533);
		when "1010011000100110" => data_out <= rom_array(42534);
		when "1010011000100111" => data_out <= rom_array(42535);
		when "1010011000101000" => data_out <= rom_array(42536);
		when "1010011000101001" => data_out <= rom_array(42537);
		when "1010011000101010" => data_out <= rom_array(42538);
		when "1010011000101011" => data_out <= rom_array(42539);
		when "1010011000101100" => data_out <= rom_array(42540);
		when "1010011000101101" => data_out <= rom_array(42541);
		when "1010011000101110" => data_out <= rom_array(42542);
		when "1010011000101111" => data_out <= rom_array(42543);
		when "1010011000110000" => data_out <= rom_array(42544);
		when "1010011000110001" => data_out <= rom_array(42545);
		when "1010011000110010" => data_out <= rom_array(42546);
		when "1010011000110011" => data_out <= rom_array(42547);
		when "1010011000110100" => data_out <= rom_array(42548);
		when "1010011000110101" => data_out <= rom_array(42549);
		when "1010011000110110" => data_out <= rom_array(42550);
		when "1010011000110111" => data_out <= rom_array(42551);
		when "1010011000111000" => data_out <= rom_array(42552);
		when "1010011000111001" => data_out <= rom_array(42553);
		when "1010011000111010" => data_out <= rom_array(42554);
		when "1010011000111011" => data_out <= rom_array(42555);
		when "1010011000111100" => data_out <= rom_array(42556);
		when "1010011000111101" => data_out <= rom_array(42557);
		when "1010011000111110" => data_out <= rom_array(42558);
		when "1010011000111111" => data_out <= rom_array(42559);
		when "1010011001000000" => data_out <= rom_array(42560);
		when "1010011001000001" => data_out <= rom_array(42561);
		when "1010011001000010" => data_out <= rom_array(42562);
		when "1010011001000011" => data_out <= rom_array(42563);
		when "1010011001000100" => data_out <= rom_array(42564);
		when "1010011001000101" => data_out <= rom_array(42565);
		when "1010011001000110" => data_out <= rom_array(42566);
		when "1010011001000111" => data_out <= rom_array(42567);
		when "1010011001001000" => data_out <= rom_array(42568);
		when "1010011001001001" => data_out <= rom_array(42569);
		when "1010011001001010" => data_out <= rom_array(42570);
		when "1010011001001011" => data_out <= rom_array(42571);
		when "1010011001001100" => data_out <= rom_array(42572);
		when "1010011001001101" => data_out <= rom_array(42573);
		when "1010011001001110" => data_out <= rom_array(42574);
		when "1010011001001111" => data_out <= rom_array(42575);
		when "1010011001010000" => data_out <= rom_array(42576);
		when "1010011001010001" => data_out <= rom_array(42577);
		when "1010011001010010" => data_out <= rom_array(42578);
		when "1010011001010011" => data_out <= rom_array(42579);
		when "1010011001010100" => data_out <= rom_array(42580);
		when "1010011001010101" => data_out <= rom_array(42581);
		when "1010011001010110" => data_out <= rom_array(42582);
		when "1010011001010111" => data_out <= rom_array(42583);
		when "1010011001011000" => data_out <= rom_array(42584);
		when "1010011001011001" => data_out <= rom_array(42585);
		when "1010011001011010" => data_out <= rom_array(42586);
		when "1010011001011011" => data_out <= rom_array(42587);
		when "1010011001011100" => data_out <= rom_array(42588);
		when "1010011001011101" => data_out <= rom_array(42589);
		when "1010011001011110" => data_out <= rom_array(42590);
		when "1010011001011111" => data_out <= rom_array(42591);
		when "1010011001100000" => data_out <= rom_array(42592);
		when "1010011001100001" => data_out <= rom_array(42593);
		when "1010011001100010" => data_out <= rom_array(42594);
		when "1010011001100011" => data_out <= rom_array(42595);
		when "1010011001100100" => data_out <= rom_array(42596);
		when "1010011001100101" => data_out <= rom_array(42597);
		when "1010011001100110" => data_out <= rom_array(42598);
		when "1010011001100111" => data_out <= rom_array(42599);
		when "1010011001101000" => data_out <= rom_array(42600);
		when "1010011001101001" => data_out <= rom_array(42601);
		when "1010011001101010" => data_out <= rom_array(42602);
		when "1010011001101011" => data_out <= rom_array(42603);
		when "1010011001101100" => data_out <= rom_array(42604);
		when "1010011001101101" => data_out <= rom_array(42605);
		when "1010011001101110" => data_out <= rom_array(42606);
		when "1010011001101111" => data_out <= rom_array(42607);
		when "1010011001110000" => data_out <= rom_array(42608);
		when "1010011001110001" => data_out <= rom_array(42609);
		when "1010011001110010" => data_out <= rom_array(42610);
		when "1010011001110011" => data_out <= rom_array(42611);
		when "1010011001110100" => data_out <= rom_array(42612);
		when "1010011001110101" => data_out <= rom_array(42613);
		when "1010011001110110" => data_out <= rom_array(42614);
		when "1010011001110111" => data_out <= rom_array(42615);
		when "1010011001111000" => data_out <= rom_array(42616);
		when "1010011001111001" => data_out <= rom_array(42617);
		when "1010011001111010" => data_out <= rom_array(42618);
		when "1010011001111011" => data_out <= rom_array(42619);
		when "1010011001111100" => data_out <= rom_array(42620);
		when "1010011001111101" => data_out <= rom_array(42621);
		when "1010011001111110" => data_out <= rom_array(42622);
		when "1010011001111111" => data_out <= rom_array(42623);
		when "1010011010000000" => data_out <= rom_array(42624);
		when "1010011010000001" => data_out <= rom_array(42625);
		when "1010011010000010" => data_out <= rom_array(42626);
		when "1010011010000011" => data_out <= rom_array(42627);
		when "1010011010000100" => data_out <= rom_array(42628);
		when "1010011010000101" => data_out <= rom_array(42629);
		when "1010011010000110" => data_out <= rom_array(42630);
		when "1010011010000111" => data_out <= rom_array(42631);
		when "1010011010001000" => data_out <= rom_array(42632);
		when "1010011010001001" => data_out <= rom_array(42633);
		when "1010011010001010" => data_out <= rom_array(42634);
		when "1010011010001011" => data_out <= rom_array(42635);
		when "1010011010001100" => data_out <= rom_array(42636);
		when "1010011010001101" => data_out <= rom_array(42637);
		when "1010011010001110" => data_out <= rom_array(42638);
		when "1010011010001111" => data_out <= rom_array(42639);
		when "1010011010010000" => data_out <= rom_array(42640);
		when "1010011010010001" => data_out <= rom_array(42641);
		when "1010011010010010" => data_out <= rom_array(42642);
		when "1010011010010011" => data_out <= rom_array(42643);
		when "1010011010010100" => data_out <= rom_array(42644);
		when "1010011010010101" => data_out <= rom_array(42645);
		when "1010011010010110" => data_out <= rom_array(42646);
		when "1010011010010111" => data_out <= rom_array(42647);
		when "1010011010011000" => data_out <= rom_array(42648);
		when "1010011010011001" => data_out <= rom_array(42649);
		when "1010011010011010" => data_out <= rom_array(42650);
		when "1010011010011011" => data_out <= rom_array(42651);
		when "1010011010011100" => data_out <= rom_array(42652);
		when "1010011010011101" => data_out <= rom_array(42653);
		when "1010011010011110" => data_out <= rom_array(42654);
		when "1010011010011111" => data_out <= rom_array(42655);
		when "1010011010100000" => data_out <= rom_array(42656);
		when "1010011010100001" => data_out <= rom_array(42657);
		when "1010011010100010" => data_out <= rom_array(42658);
		when "1010011010100011" => data_out <= rom_array(42659);
		when "1010011010100100" => data_out <= rom_array(42660);
		when "1010011010100101" => data_out <= rom_array(42661);
		when "1010011010100110" => data_out <= rom_array(42662);
		when "1010011010100111" => data_out <= rom_array(42663);
		when "1010011010101000" => data_out <= rom_array(42664);
		when "1010011010101001" => data_out <= rom_array(42665);
		when "1010011010101010" => data_out <= rom_array(42666);
		when "1010011010101011" => data_out <= rom_array(42667);
		when "1010011010101100" => data_out <= rom_array(42668);
		when "1010011010101101" => data_out <= rom_array(42669);
		when "1010011010101110" => data_out <= rom_array(42670);
		when "1010011010101111" => data_out <= rom_array(42671);
		when "1010011010110000" => data_out <= rom_array(42672);
		when "1010011010110001" => data_out <= rom_array(42673);
		when "1010011010110010" => data_out <= rom_array(42674);
		when "1010011010110011" => data_out <= rom_array(42675);
		when "1010011010110100" => data_out <= rom_array(42676);
		when "1010011010110101" => data_out <= rom_array(42677);
		when "1010011010110110" => data_out <= rom_array(42678);
		when others => data_out <= (others => '0');
		end case;
	end process;
ClockProc: process (clk, rst) is
begin
if rising_edge(clk) then
	if rst = '1' then
		count <= (others => '0');
	end if;
	if (ENABLE = '1') then
		if (unsigned(count) < rom_type'length) then
			count <= std_logic_vector(unsigned(count) + 1);
		else
			count <= (others => '0');
		end if;
	end if;
end if;
end process;
end Behavioral;