../../../../../basic/pwm/pwm.vhd