../../common/soundgates_pkg.vhd