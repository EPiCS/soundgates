../../../../basic/square/square.vhd