../../../../../basic/cordic/cordic_stage.vhd