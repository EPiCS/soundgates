../../../../basic/cordic/cordic.vhd