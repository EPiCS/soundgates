../../../../../basic/square/square.vhd