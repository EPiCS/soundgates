../../../../../basic/ramp/ramp.vhd