../../basic/triangle/triangle.vhd