../../../../../basic/triangle/triangle.vhd