-- Derived from ..\rechteck.raw
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity SampleDataRom is
Port ( clk    	 : in  STD_LOGIC;
	  	enable 	 : in STD_LOGIC;
	  	data_out : out std_logic_vector( 24 - 1 downto 0);
		rst    	 : in std_logic );
end SampleDataRom;
architecture Behavioral of SampleDataRom is
	type rom_type is array (0 to 4408) of std_logic_vector(24 - 1 downto 0);
constant rom_array : rom_type := 
( 0 => "011111111111111111111111",
1 => "011111111111111111111111",
2 => "011111111111111111111111",
3 => "011111111111111111111111",
4 => "011111111111111111111111",
5 => "011111111111111111111111",
6 => "011111111111111111111111",
7 => "011111111111111111111111",
8 => "011111111111111111111111",
9 => "011111111111111111111111",
10 => "011111111111111111111110",
11 => "011111111111111111111111",
12 => "011111111111111111111111",
13 => "011111111111111111111111",
14 => "011111111111111111111111",
15 => "011111111111111111111110",
16 => "011111111111111111111111",
17 => "011111111111111111111111",
18 => "011111111111111111111110",
19 => "011111111111111111111110",
20 => "011111111111111111111111",
21 => "011111111111111111111111",
22 => "011111111111111111111111",
23 => "011111111111111111111110",
24 => "011111111111111111111111",
25 => "011111111111111111111111",
26 => "011111111111111111111111",
27 => "011111111111111111111100",
28 => "011111111111111111111110",
29 => "011111111111111111111111",
30 => "011111111111111111111111",
31 => "011111111111111111111100",
32 => "011111111111111111111110",
33 => "011111111111111111111111",
34 => "011111111111111111111111",
35 => "011111111111111111111100",
36 => "011111111111111111111110",
37 => "011111111111111111111111",
38 => "011111111111111111111111",
39 => "011111111111111111111110",
40 => "011111111111111111111111",
41 => "011111111111111111111111",
42 => "011111111111111111111111",
43 => "011111111111111111111111",
44 => "011111111111111111111111",
45 => "011111111111111111111110",
46 => "011111111111111111111111",
47 => "011111111111111111111111",
48 => "011111111111111111111111",
49 => "011111111111111111111110",
50 => "011111111111111111111111",
51 => "011111111111111111111111",
52 => "011111111111111111111110",
53 => "011111111111111111111100",
54 => "011111111111111111111111",
55 => "011111111111111111111111",
56 => "011111111111111111111100",
57 => "011111111111111111111111",
58 => "011111111111111111111111",
59 => "011111111111111111111110",
60 => "011111111111111111111110",
61 => "011111111111111111111111",
62 => "011111111111111111111111",
63 => "011111111111111111111100",
64 => "011111111111111111111111",
65 => "011111111111111111111111",
66 => "011111111111111111111111",
67 => "011111111111111111111110",
68 => "011111111111111111111110",
69 => "011111111111111111111111",
70 => "011111111111111111111111",
71 => "011111111111111111111110",
72 => "011111111111111111111100",
73 => "011111111111111111111111",
74 => "011111111111111111111111",
75 => "011111111111111111111110",
76 => "011111111111111111111110",
77 => "011111111111111111111111",
78 => "011111111111111111111111",
79 => "011111111111111111111110",
80 => "011111111111111111111111",
81 => "011111111111111111111111",
82 => "011111111111111111111111",
83 => "011111111111111111111111",
84 => "011111111111111111111111",
85 => "011111111111111111111110",
86 => "011111111111111111111111",
87 => "011111111111111111111111",
88 => "011111111111111111111111",
89 => "011111111111111111111100",
90 => "011111111111111111111111",
91 => "011111111111111111111111",
92 => "011111111111111111111110",
93 => "011111111111111111111110",
94 => "011111111111111111111111",
95 => "011111111111111111111111",
96 => "011111111111111111111111",
97 => "011111111111111111111111",
98 => "011111111111111111111110",
99 => "011111111111111111111111",
100 => "011111111111111111111111",
101 => "100000000000000000000011",
102 => "100000000000000000000000",
103 => "100000000000000000000000",
104 => "100000000000000000000011",
105 => "100000000000000000000010",
106 => "100000000000000000000000",
107 => "100000000000000000000000",
108 => "100000000000000000000000",
109 => "100000000000000000000000",
110 => "100000000000000000000010",
111 => "100000000000000000000010",
112 => "100000000000000000000000",
113 => "100000000000000000000000",
114 => "100000000000000000000100",
115 => "100000000000000000000001",
116 => "100000000000000000000000",
117 => "100000000000000000000000",
118 => "100000000000000000000100",
119 => "100000000000000000000000",
120 => "100000000000000000000000",
121 => "100000000000000000000010",
122 => "100000000000000000000010",
123 => "100000000000000000000000",
124 => "100000000000000000000000",
125 => "100000000000000000000010",
126 => "100000000000000000000000",
127 => "100000000000000000000000",
128 => "100000000000000000000010",
129 => "100000000000000000000001",
130 => "100000000000000000000000",
131 => "100000000000000000000000",
132 => "100000000000000000000010",
133 => "100000000000000000000000",
134 => "100000000000000000000000",
135 => "100000000000000000000000",
136 => "100000000000000000000010",
137 => "100000000000000000000000",
138 => "100000000000000000000000",
139 => "100000000000000000000000",
140 => "100000000000000000000011",
141 => "100000000000000000000010",
142 => "100000000000000000000000",
143 => "100000000000000000000000",
144 => "100000000000000000000010",
145 => "100000000000000000000010",
146 => "100000000000000000000000",
147 => "100000000000000000000000",
148 => "100000000000000000000010",
149 => "100000000000000000000000",
150 => "100000000000000000000000",
151 => "100000000000000000000000",
152 => "100000000000000000000011",
153 => "100000000000000000000001",
154 => "100000000000000000000000",
155 => "100000000000000000000000",
156 => "100000000000000000000010",
157 => "100000000000000000000010",
158 => "100000000000000000000000",
159 => "100000000000000000000000",
160 => "100000000000000000000000",
161 => "100000000000000000000100",
162 => "100000000000000000000000",
163 => "100000000000000000000000",
164 => "100000000000000000000000",
165 => "100000000000000000000100",
166 => "100000000000000000000000",
167 => "100000000000000000000000",
168 => "100000000000000000000000",
169 => "100000000000000000000010",
170 => "100000000000000000000001",
171 => "100000000000000000000000",
172 => "100000000000000000000000",
173 => "100000000000000000000010",
174 => "100000000000000000000010",
175 => "100000000000000000000000",
176 => "100000000000000000000000",
177 => "100000000000000000000100",
178 => "100000000000000000000001",
179 => "100000000000000000000000",
180 => "100000000000000000000000",
181 => "100000000000000000000010",
182 => "100000000000000000000000",
183 => "100000000000000000000000",
184 => "100000000000000000000000",
185 => "100000000000000000000000",
186 => "100000000000000000000010",
187 => "100000000000000000000000",
188 => "100000000000000000000000",
189 => "100000000000000000000000",
190 => "100000000000000000000101",
191 => "100000000000000000000010",
192 => "100000000000000000000000",
193 => "100000000000000000000000",
194 => "100000000000000000000100",
195 => "100000000000000000000010",
196 => "100000000000000000000000",
197 => "100000000000000000000000",
198 => "100000000000000000000011",
199 => "100000000000000000000000",
200 => "100000000000000000000000",
201 => "011111111111111111111111",
202 => "011111111111111111111111",
203 => "011111111111111111111110",
204 => "011111111111111111111110",
205 => "011111111111111111111111",
206 => "011111111111111111111111",
207 => "011111111111111111111111",
208 => "011111111111111111111111",
209 => "011111111111111111111111",
210 => "011111111111111111111101",
211 => "011111111111111111111110",
212 => "011111111111111111111111",
213 => "011111111111111111111111",
214 => "011111111111111111111110",
215 => "011111111111111111111110",
216 => "011111111111111111111111",
217 => "011111111111111111111111",
218 => "011111111111111111111111",
219 => "011111111111111111111100",
220 => "011111111111111111111111",
221 => "011111111111111111111111",
222 => "011111111111111111111111",
223 => "011111111111111111111100",
224 => "011111111111111111111111",
225 => "011111111111111111111111",
226 => "011111111111111111111111",
227 => "011111111111111111111110",
228 => "011111111111111111111111",
229 => "011111111111111111111111",
230 => "011111111111111111111111",
231 => "011111111111111111111110",
232 => "011111111111111111111111",
233 => "011111111111111111111111",
234 => "011111111111111111111111",
235 => "011111111111111111111110",
236 => "011111111111111111111111",
237 => "011111111111111111111111",
238 => "011111111111111111111110",
239 => "011111111111111111111111",
240 => "011111111111111111111111",
241 => "011111111111111111111110",
242 => "011111111111111111111110",
243 => "011111111111111111111111",
244 => "011111111111111111111111",
245 => "011111111111111111111100",
246 => "011111111111111111111111",
247 => "011111111111111111111111",
248 => "011111111111111111111111",
249 => "011111111111111111111100",
250 => "011111111111111111111111",
251 => "011111111111111111111111",
252 => "011111111111111111111111",
253 => "011111111111111111111100",
254 => "011111111111111111111111",
255 => "011111111111111111111111",
256 => "011111111111111111111111",
257 => "011111111111111111111110",
258 => "011111111111111111111110",
259 => "011111111111111111111111",
260 => "011111111111111111111111",
261 => "011111111111111111111111",
262 => "011111111111111111111111",
263 => "011111111111111111111101",
264 => "011111111111111111111111",
265 => "011111111111111111111111",
266 => "011111111111111111111111",
267 => "011111111111111111111101",
268 => "011111111111111111111111",
269 => "011111111111111111111111",
270 => "011111111111111111111111",
271 => "011111111111111111111110",
272 => "011111111111111111111111",
273 => "011111111111111111111111",
274 => "011111111111111111111110",
275 => "011111111111111111111111",
276 => "011111111111111111111111",
277 => "011111111111111111111111",
278 => "011111111111111111111111",
279 => "011111111111111111111111",
280 => "011111111111111111111111",
281 => "011111111111111111111111",
282 => "011111111111111111111110",
283 => "011111111111111111111111",
284 => "011111111111111111111111",
285 => "011111111111111111111111",
286 => "011111111111111111111110",
287 => "011111111111111111111111",
288 => "011111111111111111111111",
289 => "011111111111111111111110",
290 => "011111111111111111111111",
291 => "011111111111111111111111",
292 => "011111111111111111111110",
293 => "011111111111111111111111",
294 => "011111111111111111111111",
295 => "011111111111111111111111",
296 => "011111111111111111111111",
297 => "011111111111111111111111",
298 => "011111111111111111111110",
299 => "011111111111111111111111",
300 => "011111111111111111111111",
301 => "100000000000000000000000",
302 => "100000000000000000000000",
303 => "100000000000000000000001",
304 => "100000000000000000000011",
305 => "100000000000000000000000",
306 => "100000000000000000000000",
307 => "100000000000000000000000",
308 => "100000000000000000000000",
309 => "100000000000000000000010",
310 => "100000000000000000000000",
311 => "100000000000000000000000",
312 => "100000000000000000000000",
313 => "100000000000000000000011",
314 => "100000000000000000000010",
315 => "100000000000000000000000",
316 => "100000000000000000000000",
317 => "100000000000000000000010",
318 => "100000000000000000000101",
319 => "100000000000000000000000",
320 => "100000000000000000000000",
321 => "100000000000000000000010",
322 => "100000000000000000000100",
323 => "100000000000000000000000",
324 => "100000000000000000000000",
325 => "100000000000000000000011",
326 => "100000000000000000000000",
327 => "100000000000000000000000",
328 => "100000000000000000000001",
329 => "100000000000000000000010",
330 => "100000000000000000000000",
331 => "100000000000000000000000",
332 => "100000000000000000000000",
333 => "100000000000000000000010",
334 => "100000000000000000000001",
335 => "100000000000000000000000",
336 => "100000000000000000000000",
337 => "100000000000000000000100",
338 => "100000000000000000000010",
339 => "100000000000000000000000",
340 => "100000000000000000000000",
341 => "100000000000000000000100",
342 => "100000000000000000000001",
343 => "100000000000000000000000",
344 => "100000000000000000000000",
345 => "100000000000000000000001",
346 => "100000000000000000000100",
347 => "100000000000000000000000",
348 => "100000000000000000000000",
349 => "100000000000000000000000",
350 => "100000000000000000000101",
351 => "100000000000000000000000",
352 => "100000000000000000000000",
353 => "100000000000000000000010",
354 => "100000000000000000000010",
355 => "100000000000000000000000",
356 => "100000000000000000000000",
357 => "100000000000000000000010",
358 => "100000000000000000000000",
359 => "100000000000000000000000",
360 => "100000000000000000000000",
361 => "100000000000000000000000",
362 => "100000000000000000000000",
363 => "100000000000000000000010",
364 => "100000000000000000000000",
365 => "100000000000000000000000",
366 => "100000000000000000000000",
367 => "100000000000000000000000",
368 => "100000000000000000000000",
369 => "100000000000000000000010",
370 => "100000000000000000000000",
371 => "100000000000000000000000",
372 => "100000000000000000000000",
373 => "100000000000000000000000",
374 => "100000000000000000000000",
375 => "100000000000000000000001",
376 => "100000000000000000000000",
377 => "100000000000000000000000",
378 => "100000000000000000000001",
379 => "100000000000000000000100",
380 => "100000000000000000000000",
381 => "100000000000000000000000",
382 => "100000000000000000000010",
383 => "100000000000000000000011",
384 => "100000000000000000000000",
385 => "100000000000000000000000",
386 => "100000000000000000000010",
387 => "100000000000000000000010",
388 => "100000000000000000000000",
389 => "100000000000000000000000",
390 => "100000000000000000000010",
391 => "100000000000000000000010",
392 => "100000000000000000000000",
393 => "100000000000000000000000",
394 => "100000000000000000000010",
395 => "100000000000000000000010",
396 => "100000000000000000000000",
397 => "100000000000000000000000",
398 => "100000000000000000000000",
399 => "100000000000000000000000",
400 => "100000000000000000000100",
401 => "011111111111111111111111",
402 => "011111111111111111111100",
403 => "011111111111111111111100",
404 => "011111111111111111111111",
405 => "011111111111111111111111",
406 => "011111111111111111111111",
407 => "011111111111111111111111",
408 => "011111111111111111111110",
409 => "011111111111111111111111",
410 => "011111111111111111111111",
411 => "011111111111111111111111",
412 => "011111111111111111111101",
413 => "011111111111111111111111",
414 => "011111111111111111111111",
415 => "011111111111111111111111",
416 => "011111111111111111111110",
417 => "011111111111111111111111",
418 => "011111111111111111111111",
419 => "011111111111111111111110",
420 => "011111111111111111111111",
421 => "011111111111111111111111",
422 => "011111111111111111111111",
423 => "011111111111111111111100",
424 => "011111111111111111111111",
425 => "011111111111111111111111",
426 => "011111111111111111111111",
427 => "011111111111111111111010",
428 => "011111111111111111111111",
429 => "011111111111111111111111",
430 => "011111111111111111111111",
431 => "011111111111111111111100",
432 => "011111111111111111111111",
433 => "011111111111111111111111",
434 => "011111111111111111111111",
435 => "011111111111111111111101",
436 => "011111111111111111111111",
437 => "011111111111111111111111",
438 => "011111111111111111111110",
439 => "011111111111111111111100",
440 => "011111111111111111111111",
441 => "011111111111111111111111",
442 => "011111111111111111111110",
443 => "011111111111111111111100",
444 => "011111111111111111111111",
445 => "011111111111111111111111",
446 => "011111111111111111111110",
447 => "011111111111111111111101",
448 => "011111111111111111111111",
449 => "011111111111111111111111",
450 => "011111111111111111111111",
451 => "011111111111111111111111",
452 => "011111111111111111111110",
453 => "011111111111111111111111",
454 => "011111111111111111111111",
455 => "011111111111111111111111",
456 => "011111111111111111111101",
457 => "011111111111111111111111",
458 => "011111111111111111111111",
459 => "011111111111111111111111",
460 => "011111111111111111111111",
461 => "011111111111111111111111",
462 => "011111111111111111111110",
463 => "011111111111111111111111",
464 => "011111111111111111111111",
465 => "011111111111111111111111",
466 => "011111111111111111111110",
467 => "011111111111111111111111",
468 => "011111111111111111111111",
469 => "011111111111111111111111",
470 => "011111111111111111111101",
471 => "011111111111111111111110",
472 => "011111111111111111111111",
473 => "011111111111111111111111",
474 => "011111111111111111111110",
475 => "011111111111111111111110",
476 => "011111111111111111111111",
477 => "011111111111111111111111",
478 => "011111111111111111111110",
479 => "011111111111111111111111",
480 => "011111111111111111111111",
481 => "011111111111111111111111",
482 => "011111111111111111111010",
483 => "011111111111111111111111",
484 => "011111111111111111111111",
485 => "011111111111111111111110",
486 => "011111111111111111111100",
487 => "011111111111111111111111",
488 => "011111111111111111111111",
489 => "011111111111111111111111",
490 => "011111111111111111111111",
491 => "011111111111111111111111",
492 => "011111111111111111111110",
493 => "011111111111111111111111",
494 => "011111111111111111111111",
495 => "011111111111111111111111",
496 => "011111111111111111111110",
497 => "011111111111111111111111",
498 => "011111111111111111111111",
499 => "011111111111111111111111",
500 => "011111111111111111111100",
501 => "100000000000000000000001",
502 => "100000000000000000000101",
503 => "100000000000000000000000",
504 => "100000000000000000000000",
505 => "100000000000000000000000",
506 => "100000000000000000000011",
507 => "100000000000000000000010",
508 => "100000000000000000000000",
509 => "100000000000000000000000",
510 => "100000000000000000000000",
511 => "100000000000000000000001",
512 => "100000000000000000000100",
513 => "100000000000000000000000",
514 => "100000000000000000000000",
515 => "100000000000000000000000",
516 => "100000000000000000000100",
517 => "100000000000000000000001",
518 => "100000000000000000000000",
519 => "100000000000000000000000",
520 => "100000000000000000000000",
521 => "100000000000000000000000",
522 => "100000000000000000000011",
523 => "100000000000000000000000",
524 => "100000000000000000000000",
525 => "100000000000000000000000",
526 => "100000000000000000000110",
527 => "100000000000000000000000",
528 => "100000000000000000000000",
529 => "100000000000000000000010",
530 => "100000000000000000000100",
531 => "100000000000000000000000",
532 => "100000000000000000000000",
533 => "100000000000000000000010",
534 => "100000000000000000000010",
535 => "100000000000000000000000",
536 => "100000000000000000000000",
537 => "100000000000000000000000",
538 => "100000000000000000000010",
539 => "100000000000000000000010",
540 => "100000000000000000000000",
541 => "100000000000000000000000",
542 => "100000000000000000000100",
543 => "100000000000000000000000",
544 => "100000000000000000000000",
545 => "100000000000000000000010",
546 => "100000000000000000000100",
547 => "100000000000000000000000",
548 => "100000000000000000000000",
549 => "100000000000000000000110",
550 => "100000000000000000000000",
551 => "100000000000000000000000",
552 => "100000000000000000000100",
553 => "100000000000000000000100",
554 => "100000000000000000000000",
555 => "100000000000000000000000",
556 => "100000000000000000000110",
557 => "100000000000000000000000",
558 => "100000000000000000000000",
559 => "100000000000000000000010",
560 => "100000000000000000000010",
561 => "100000000000000000000000",
562 => "100000000000000000000000",
563 => "100000000000000000000001",
564 => "100000000000000000000000",
565 => "100000000000000000000000",
566 => "100000000000000000000010",
567 => "100000000000000000000000",
568 => "100000000000000000000000",
569 => "100000000000000000000000",
570 => "100000000000000000000001",
571 => "100000000000000000000000",
572 => "100000000000000000000000",
573 => "100000000000000000000000",
574 => "100000000000000000000000",
575 => "100000000000000000000000",
576 => "100000000000000000000000",
577 => "100000000000000000000010",
578 => "100000000000000000000000",
579 => "100000000000000000000000",
580 => "100000000000000000000000",
581 => "100000000000000000000011",
582 => "100000000000000000000001",
583 => "100000000000000000000000",
584 => "100000000000000000000000",
585 => "100000000000000000000100",
586 => "100000000000000000000000",
587 => "100000000000000000000000",
588 => "100000000000000000000010",
589 => "100000000000000000000010",
590 => "100000000000000000000000",
591 => "100000000000000000000000",
592 => "100000000000000000000001",
593 => "100000000000000000000001",
594 => "100000000000000000000000",
595 => "100000000000000000000000",
596 => "100000000000000000000000",
597 => "100000000000000000000000",
598 => "100000000000000000000000",
599 => "100000000000000000000010",
600 => "100000000000000000000000",
601 => "011111111111111111111101",
602 => "011111111111111111111111",
603 => "011111111111111111111111",
604 => "011111111111111111111111",
605 => "011111111111111111111110",
606 => "011111111111111111111111",
607 => "011111111111111111111111",
608 => "011111111111111111111111",
609 => "011111111111111111111111",
610 => "011111111111111111111111",
611 => "011111111111111111111111",
612 => "011111111111111111111111",
613 => "011111111111111111111111",
614 => "011111111111111111111111",
615 => "011111111111111111111111",
616 => "011111111111111111111111",
617 => "011111111111111111111110",
618 => "011111111111111111111111",
619 => "011111111111111111111111",
620 => "011111111111111111111111",
621 => "011111111111111111111110",
622 => "011111111111111111111111",
623 => "011111111111111111111111",
624 => "011111111111111111111111",
625 => "011111111111111111111111",
626 => "011111111111111111111111",
627 => "011111111111111111111110",
628 => "011111111111111111111100",
629 => "011111111111111111111111",
630 => "011111111111111111111111",
631 => "011111111111111111111110",
632 => "011111111111111111111100",
633 => "011111111111111111111111",
634 => "011111111111111111111111",
635 => "011111111111111111111111",
636 => "011111111111111111111110",
637 => "011111111111111111111111",
638 => "011111111111111111111111",
639 => "011111111111111111111111",
640 => "011111111111111111111110",
641 => "011111111111111111111111",
642 => "011111111111111111111111",
643 => "011111111111111111111101",
644 => "011111111111111111111110",
645 => "011111111111111111111111",
646 => "011111111111111111111111",
647 => "011111111111111111111110",
648 => "011111111111111111111110",
649 => "011111111111111111111111",
650 => "011111111111111111111111",
651 => "011111111111111111111111",
652 => "011111111111111111111110",
653 => "011111111111111111111111",
654 => "011111111111111111111111",
655 => "011111111111111111111111",
656 => "011111111111111111111111",
657 => "011111111111111111111111",
658 => "011111111111111111111111",
659 => "011111111111111111111110",
660 => "011111111111111111111110",
661 => "011111111111111111111111",
662 => "011111111111111111111111",
663 => "011111111111111111111111",
664 => "011111111111111111111110",
665 => "011111111111111111111111",
666 => "011111111111111111111111",
667 => "011111111111111111111111",
668 => "011111111111111111111111",
669 => "011111111111111111111110",
670 => "011111111111111111111111",
671 => "011111111111111111111111",
672 => "011111111111111111111111",
673 => "011111111111111111111111",
674 => "011111111111111111111111",
675 => "011111111111111111111111",
676 => "011111111111111111111111",
677 => "011111111111111111111111",
678 => "011111111111111111111111",
679 => "011111111111111111111111",
680 => "011111111111111111111111",
681 => "011111111111111111111111",
682 => "011111111111111111111111",
683 => "011111111111111111111111",
684 => "011111111111111111111111",
685 => "011111111111111111111111",
686 => "011111111111111111111111",
687 => "011111111111111111111111",
688 => "011111111111111111111111",
689 => "011111111111111111111110",
690 => "011111111111111111111111",
691 => "011111111111111111111111",
692 => "011111111111111111111110",
693 => "011111111111111111111110",
694 => "011111111111111111111111",
695 => "011111111111111111111111",
696 => "011111111111111111111100",
697 => "011111111111111111111111",
698 => "011111111111111111111111",
699 => "011111111111111111111111",
700 => "011111111111111111111100",
701 => "100000000000000000000000",
702 => "100000000000000000000010",
703 => "100000000000000000000001",
704 => "100000000000000000000000",
705 => "100000000000000000000000",
706 => "100000000000000000000000",
707 => "100000000000000000000001",
708 => "100000000000000000000000",
709 => "100000000000000000000000",
710 => "100000000000000000000000",
711 => "100000000000000000000000",
712 => "100000000000000000000000",
713 => "100000000000000000000000",
714 => "100000000000000000000000",
715 => "100000000000000000000000",
716 => "100000000000000000000010",
717 => "100000000000000000000000",
718 => "100000000000000000000000",
719 => "100000000000000000000000",
720 => "100000000000000000000010",
721 => "100000000000000000000010",
722 => "100000000000000000000000",
723 => "100000000000000000000000",
724 => "100000000000000000000000",
725 => "100000000000000000000010",
726 => "100000000000000000000001",
727 => "100000000000000000000000",
728 => "100000000000000000000000",
729 => "100000000000000000000000",
730 => "100000000000000000000010",
731 => "100000000000000000000000",
732 => "100000000000000000000000",
733 => "100000000000000000000000",
734 => "100000000000000000000100",
735 => "100000000000000000000010",
736 => "100000000000000000000000",
737 => "100000000000000000000000",
738 => "100000000000000000000100",
739 => "100000000000000000000010",
740 => "100000000000000000000000",
741 => "100000000000000000000000",
742 => "100000000000000000000010",
743 => "100000000000000000000000",
744 => "100000000000000000000000",
745 => "100000000000000000000010",
746 => "100000000000000000000000",
747 => "100000000000000000000000",
748 => "100000000000000000000010",
749 => "100000000000000000000000",
750 => "100000000000000000000000",
751 => "100000000000000000000000",
752 => "100000000000000000000011",
753 => "100000000000000000000000",
754 => "100000000000000000000000",
755 => "100000000000000000000001",
756 => "100000000000000000000100",
757 => "100000000000000000000000",
758 => "100000000000000000000000",
759 => "100000000000000000000001",
760 => "100000000000000000000100",
761 => "100000000000000000000000",
762 => "100000000000000000000000",
763 => "100000000000000000000010",
764 => "100000000000000000000010",
765 => "100000000000000000000000",
766 => "100000000000000000000000",
767 => "100000000000000000000010",
768 => "100000000000000000000010",
769 => "100000000000000000000000",
770 => "100000000000000000000000",
771 => "100000000000000000000001",
772 => "100000000000000000000001",
773 => "100000000000000000000000",
774 => "100000000000000000000000",
775 => "100000000000000000000001",
776 => "100000000000000000000000",
777 => "100000000000000000000000",
778 => "100000000000000000000000",
779 => "100000000000000000000010",
780 => "100000000000000000000010",
781 => "100000000000000000000000",
782 => "100000000000000000000000",
783 => "100000000000000000000001",
784 => "100000000000000000000000",
785 => "100000000000000000000000",
786 => "100000000000000000000010",
787 => "100000000000000000000001",
788 => "100000000000000000000000",
789 => "100000000000000000000000",
790 => "100000000000000000000010",
791 => "100000000000000000000010",
792 => "100000000000000000000000",
793 => "100000000000000000000000",
794 => "100000000000000000000000",
795 => "100000000000000000000001",
796 => "100000000000000000000001",
797 => "100000000000000000000000",
798 => "100000000000000000000000",
799 => "100000000000000000000000",
800 => "100000000000000000000000",
801 => "011111111111111111111111",
802 => "011111111111111111111111",
803 => "011111111111111111111111",
804 => "011111111111111111111011",
805 => "011111111111111111111111",
806 => "011111111111111111111111",
807 => "011111111111111111111111",
808 => "011111111111111111111101",
809 => "011111111111111111111111",
810 => "011111111111111111111111",
811 => "011111111111111111111111",
812 => "011111111111111111111111",
813 => "011111111111111111111111",
814 => "011111111111111111111111",
815 => "011111111111111111111111",
816 => "011111111111111111111111",
817 => "011111111111111111111111",
818 => "011111111111111111111111",
819 => "011111111111111111111111",
820 => "011111111111111111111111",
821 => "011111111111111111111111",
822 => "011111111111111111111111",
823 => "011111111111111111111111",
824 => "011111111111111111111111",
825 => "011111111111111111111111",
826 => "011111111111111111111111",
827 => "011111111111111111111111",
828 => "011111111111111111111111",
829 => "011111111111111111111111",
830 => "011111111111111111111111",
831 => "011111111111111111111111",
832 => "011111111111111111111111",
833 => "011111111111111111111111",
834 => "011111111111111111111111",
835 => "011111111111111111111111",
836 => "011111111111111111111111",
837 => "011111111111111111111110",
838 => "011111111111111111111111",
839 => "011111111111111111111111",
840 => "011111111111111111111111",
841 => "011111111111111111111100",
842 => "011111111111111111111111",
843 => "011111111111111111111111",
844 => "011111111111111111111111",
845 => "011111111111111111111110",
846 => "011111111111111111111111",
847 => "011111111111111111111111",
848 => "011111111111111111111111",
849 => "011111111111111111111111",
850 => "011111111111111111111111",
851 => "011111111111111111111110",
852 => "011111111111111111111111",
853 => "011111111111111111111111",
854 => "011111111111111111111111",
855 => "011111111111111111111111",
856 => "011111111111111111111111",
857 => "011111111111111111111111",
858 => "011111111111111111111111",
859 => "011111111111111111111111",
860 => "011111111111111111111111",
861 => "011111111111111111111110",
862 => "011111111111111111111111",
863 => "011111111111111111111111",
864 => "011111111111111111111111",
865 => "011111111111111111111100",
866 => "011111111111111111111111",
867 => "011111111111111111111111",
868 => "011111111111111111111111",
869 => "011111111111111111111100",
870 => "011111111111111111111111",
871 => "011111111111111111111111",
872 => "011111111111111111111111",
873 => "011111111111111111111110",
874 => "011111111111111111111111",
875 => "011111111111111111111111",
876 => "011111111111111111111111",
877 => "011111111111111111111111",
878 => "011111111111111111111111",
879 => "011111111111111111111111",
880 => "011111111111111111111111",
881 => "011111111111111111111110",
882 => "011111111111111111111111",
883 => "011111111111111111111111",
884 => "011111111111111111111111",
885 => "011111111111111111111110",
886 => "011111111111111111111111",
887 => "011111111111111111111111",
888 => "011111111111111111111111",
889 => "011111111111111111111111",
890 => "011111111111111111111111",
891 => "011111111111111111111111",
892 => "011111111111111111111111",
893 => "011111111111111111111111",
894 => "011111111111111111111111",
895 => "011111111111111111111111",
896 => "011111111111111111111111",
897 => "011111111111111111111111",
898 => "011111111111111111111111",
899 => "011111111111111111111111",
900 => "011111111111111111111111",
901 => "011111111111111111111111",
902 => "011111111111111111111110",
903 => "100000000000000000000000",
904 => "100000000000000000000010",
905 => "100000000000000000000000",
906 => "100000000000000000000000",
907 => "100000000000000000000000",
908 => "100000000000000000000010",
909 => "100000000000000000000000",
910 => "100000000000000000000000",
911 => "100000000000000000000000",
912 => "100000000000000000000000",
913 => "100000000000000000000000",
914 => "100000000000000000000000",
915 => "100000000000000000000000",
916 => "100000000000000000000001",
917 => "100000000000000000000000",
918 => "100000000000000000000000",
919 => "100000000000000000000010",
920 => "100000000000000000000001",
921 => "100000000000000000000000",
922 => "100000000000000000000000",
923 => "100000000000000000000010",
924 => "100000000000000000000000",
925 => "100000000000000000000000",
926 => "100000000000000000000010",
927 => "100000000000000000000001",
928 => "100000000000000000000000",
929 => "100000000000000000000000",
930 => "100000000000000000000010",
931 => "100000000000000000000001",
932 => "100000000000000000000000",
933 => "100000000000000000000000",
934 => "100000000000000000000001",
935 => "100000000000000000000000",
936 => "100000000000000000000000",
937 => "100000000000000000000000",
938 => "100000000000000000000010",
939 => "100000000000000000000001",
940 => "100000000000000000000000",
941 => "100000000000000000000000",
942 => "100000000000000000000010",
943 => "100000000000000000000010",
944 => "100000000000000000000000",
945 => "100000000000000000000000",
946 => "100000000000000000000010",
947 => "100000000000000000000010",
948 => "100000000000000000000000",
949 => "100000000000000000000000",
950 => "100000000000000000000100",
951 => "100000000000000000000010",
952 => "100000000000000000000000",
953 => "100000000000000000000000",
954 => "100000000000000000000110",
955 => "100000000000000000000010",
956 => "100000000000000000000000",
957 => "100000000000000000000000",
958 => "100000000000000000000101",
959 => "100000000000000000000000",
960 => "100000000000000000000000",
961 => "100000000000000000000011",
962 => "100000000000000000000010",
963 => "100000000000000000000000",
964 => "100000000000000000000000",
965 => "100000000000000000000011",
966 => "100000000000000000000000",
967 => "100000000000000000000000",
968 => "100000000000000000000001",
969 => "100000000000000000000001",
970 => "100000000000000000000000",
971 => "100000000000000000000000",
972 => "100000000000000000000010",
973 => "100000000000000000000000",
974 => "100000000000000000000000",
975 => "100000000000000000000001",
976 => "100000000000000000000010",
977 => "100000000000000000000000",
978 => "100000000000000000000000",
979 => "100000000000000000000010",
980 => "100000000000000000000010",
981 => "100000000000000000000000",
982 => "100000000000000000000000",
983 => "100000000000000000000000",
984 => "100000000000000000000010",
985 => "100000000000000000000000",
986 => "100000000000000000000000",
987 => "100000000000000000000000",
988 => "100000000000000000000010",
989 => "100000000000000000000000",
990 => "100000000000000000000000",
991 => "100000000000000000000000",
992 => "100000000000000000000010",
993 => "100000000000000000000001",
994 => "100000000000000000000000",
995 => "100000000000000000000000",
996 => "100000000000000000000011",
997 => "100000000000000000000010",
998 => "100000000000000000000000",
999 => "100000000000000000000000",
1000 => "100000000000000000000100",
1001 => "100000000000000000000000",
1002 => "100000000000000000000000",
1003 => "011111111111111111111111",
1004 => "011111111111111111111111",
1005 => "011111111111111111111101",
1006 => "011111111111111111111110",
1007 => "011111111111111111111111",
1008 => "011111111111111111111111",
1009 => "011111111111111111111111",
1010 => "011111111111111111111111",
1011 => "011111111111111111111111",
1012 => "011111111111111111111101",
1013 => "011111111111111111111111",
1014 => "011111111111111111111111",
1015 => "011111111111111111111110",
1016 => "011111111111111111111101",
1017 => "011111111111111111111111",
1018 => "011111111111111111111111",
1019 => "011111111111111111111110",
1020 => "011111111111111111111110",
1021 => "011111111111111111111111",
1022 => "011111111111111111111111",
1023 => "011111111111111111111111",
1024 => "011111111111111111111110",
1025 => "011111111111111111111111",
1026 => "011111111111111111111111",
1027 => "011111111111111111111111",
1028 => "011111111111111111111101",
1029 => "011111111111111111111101",
1030 => "011111111111111111111111",
1031 => "011111111111111111111111",
1032 => "011111111111111111111100",
1033 => "011111111111111111111100",
1034 => "011111111111111111111111",
1035 => "011111111111111111111111",
1036 => "011111111111111111111110",
1037 => "011111111111111111111110",
1038 => "011111111111111111111111",
1039 => "011111111111111111111111",
1040 => "011111111111111111111111",
1041 => "011111111111111111111110",
1042 => "011111111111111111111110",
1043 => "011111111111111111111111",
1044 => "011111111111111111111111",
1045 => "011111111111111111111101",
1046 => "011111111111111111111110",
1047 => "011111111111111111111111",
1048 => "011111111111111111111111",
1049 => "011111111111111111111110",
1050 => "011111111111111111111111",
1051 => "011111111111111111111111",
1052 => "011111111111111111111111",
1053 => "011111111111111111111111",
1054 => "011111111111111111111111",
1055 => "011111111111111111111111",
1056 => "011111111111111111111111",
1057 => "011111111111111111111111",
1058 => "011111111111111111111111",
1059 => "011111111111111111111111",
1060 => "011111111111111111111111",
1061 => "011111111111111111111111",
1062 => "011111111111111111111111",
1063 => "011111111111111111111111",
1064 => "011111111111111111111111",
1065 => "011111111111111111111111",
1066 => "011111111111111111111111",
1067 => "011111111111111111111111",
1068 => "011111111111111111111111",
1069 => "011111111111111111111111",
1070 => "011111111111111111111111",
1071 => "011111111111111111111111",
1072 => "011111111111111111111111",
1073 => "011111111111111111111110",
1074 => "011111111111111111111110",
1075 => "011111111111111111111111",
1076 => "011111111111111111111111",
1077 => "011111111111111111111111",
1078 => "011111111111111111111110",
1079 => "011111111111111111111111",
1080 => "011111111111111111111111",
1081 => "011111111111111111111111",
1082 => "011111111111111111111111",
1083 => "011111111111111111111111",
1084 => "011111111111111111111111",
1085 => "011111111111111111111110",
1086 => "011111111111111111111111",
1087 => "011111111111111111111111",
1088 => "011111111111111111111111",
1089 => "011111111111111111111110",
1090 => "011111111111111111111110",
1091 => "011111111111111111111111",
1092 => "011111111111111111111111",
1093 => "011111111111111111111111",
1094 => "011111111111111111111110",
1095 => "011111111111111111111101",
1096 => "011111111111111111111111",
1097 => "011111111111111111111111",
1098 => "011111111111111111111110",
1099 => "011111111111111111111110",
1100 => "011111111111111111111111",
1101 => "011111111111111111111111",
1102 => "011111111111111111111110",
1103 => "100000000000000000000000",
1104 => "100000000000000000000010",
1105 => "100000000000000000000000",
1106 => "100000000000000000000000",
1107 => "100000000000000000000000",
1108 => "100000000000000000000000",
1109 => "100000000000000000000000",
1110 => "100000000000000000000000",
1111 => "100000000000000000000000",
1112 => "100000000000000000000001",
1113 => "100000000000000000000000",
1114 => "100000000000000000000000",
1115 => "100000000000000000000001",
1116 => "100000000000000000000100",
1117 => "100000000000000000000000",
1118 => "100000000000000000000000",
1119 => "100000000000000000000010",
1120 => "100000000000000000000000",
1121 => "100000000000000000000000",
1122 => "100000000000000000000001",
1123 => "100000000000000000000000",
1124 => "100000000000000000000000",
1125 => "100000000000000000000001",
1126 => "100000000000000000000000",
1127 => "100000000000000000000000",
1128 => "100000000000000000000100",
1129 => "100000000000000000000000",
1130 => "100000000000000000000000",
1131 => "100000000000000000000001",
1132 => "100000000000000000000010",
1133 => "100000000000000000000000",
1134 => "100000000000000000000000",
1135 => "100000000000000000000000",
1136 => "100000000000000000000000",
1137 => "100000000000000000000001",
1138 => "100000000000000000000000",
1139 => "100000000000000000000000",
1140 => "100000000000000000000010",
1141 => "100000000000000000000101",
1142 => "100000000000000000000000",
1143 => "100000000000000000000000",
1144 => "100000000000000000000011",
1145 => "100000000000000000000100",
1146 => "100000000000000000000000",
1147 => "100000000000000000000000",
1148 => "100000000000000000000000",
1149 => "100000000000000000000001",
1150 => "100000000000000000000100",
1151 => "100000000000000000000000",
1152 => "100000000000000000000000",
1153 => "100000000000000000000000",
1154 => "100000000000000000000110",
1155 => "100000000000000000000000",
1156 => "100000000000000000000000",
1157 => "100000000000000000000000",
1158 => "100000000000000000000011",
1159 => "100000000000000000000000",
1160 => "100000000000000000000000",
1161 => "100000000000000000000000",
1162 => "100000000000000000000000",
1163 => "100000000000000000000000",
1164 => "100000000000000000000010",
1165 => "100000000000000000000001",
1166 => "100000000000000000000000",
1167 => "100000000000000000000000",
1168 => "100000000000000000000011",
1169 => "100000000000000000000010",
1170 => "100000000000000000000000",
1171 => "100000000000000000000000",
1172 => "100000000000000000000011",
1173 => "100000000000000000000010",
1174 => "100000000000000000000000",
1175 => "100000000000000000000000",
1176 => "100000000000000000000011",
1177 => "100000000000000000000010",
1178 => "100000000000000000000000",
1179 => "100000000000000000000000",
1180 => "100000000000000000000010",
1181 => "100000000000000000000010",
1182 => "100000000000000000000000",
1183 => "100000000000000000000000",
1184 => "100000000000000000000000",
1185 => "100000000000000000000010",
1186 => "100000000000000000000000",
1187 => "100000000000000000000000",
1188 => "100000000000000000000000",
1189 => "100000000000000000000000",
1190 => "100000000000000000000000",
1191 => "100000000000000000000001",
1192 => "100000000000000000000000",
1193 => "100000000000000000000000",
1194 => "100000000000000000000000",
1195 => "100000000000000000000010",
1196 => "100000000000000000000000",
1197 => "100000000000000000000000",
1198 => "100000000000000000000000",
1199 => "100000000000000000000100",
1200 => "100000000000000000000000",
1201 => "100000000000000000000000",
1202 => "100000000000000000000000",
1203 => "011111111111111111111111",
1204 => "011111111111111111111111",
1205 => "011111111111111111111100",
1206 => "011111111111111111111111",
1207 => "011111111111111111111111",
1208 => "011111111111111111111110",
1209 => "011111111111111111111110",
1210 => "011111111111111111111111",
1211 => "011111111111111111111111",
1212 => "011111111111111111111111",
1213 => "011111111111111111111111",
1214 => "011111111111111111111111",
1215 => "011111111111111111111110",
1216 => "011111111111111111111111",
1217 => "011111111111111111111111",
1218 => "011111111111111111111111",
1219 => "011111111111111111111110",
1220 => "011111111111111111111111",
1221 => "011111111111111111111111",
1222 => "011111111111111111111111",
1223 => "011111111111111111111110",
1224 => "011111111111111111111111",
1225 => "011111111111111111111111",
1226 => "011111111111111111111110",
1227 => "011111111111111111111111",
1228 => "011111111111111111111111",
1229 => "011111111111111111111111",
1230 => "011111111111111111111110",
1231 => "011111111111111111111111",
1232 => "011111111111111111111111",
1233 => "011111111111111111111110",
1234 => "011111111111111111111101",
1235 => "011111111111111111111111",
1236 => "011111111111111111111111",
1237 => "011111111111111111111110",
1238 => "011111111111111111111011",
1239 => "011111111111111111111111",
1240 => "011111111111111111111111",
1241 => "011111111111111111111110",
1242 => "011111111111111111111110",
1243 => "011111111111111111111111",
1244 => "011111111111111111111111",
1245 => "011111111111111111111110",
1246 => "011111111111111111111111",
1247 => "011111111111111111111111",
1248 => "011111111111111111111111",
1249 => "011111111111111111111111",
1250 => "011111111111111111111100",
1251 => "011111111111111111111110",
1252 => "011111111111111111111111",
1253 => "011111111111111111111111",
1254 => "011111111111111111111011",
1255 => "011111111111111111111110",
1256 => "011111111111111111111111",
1257 => "011111111111111111111111",
1258 => "011111111111111111111110",
1259 => "011111111111111111111110",
1260 => "011111111111111111111111",
1261 => "011111111111111111111111",
1262 => "011111111111111111111111",
1263 => "011111111111111111111111",
1264 => "011111111111111111111110",
1265 => "011111111111111111111111",
1266 => "011111111111111111111111",
1267 => "011111111111111111111111",
1268 => "011111111111111111111111",
1269 => "011111111111111111111111",
1270 => "011111111111111111111110",
1271 => "011111111111111111111111",
1272 => "011111111111111111111111",
1273 => "011111111111111111111110",
1274 => "011111111111111111111111",
1275 => "011111111111111111111111",
1276 => "011111111111111111111111",
1277 => "011111111111111111111111",
1278 => "011111111111111111111111",
1279 => "011111111111111111111111",
1280 => "011111111111111111111111",
1281 => "011111111111111111111111",
1282 => "011111111111111111111110",
1283 => "011111111111111111111110",
1284 => "011111111111111111111111",
1285 => "011111111111111111111111",
1286 => "011111111111111111111101",
1287 => "011111111111111111111111",
1288 => "011111111111111111111111",
1289 => "011111111111111111111110",
1290 => "011111111111111111111111",
1291 => "011111111111111111111111",
1292 => "011111111111111111111101",
1293 => "011111111111111111111111",
1294 => "011111111111111111111111",
1295 => "011111111111111111111111",
1296 => "011111111111111111111110",
1297 => "011111111111111111111111",
1298 => "011111111111111111111111",
1299 => "011111111111111111111100",
1300 => "011111111111111111111110",
1301 => "011111111111111111111111",
1302 => "011111111111111111111111",
1303 => "100000000000000000000000",
1304 => "100000000000000000000000",
1305 => "100000000000000000000010",
1306 => "100000000000000000000110",
1307 => "100000000000000000000000",
1308 => "100000000000000000000000",
1309 => "100000000000000000000000",
1310 => "100000000000000000000010",
1311 => "100000000000000000000000",
1312 => "100000000000000000000000",
1313 => "100000000000000000000010",
1314 => "100000000000000000000000",
1315 => "100000000000000000000000",
1316 => "100000000000000000000000",
1317 => "100000000000000000000000",
1318 => "100000000000000000000010",
1319 => "100000000000000000000010",
1320 => "100000000000000000000000",
1321 => "100000000000000000000000",
1322 => "100000000000000000000011",
1323 => "100000000000000000000100",
1324 => "100000000000000000000000",
1325 => "100000000000000000000000",
1326 => "100000000000000000000010",
1327 => "100000000000000000000010",
1328 => "100000000000000000000000",
1329 => "100000000000000000000000",
1330 => "100000000000000000000010",
1331 => "100000000000000000000001",
1332 => "100000000000000000000000",
1333 => "100000000000000000000001",
1334 => "100000000000000000000010",
1335 => "100000000000000000000000",
1336 => "100000000000000000000000",
1337 => "100000000000000000000000",
1338 => "100000000000000000000000",
1339 => "100000000000000000000000",
1340 => "100000000000000000000000",
1341 => "100000000000000000000000",
1342 => "100000000000000000000001",
1343 => "100000000000000000000010",
1344 => "100000000000000000000000",
1345 => "100000000000000000000000",
1346 => "100000000000000000000010",
1347 => "100000000000000000000001",
1348 => "100000000000000000000000",
1349 => "100000000000000000000000",
1350 => "100000000000000000000000",
1351 => "100000000000000000000000",
1352 => "100000000000000000000010",
1353 => "100000000000000000000100",
1354 => "100000000000000000000000",
1355 => "100000000000000000000000",
1356 => "100000000000000000000010",
1357 => "100000000000000000000010",
1358 => "100000000000000000000000",
1359 => "100000000000000000000000",
1360 => "100000000000000000000000",
1361 => "100000000000000000000000",
1362 => "100000000000000000000001",
1363 => "100000000000000000000010",
1364 => "100000000000000000000000",
1365 => "100000000000000000000000",
1366 => "100000000000000000000011",
1367 => "100000000000000000000000",
1368 => "100000000000000000000000",
1369 => "100000000000000000000000",
1370 => "100000000000000000000100",
1371 => "100000000000000000000000",
1372 => "100000000000000000000000",
1373 => "100000000000000000000000",
1374 => "100000000000000000000011",
1375 => "100000000000000000000000",
1376 => "100000000000000000000000",
1377 => "100000000000000000000000",
1378 => "100000000000000000000010",
1379 => "100000000000000000000000",
1380 => "100000000000000000000000",
1381 => "100000000000000000000000",
1382 => "100000000000000000000000",
1383 => "100000000000000000000010",
1384 => "100000000000000000000001",
1385 => "100000000000000000000000",
1386 => "100000000000000000000000",
1387 => "100000000000000000000100",
1388 => "100000000000000000000010",
1389 => "100000000000000000000000",
1390 => "100000000000000000000000",
1391 => "100000000000000000000010",
1392 => "100000000000000000000010",
1393 => "100000000000000000000000",
1394 => "100000000000000000000000",
1395 => "100000000000000000000010",
1396 => "100000000000000000000010",
1397 => "100000000000000000000000",
1398 => "100000000000000000000000",
1399 => "100000000000000000000010",
1400 => "100000000000000000000010",
1401 => "100000000000000000000000",
1402 => "100000000000000000000000",
1403 => "011111111111111111111111",
1404 => "011111111111111111111111",
1405 => "011111111111111111111111",
1406 => "011111111111111111111110",
1407 => "011111111111111111111110",
1408 => "011111111111111111111111",
1409 => "011111111111111111111111",
1410 => "011111111111111111111111",
1411 => "011111111111111111111110",
1412 => "011111111111111111111111",
1413 => "011111111111111111111111",
1414 => "011111111111111111111111",
1415 => "011111111111111111111101",
1416 => "011111111111111111111111",
1417 => "011111111111111111111111",
1418 => "011111111111111111111111",
1419 => "011111111111111111111101",
1420 => "011111111111111111111111",
1421 => "011111111111111111111111",
1422 => "011111111111111111111111",
1423 => "011111111111111111111111",
1424 => "011111111111111111111111",
1425 => "011111111111111111111111",
1426 => "011111111111111111111111",
1427 => "011111111111111111111111",
1428 => "011111111111111111111111",
1429 => "011111111111111111111111",
1430 => "011111111111111111111111",
1431 => "011111111111111111111111",
1432 => "011111111111111111111111",
1433 => "011111111111111111111111",
1434 => "011111111111111111111111",
1435 => "011111111111111111111111",
1436 => "011111111111111111111110",
1437 => "011111111111111111111111",
1438 => "011111111111111111111111",
1439 => "011111111111111111111110",
1440 => "011111111111111111111110",
1441 => "011111111111111111111111",
1442 => "011111111111111111111111",
1443 => "011111111111111111111110",
1444 => "011111111111111111111111",
1445 => "011111111111111111111111",
1446 => "011111111111111111111110",
1447 => "011111111111111111111111",
1448 => "011111111111111111111111",
1449 => "011111111111111111111111",
1450 => "011111111111111111111100",
1451 => "011111111111111111111111",
1452 => "011111111111111111111111",
1453 => "011111111111111111111110",
1454 => "011111111111111111111100",
1455 => "011111111111111111111111",
1456 => "011111111111111111111111",
1457 => "011111111111111111111100",
1458 => "011111111111111111111110",
1459 => "011111111111111111111111",
1460 => "011111111111111111111111",
1461 => "011111111111111111111110",
1462 => "011111111111111111111111",
1463 => "011111111111111111111111",
1464 => "011111111111111111111111",
1465 => "011111111111111111111111",
1466 => "011111111111111111111111",
1467 => "011111111111111111111101",
1468 => "011111111111111111111110",
1469 => "011111111111111111111111",
1470 => "011111111111111111111111",
1471 => "011111111111111111111111",
1472 => "011111111111111111111101",
1473 => "011111111111111111111111",
1474 => "011111111111111111111111",
1475 => "011111111111111111111111",
1476 => "011111111111111111111110",
1477 => "011111111111111111111111",
1478 => "011111111111111111111111",
1479 => "011111111111111111111110",
1480 => "011111111111111111111111",
1481 => "011111111111111111111111",
1482 => "011111111111111111111111",
1483 => "011111111111111111111110",
1484 => "011111111111111111111111",
1485 => "011111111111111111111111",
1486 => "011111111111111111111111",
1487 => "011111111111111111111111",
1488 => "011111111111111111111111",
1489 => "011111111111111111111110",
1490 => "011111111111111111111111",
1491 => "011111111111111111111111",
1492 => "011111111111111111111111",
1493 => "011111111111111111111100",
1494 => "011111111111111111111111",
1495 => "011111111111111111111111",
1496 => "011111111111111111111111",
1497 => "011111111111111111111100",
1498 => "011111111111111111111111",
1499 => "011111111111111111111111",
1500 => "011111111111111111111111",
1501 => "011111111111111111111110",
1502 => "011111111111111111111111",
1503 => "100000000000000000000001",
1504 => "100000000000000000000001",
1505 => "100000000000000000000000",
1506 => "100000000000000000000000",
1507 => "100000000000000000000000",
1508 => "100000000000000000000001",
1509 => "100000000000000000000010",
1510 => "100000000000000000000000",
1511 => "100000000000000000000000",
1512 => "100000000000000000000000",
1513 => "100000000000000000000100",
1514 => "100000000000000000000010",
1515 => "100000000000000000000000",
1516 => "100000000000000000000000",
1517 => "100000000000000000000100",
1518 => "100000000000000000000100",
1519 => "100000000000000000000000",
1520 => "100000000000000000000000",
1521 => "100000000000000000000110",
1522 => "100000000000000000000011",
1523 => "100000000000000000000000",
1524 => "100000000000000000000000",
1525 => "100000000000000000000110",
1526 => "100000000000000000000001",
1527 => "100000000000000000000000",
1528 => "100000000000000000000001",
1529 => "100000000000000000000100",
1530 => "100000000000000000000000",
1531 => "100000000000000000000000",
1532 => "100000000000000000000010",
1533 => "100000000000000000000100",
1534 => "100000000000000000000000",
1535 => "100000000000000000000000",
1536 => "100000000000000000000010",
1537 => "100000000000000000000001",
1538 => "100000000000000000000000",
1539 => "100000000000000000000000",
1540 => "100000000000000000000010",
1541 => "100000000000000000000000",
1542 => "100000000000000000000000",
1543 => "100000000000000000000000",
1544 => "100000000000000000000010",
1545 => "100000000000000000000010",
1546 => "100000000000000000000000",
1547 => "100000000000000000000000",
1548 => "100000000000000000000001",
1549 => "100000000000000000000000",
1550 => "100000000000000000000000",
1551 => "100000000000000000000010",
1552 => "100000000000000000000000",
1553 => "100000000000000000000000",
1554 => "100000000000000000000001",
1555 => "100000000000000000000100",
1556 => "100000000000000000000000",
1557 => "100000000000000000000000",
1558 => "100000000000000000000010",
1559 => "100000000000000000000000",
1560 => "100000000000000000000000",
1561 => "100000000000000000000010",
1562 => "100000000000000000000010",
1563 => "100000000000000000000000",
1564 => "100000000000000000000000",
1565 => "100000000000000000000001",
1566 => "100000000000000000000000",
1567 => "100000000000000000000000",
1568 => "100000000000000000000001",
1569 => "100000000000000000000000",
1570 => "100000000000000000000000",
1571 => "100000000000000000000000",
1572 => "100000000000000000000000",
1573 => "100000000000000000000000",
1574 => "100000000000000000000010",
1575 => "100000000000000000000010",
1576 => "100000000000000000000000",
1577 => "100000000000000000000000",
1578 => "100000000000000000000010",
1579 => "100000000000000000000010",
1580 => "100000000000000000000000",
1581 => "100000000000000000000000",
1582 => "100000000000000000000000",
1583 => "100000000000000000000000",
1584 => "100000000000000000000001",
1585 => "100000000000000000000010",
1586 => "100000000000000000000000",
1587 => "100000000000000000000000",
1588 => "100000000000000000000010",
1589 => "100000000000000000000010",
1590 => "100000000000000000000000",
1591 => "100000000000000000000000",
1592 => "100000000000000000000000",
1593 => "100000000000000000000010",
1594 => "100000000000000000000010",
1595 => "100000000000000000000000",
1596 => "100000000000000000000000",
1597 => "100000000000000000000001",
1598 => "100000000000000000000100",
1599 => "100000000000000000000000",
1600 => "100000000000000000000000",
1601 => "100000000000000000000000",
1602 => "100000000000000000000010",
1603 => "011111111111111111111111",
1604 => "011111111111111111111111",
1605 => "011111111111111111111110",
1606 => "011111111111111111111111",
1607 => "011111111111111111111111",
1608 => "011111111111111111111110",
1609 => "011111111111111111111100",
1610 => "011111111111111111111111",
1611 => "011111111111111111111111",
1612 => "011111111111111111111110",
1613 => "011111111111111111111110",
1614 => "011111111111111111111111",
1615 => "011111111111111111111111",
1616 => "011111111111111111111111",
1617 => "011111111111111111111111",
1618 => "011111111111111111111110",
1619 => "011111111111111111111110",
1620 => "011111111111111111111111",
1621 => "011111111111111111111111",
1622 => "011111111111111111111110",
1623 => "011111111111111111111110",
1624 => "011111111111111111111111",
1625 => "011111111111111111111111",
1626 => "011111111111111111111111",
1627 => "011111111111111111111110",
1628 => "011111111111111111111101",
1629 => "011111111111111111111111",
1630 => "011111111111111111111111",
1631 => "011111111111111111111111",
1632 => "011111111111111111111110",
1633 => "011111111111111111111110",
1634 => "011111111111111111111111",
1635 => "011111111111111111111111",
1636 => "011111111111111111111111",
1637 => "011111111111111111111101",
1638 => "011111111111111111111111",
1639 => "011111111111111111111111",
1640 => "011111111111111111111111",
1641 => "011111111111111111111101",
1642 => "011111111111111111111111",
1643 => "011111111111111111111111",
1644 => "011111111111111111111111",
1645 => "011111111111111111111111",
1646 => "011111111111111111111111",
1647 => "011111111111111111111111",
1648 => "011111111111111111111111",
1649 => "011111111111111111111110",
1650 => "011111111111111111111111",
1651 => "011111111111111111111111",
1652 => "011111111111111111111111",
1653 => "011111111111111111111111",
1654 => "011111111111111111111111",
1655 => "011111111111111111111111",
1656 => "011111111111111111111111",
1657 => "011111111111111111111111",
1658 => "011111111111111111111111",
1659 => "011111111111111111111111",
1660 => "011111111111111111111111",
1661 => "011111111111111111111110",
1662 => "011111111111111111111111",
1663 => "011111111111111111111111",
1664 => "011111111111111111111111",
1665 => "011111111111111111111110",
1666 => "011111111111111111111111",
1667 => "011111111111111111111111",
1668 => "011111111111111111111111",
1669 => "011111111111111111111111",
1670 => "011111111111111111111111",
1671 => "011111111111111111111111",
1672 => "011111111111111111111111",
1673 => "011111111111111111111111",
1674 => "011111111111111111111111",
1675 => "011111111111111111111111",
1676 => "011111111111111111111111",
1677 => "011111111111111111111111",
1678 => "011111111111111111111110",
1679 => "011111111111111111111111",
1680 => "011111111111111111111111",
1681 => "011111111111111111111111",
1682 => "011111111111111111111110",
1683 => "011111111111111111111111",
1684 => "011111111111111111111111",
1685 => "011111111111111111111111",
1686 => "011111111111111111111111",
1687 => "011111111111111111111111",
1688 => "011111111111111111111111",
1689 => "011111111111111111111011",
1690 => "011111111111111111111111",
1691 => "011111111111111111111111",
1692 => "011111111111111111111111",
1693 => "011111111111111111111100",
1694 => "011111111111111111111111",
1695 => "011111111111111111111111",
1696 => "011111111111111111111111",
1697 => "011111111111111111111111",
1698 => "011111111111111111111111",
1699 => "011111111111111111111111",
1700 => "011111111111111111111111",
1701 => "011111111111111111111111",
1702 => "011111111111111111111111",
1703 => "100000000000000000000000",
1704 => "100000000000000000000000",
1705 => "100000000000000000000010",
1706 => "100000000000000000000001",
1707 => "100000000000000000000001",
1708 => "100000000000000000000000",
1709 => "100000000000000000000000",
1710 => "100000000000000000000010",
1711 => "100000000000000000000011",
1712 => "100000000000000000000000",
1713 => "100000000000000000000000",
1714 => "100000000000000000000000",
1715 => "100000000000000000000000",
1716 => "100000000000000000000000",
1717 => "100000000000000000000010",
1718 => "100000000000000000000000",
1719 => "100000000000000000000000",
1720 => "100000000000000000000000",
1721 => "100000000000000000000010",
1722 => "100000000000000000000000",
1723 => "100000000000000000000000",
1724 => "100000000000000000000001",
1725 => "100000000000000000000010",
1726 => "100000000000000000000000",
1727 => "100000000000000000000000",
1728 => "100000000000000000000010",
1729 => "100000000000000000000000",
1730 => "100000000000000000000000",
1731 => "100000000000000000000010",
1732 => "100000000000000000000000",
1733 => "100000000000000000000000",
1734 => "100000000000000000000000",
1735 => "100000000000000000000010",
1736 => "100000000000000000000000",
1737 => "100000000000000000000000",
1738 => "100000000000000000000000",
1739 => "100000000000000000000001",
1740 => "100000000000000000000010",
1741 => "100000000000000000000000",
1742 => "100000000000000000000000",
1743 => "100000000000000000000000",
1744 => "100000000000000000000010",
1745 => "100000000000000000000000",
1746 => "100000000000000000000000",
1747 => "100000000000000000000010",
1748 => "100000000000000000000001",
1749 => "100000000000000000000000",
1750 => "100000000000000000000000",
1751 => "100000000000000000000100",
1752 => "100000000000000000000000",
1753 => "100000000000000000000000",
1754 => "100000000000000000000000",
1755 => "100000000000000000000011",
1756 => "100000000000000000000000",
1757 => "100000000000000000000000",
1758 => "100000000000000000000001",
1759 => "100000000000000000000011",
1760 => "100000000000000000000000",
1761 => "100000000000000000000000",
1762 => "100000000000000000000000",
1763 => "100000000000000000000010",
1764 => "100000000000000000000100",
1765 => "100000000000000000000000",
1766 => "100000000000000000000000",
1767 => "100000000000000000000010",
1768 => "100000000000000000000011",
1769 => "100000000000000000000000",
1770 => "100000000000000000000000",
1771 => "100000000000000000000100",
1772 => "100000000000000000000000",
1773 => "100000000000000000000000",
1774 => "100000000000000000000010",
1775 => "100000000000000000000100",
1776 => "100000000000000000000000",
1777 => "100000000000000000000000",
1778 => "100000000000000000000001",
1779 => "100000000000000000000010",
1780 => "100000000000000000000000",
1781 => "100000000000000000000000",
1782 => "100000000000000000000010",
1783 => "100000000000000000000001",
1784 => "100000000000000000000000",
1785 => "100000000000000000000000",
1786 => "100000000000000000000010",
1787 => "100000000000000000000000",
1788 => "100000000000000000000000",
1789 => "100000000000000000000010",
1790 => "100000000000000000000010",
1791 => "100000000000000000000000",
1792 => "100000000000000000000000",
1793 => "100000000000000000000011",
1794 => "100000000000000000000011",
1795 => "100000000000000000000000",
1796 => "100000000000000000000000",
1797 => "100000000000000000000010",
1798 => "100000000000000000000001",
1799 => "100000000000000000000000",
1800 => "100000000000000000000000",
1801 => "100000000000000000000010",
1802 => "100000000000000000000000",
1803 => "100000000000000000000000",
1804 => "100000000000000000000010",
1805 => "011111111111111111111111",
1806 => "011111111111111111111111",
1807 => "011111111111111111111110",
1808 => "011111111111111111111111",
1809 => "011111111111111111111111",
1810 => "011111111111111111111111",
1811 => "011111111111111111111110",
1812 => "011111111111111111111111",
1813 => "011111111111111111111111",
1814 => "011111111111111111111111",
1815 => "011111111111111111111111",
1816 => "011111111111111111111111",
1817 => "011111111111111111111110",
1818 => "011111111111111111111111",
1819 => "011111111111111111111111",
1820 => "011111111111111111111111",
1821 => "011111111111111111111100",
1822 => "011111111111111111111111",
1823 => "011111111111111111111111",
1824 => "011111111111111111111111",
1825 => "011111111111111111111101",
1826 => "011111111111111111111111",
1827 => "011111111111111111111111",
1828 => "011111111111111111111101",
1829 => "011111111111111111111110",
1830 => "011111111111111111111111",
1831 => "011111111111111111111111",
1832 => "011111111111111111111101",
1833 => "011111111111111111111110",
1834 => "011111111111111111111111",
1835 => "011111111111111111111111",
1836 => "011111111111111111111110",
1837 => "011111111111111111111101",
1838 => "011111111111111111111111",
1839 => "011111111111111111111111",
1840 => "011111111111111111111110",
1841 => "011111111111111111111111",
1842 => "011111111111111111111111",
1843 => "011111111111111111111110",
1844 => "011111111111111111111010",
1845 => "011111111111111111111111",
1846 => "011111111111111111111111",
1847 => "011111111111111111111101",
1848 => "011111111111111111111010",
1849 => "011111111111111111111111",
1850 => "011111111111111111111111",
1851 => "011111111111111111111110",
1852 => "011111111111111111111100",
1853 => "011111111111111111111111",
1854 => "011111111111111111111111",
1855 => "011111111111111111111110",
1856 => "011111111111111111111110",
1857 => "011111111111111111111111",
1858 => "011111111111111111111111",
1859 => "011111111111111111111110",
1860 => "011111111111111111111101",
1861 => "011111111111111111111111",
1862 => "011111111111111111111111",
1863 => "011111111111111111111110",
1864 => "011111111111111111111111",
1865 => "011111111111111111111111",
1866 => "011111111111111111111111",
1867 => "011111111111111111111111",
1868 => "011111111111111111111111",
1869 => "011111111111111111111111",
1870 => "011111111111111111111111",
1871 => "011111111111111111111111",
1872 => "011111111111111111111111",
1873 => "011111111111111111111110",
1874 => "011111111111111111111111",
1875 => "011111111111111111111111",
1876 => "011111111111111111111111",
1877 => "011111111111111111111110",
1878 => "011111111111111111111111",
1879 => "011111111111111111111111",
1880 => "011111111111111111111110",
1881 => "011111111111111111111111",
1882 => "011111111111111111111111",
1883 => "011111111111111111111111",
1884 => "011111111111111111111111",
1885 => "011111111111111111111111",
1886 => "011111111111111111111111",
1887 => "011111111111111111111111",
1888 => "011111111111111111111111",
1889 => "011111111111111111111111",
1890 => "011111111111111111111111",
1891 => "011111111111111111111111",
1892 => "011111111111111111111111",
1893 => "011111111111111111111111",
1894 => "011111111111111111111111",
1895 => "011111111111111111111111",
1896 => "011111111111111111111111",
1897 => "011111111111111111111111",
1898 => "011111111111111111111111",
1899 => "011111111111111111111111",
1900 => "011111111111111111111111",
1901 => "011111111111111111111110",
1902 => "011111111111111111111111",
1903 => "011111111111111111111111",
1904 => "011111111111111111111110",
1905 => "100000000000000000000000",
1906 => "100000000000000000000010",
1907 => "100000000000000000000000",
1908 => "100000000000000000000000",
1909 => "100000000000000000000001",
1910 => "100000000000000000000000",
1911 => "100000000000000000000000",
1912 => "100000000000000000000010",
1913 => "100000000000000000000010",
1914 => "100000000000000000000000",
1915 => "100000000000000000000000",
1916 => "100000000000000000000011",
1917 => "100000000000000000000010",
1918 => "100000000000000000000000",
1919 => "100000000000000000000000",
1920 => "100000000000000000000010",
1921 => "100000000000000000000000",
1922 => "100000000000000000000000",
1923 => "100000000000000000000001",
1924 => "100000000000000000000000",
1925 => "100000000000000000000000",
1926 => "100000000000000000000010",
1927 => "100000000000000000000001",
1928 => "100000000000000000000000",
1929 => "100000000000000000000000",
1930 => "100000000000000000000011",
1931 => "100000000000000000000000",
1932 => "100000000000000000000000",
1933 => "100000000000000000000000",
1934 => "100000000000000000000000",
1935 => "100000000000000000000000",
1936 => "100000000000000000000010",
1937 => "100000000000000000000010",
1938 => "100000000000000000000000",
1939 => "100000000000000000000000",
1940 => "100000000000000000000010",
1941 => "100000000000000000000100",
1942 => "100000000000000000000000",
1943 => "100000000000000000000000",
1944 => "100000000000000000000001",
1945 => "100000000000000000000110",
1946 => "100000000000000000000000",
1947 => "100000000000000000000000",
1948 => "100000000000000000000000",
1949 => "100000000000000000000110",
1950 => "100000000000000000000010",
1951 => "100000000000000000000000",
1952 => "100000000000000000000000",
1953 => "100000000000000000000100",
1954 => "100000000000000000000101",
1955 => "100000000000000000000000",
1956 => "100000000000000000000000",
1957 => "100000000000000000000001",
1958 => "100000000000000000000110",
1959 => "100000000000000000000000",
1960 => "100000000000000000000000",
1961 => "100000000000000000000000",
1962 => "100000000000000000000100",
1963 => "100000000000000000000000",
1964 => "100000000000000000000000",
1965 => "100000000000000000000000",
1966 => "100000000000000000000010",
1967 => "100000000000000000000000",
1968 => "100000000000000000000000",
1969 => "100000000000000000000000",
1970 => "100000000000000000000000",
1971 => "100000000000000000000010",
1972 => "100000000000000000000000",
1973 => "100000000000000000000000",
1974 => "100000000000000000000000",
1975 => "100000000000000000000000",
1976 => "100000000000000000000000",
1977 => "100000000000000000000001",
1978 => "100000000000000000000001",
1979 => "100000000000000000000000",
1980 => "100000000000000000000000",
1981 => "100000000000000000000010",
1982 => "100000000000000000000011",
1983 => "100000000000000000000000",
1984 => "100000000000000000000000",
1985 => "100000000000000000000010",
1986 => "100000000000000000000010",
1987 => "100000000000000000000000",
1988 => "100000000000000000000000",
1989 => "100000000000000000000100",
1990 => "100000000000000000000000",
1991 => "100000000000000000000000",
1992 => "100000000000000000000010",
1993 => "100000000000000000000110",
1994 => "100000000000000000000000",
1995 => "100000000000000000000000",
1996 => "100000000000000000000001",
1997 => "100000000000000000000100",
1998 => "100000000000000000000000",
1999 => "100000000000000000000000",
2000 => "100000000000000000000000",
2001 => "100000000000000000000000",
2002 => "100000000000000000000000",
2003 => "100000000000000000000010",
2004 => "100000000000000000000000",
2005 => "011111111111111111111101",
2006 => "011111111111111111111111",
2007 => "011111111111111111111111",
2008 => "011111111111111111111111",
2009 => "011111111111111111111111",
2010 => "011111111111111111111111",
2011 => "011111111111111111111111",
2012 => "011111111111111111111111",
2013 => "011111111111111111111111",
2014 => "011111111111111111111111",
2015 => "011111111111111111111111",
2016 => "011111111111111111111111",
2017 => "011111111111111111111110",
2018 => "011111111111111111111111",
2019 => "011111111111111111111111",
2020 => "011111111111111111111111",
2021 => "011111111111111111111101",
2022 => "011111111111111111111111",
2023 => "011111111111111111111111",
2024 => "011111111111111111111110",
2025 => "011111111111111111111110",
2026 => "011111111111111111111111",
2027 => "011111111111111111111111",
2028 => "011111111111111111111100",
2029 => "011111111111111111111110",
2030 => "011111111111111111111111",
2031 => "011111111111111111111111",
2032 => "011111111111111111111101",
2033 => "011111111111111111111110",
2034 => "011111111111111111111111",
2035 => "011111111111111111111111",
2036 => "011111111111111111111111",
2037 => "011111111111111111111111",
2038 => "011111111111111111111110",
2039 => "011111111111111111111111",
2040 => "011111111111111111111111",
2041 => "011111111111111111111110",
2042 => "011111111111111111111111",
2043 => "011111111111111111111111",
2044 => "011111111111111111111111",
2045 => "011111111111111111111111",
2046 => "011111111111111111111111",
2047 => "011111111111111111111111",
2048 => "011111111111111111111111",
2049 => "011111111111111111111110",
2050 => "011111111111111111111111",
2051 => "011111111111111111111111",
2052 => "011111111111111111111111",
2053 => "011111111111111111111101",
2054 => "011111111111111111111111",
2055 => "011111111111111111111111",
2056 => "011111111111111111111111",
2057 => "011111111111111111111111",
2058 => "011111111111111111111101",
2059 => "011111111111111111111110",
2060 => "011111111111111111111111",
2061 => "011111111111111111111111",
2062 => "011111111111111111111100",
2063 => "011111111111111111111101",
2064 => "011111111111111111111111",
2065 => "011111111111111111111111",
2066 => "011111111111111111111111",
2067 => "011111111111111111111110",
2068 => "011111111111111111111111",
2069 => "011111111111111111111111",
2070 => "011111111111111111111111",
2071 => "011111111111111111111110",
2072 => "011111111111111111111111",
2073 => "011111111111111111111111",
2074 => "011111111111111111111111",
2075 => "011111111111111111111110",
2076 => "011111111111111111111111",
2077 => "011111111111111111111111",
2078 => "011111111111111111111111",
2079 => "011111111111111111111111",
2080 => "011111111111111111111111",
2081 => "011111111111111111111111",
2082 => "011111111111111111111111",
2083 => "011111111111111111111111",
2084 => "011111111111111111111111",
2085 => "011111111111111111111111",
2086 => "011111111111111111111111",
2087 => "011111111111111111111100",
2088 => "011111111111111111111111",
2089 => "011111111111111111111111",
2090 => "011111111111111111111110",
2091 => "011111111111111111111111",
2092 => "011111111111111111111111",
2093 => "011111111111111111111111",
2094 => "011111111111111111111100",
2095 => "011111111111111111111111",
2096 => "011111111111111111111111",
2097 => "011111111111111111111110",
2098 => "011111111111111111111010",
2099 => "011111111111111111111111",
2100 => "011111111111111111111111",
2101 => "011111111111111111111101",
2102 => "011111111111111111111110",
2103 => "011111111111111111111111",
2104 => "011111111111111111111111",
2105 => "100000000000000000000000",
2106 => "100000000000000000000000",
2107 => "100000000000000000000100",
2108 => "100000000000000000000000",
2109 => "100000000000000000000000",
2110 => "100000000000000000000000",
2111 => "100000000000000000000100",
2112 => "100000000000000000000001",
2113 => "100000000000000000000000",
2114 => "100000000000000000000000",
2115 => "100000000000000000000010",
2116 => "100000000000000000000000",
2117 => "100000000000000000000000",
2118 => "100000000000000000000000",
2119 => "100000000000000000000000",
2120 => "100000000000000000000000",
2121 => "100000000000000000000001",
2122 => "100000000000000000000000",
2123 => "100000000000000000000000",
2124 => "100000000000000000000000",
2125 => "100000000000000000000000",
2126 => "100000000000000000000000",
2127 => "100000000000000000000010",
2128 => "100000000000000000000011",
2129 => "100000000000000000000000",
2130 => "100000000000000000000000",
2131 => "100000000000000000000000",
2132 => "100000000000000000000010",
2133 => "100000000000000000000000",
2134 => "100000000000000000000000",
2135 => "100000000000000000000000",
2136 => "100000000000000000000010",
2137 => "100000000000000000000010",
2138 => "100000000000000000000000",
2139 => "100000000000000000000000",
2140 => "100000000000000000000010",
2141 => "100000000000000000000010",
2142 => "100000000000000000000000",
2143 => "100000000000000000000000",
2144 => "100000000000000000000010",
2145 => "100000000000000000000001",
2146 => "100000000000000000000000",
2147 => "100000000000000000000001",
2148 => "100000000000000000000001",
2149 => "100000000000000000000000",
2150 => "100000000000000000000000",
2151 => "100000000000000000000010",
2152 => "100000000000000000000001",
2153 => "100000000000000000000000",
2154 => "100000000000000000000000",
2155 => "100000000000000000000001",
2156 => "100000000000000000000010",
2157 => "100000000000000000000000",
2158 => "100000000000000000000000",
2159 => "100000000000000000000000",
2160 => "100000000000000000000001",
2161 => "100000000000000000000000",
2162 => "100000000000000000000001",
2163 => "100000000000000000000000",
2164 => "100000000000000000000000",
2165 => "100000000000000000000000",
2166 => "100000000000000000000010",
2167 => "100000000000000000000000",
2168 => "100000000000000000000000",
2169 => "100000000000000000000000",
2170 => "100000000000000000000000",
2171 => "100000000000000000000000",
2172 => "100000000000000000000010",
2173 => "100000000000000000000001",
2174 => "100000000000000000000000",
2175 => "100000000000000000000000",
2176 => "100000000000000000000010",
2177 => "100000000000000000000000",
2178 => "100000000000000000000000",
2179 => "100000000000000000000000",
2180 => "100000000000000000000010",
2181 => "100000000000000000000000",
2182 => "100000000000000000000000",
2183 => "100000000000000000000001",
2184 => "100000000000000000000000",
2185 => "100000000000000000000000",
2186 => "100000000000000000000100",
2187 => "100000000000000000000000",
2188 => "100000000000000000000000",
2189 => "100000000000000000000000",
2190 => "100000000000000000000010",
2191 => "100000000000000000000000",
2192 => "100000000000000000000000",
2193 => "100000000000000000000000",
2194 => "100000000000000000000000",
2195 => "100000000000000000000000",
2196 => "100000000000000000000000",
2197 => "100000000000000000000000",
2198 => "100000000000000000000010",
2199 => "100000000000000000000010",
2200 => "100000000000000000000000",
2201 => "100000000000000000000000",
2202 => "100000000000000000000010",
2203 => "100000000000000000000010",
2204 => "100000000000000000000000",
2205 => "011111111111111111111110",
2206 => "011111111111111111111110",
2207 => "011111111111111111111111",
2208 => "011111111111111111111111",
2209 => "011111111111111111111111",
2210 => "011111111111111111111111",
2211 => "011111111111111111111111",
2212 => "011111111111111111111110",
2213 => "011111111111111111111110",
2214 => "011111111111111111111111",
2215 => "011111111111111111111111",
2216 => "011111111111111111111110",
2217 => "011111111111111111111111",
2218 => "011111111111111111111111",
2219 => "011111111111111111111111",
2220 => "011111111111111111111111",
2221 => "011111111111111111111111",
2222 => "011111111111111111111111",
2223 => "011111111111111111111111",
2224 => "011111111111111111111111",
2225 => "011111111111111111111100",
2226 => "011111111111111111111111",
2227 => "011111111111111111111111",
2228 => "011111111111111111111111",
2229 => "011111111111111111111100",
2230 => "011111111111111111111110",
2231 => "011111111111111111111111",
2232 => "011111111111111111111111",
2233 => "011111111111111111111111",
2234 => "011111111111111111111011",
2235 => "011111111111111111111111",
2236 => "011111111111111111111111",
2237 => "011111111111111111111111",
2238 => "011111111111111111111100",
2239 => "011111111111111111111111",
2240 => "011111111111111111111111",
2241 => "011111111111111111111110",
2242 => "011111111111111111111111",
2243 => "011111111111111111111111",
2244 => "011111111111111111111111",
2245 => "011111111111111111111110",
2246 => "011111111111111111111110",
2247 => "011111111111111111111111",
2248 => "011111111111111111111111",
2249 => "011111111111111111111110",
2250 => "011111111111111111111101",
2251 => "011111111111111111111111",
2252 => "011111111111111111111111",
2253 => "011111111111111111111111",
2254 => "011111111111111111111110",
2255 => "011111111111111111111111",
2256 => "011111111111111111111111",
2257 => "011111111111111111111111",
2258 => "011111111111111111111111",
2259 => "011111111111111111111111",
2260 => "011111111111111111111111",
2261 => "011111111111111111111111",
2262 => "011111111111111111111110",
2263 => "011111111111111111111111",
2264 => "011111111111111111111111",
2265 => "011111111111111111111111",
2266 => "011111111111111111111100",
2267 => "011111111111111111111111",
2268 => "011111111111111111111111",
2269 => "011111111111111111111111",
2270 => "011111111111111111111111",
2271 => "011111111111111111111111",
2272 => "011111111111111111111111",
2273 => "011111111111111111111111",
2274 => "011111111111111111111111",
2275 => "011111111111111111111110",
2276 => "011111111111111111111110",
2277 => "011111111111111111111111",
2278 => "011111111111111111111111",
2279 => "011111111111111111111100",
2280 => "011111111111111111111110",
2281 => "011111111111111111111111",
2282 => "011111111111111111111111",
2283 => "011111111111111111111110",
2284 => "011111111111111111111110",
2285 => "011111111111111111111111",
2286 => "011111111111111111111111",
2287 => "011111111111111111111111",
2288 => "011111111111111111111111",
2289 => "011111111111111111111110",
2290 => "011111111111111111111111",
2291 => "011111111111111111111111",
2292 => "011111111111111111111111",
2293 => "011111111111111111111111",
2294 => "011111111111111111111111",
2295 => "011111111111111111111110",
2296 => "011111111111111111111111",
2297 => "011111111111111111111111",
2298 => "011111111111111111111111",
2299 => "011111111111111111111110",
2300 => "011111111111111111111111",
2301 => "011111111111111111111111",
2302 => "011111111111111111111110",
2303 => "011111111111111111111110",
2304 => "011111111111111111111111",
2305 => "100000000000000000000010",
2306 => "100000000000000000000000",
2307 => "100000000000000000000000",
2308 => "100000000000000000000010",
2309 => "100000000000000000000010",
2310 => "100000000000000000000000",
2311 => "100000000000000000000000",
2312 => "100000000000000000000000",
2313 => "100000000000000000000100",
2314 => "100000000000000000000000",
2315 => "100000000000000000000000",
2316 => "100000000000000000000000",
2317 => "100000000000000000000011",
2318 => "100000000000000000000000",
2319 => "100000000000000000000000",
2320 => "100000000000000000000010",
2321 => "100000000000000000000000",
2322 => "100000000000000000000000",
2323 => "100000000000000000000010",
2324 => "100000000000000000000010",
2325 => "100000000000000000000000",
2326 => "100000000000000000000000",
2327 => "100000000000000000000011",
2328 => "100000000000000000000010",
2329 => "100000000000000000000000",
2330 => "100000000000000000000000",
2331 => "100000000000000000000100",
2332 => "100000000000000000000010",
2333 => "100000000000000000000000",
2334 => "100000000000000000000000",
2335 => "100000000000000000000010",
2336 => "100000000000000000000010",
2337 => "100000000000000000000000",
2338 => "100000000000000000000000",
2339 => "100000000000000000000001",
2340 => "100000000000000000000010",
2341 => "100000000000000000000000",
2342 => "100000000000000000000000",
2343 => "100000000000000000000000",
2344 => "100000000000000000000010",
2345 => "100000000000000000000010",
2346 => "100000000000000000000000",
2347 => "100000000000000000000000",
2348 => "100000000000000000000011",
2349 => "100000000000000000000010",
2350 => "100000000000000000000000",
2351 => "100000000000000000000000",
2352 => "100000000000000000000001",
2353 => "100000000000000000000000",
2354 => "100000000000000000000001",
2355 => "100000000000000000000100",
2356 => "100000000000000000000000",
2357 => "100000000000000000000000",
2358 => "100000000000000000000010",
2359 => "100000000000000000000100",
2360 => "100000000000000000000000",
2361 => "100000000000000000000000",
2362 => "100000000000000000000010",
2363 => "100000000000000000000010",
2364 => "100000000000000000000000",
2365 => "100000000000000000000000",
2366 => "100000000000000000000010",
2367 => "100000000000000000000001",
2368 => "100000000000000000000000",
2369 => "100000000000000000000000",
2370 => "100000000000000000000001",
2371 => "100000000000000000000001",
2372 => "100000000000000000000000",
2373 => "100000000000000000000000",
2374 => "100000000000000000000000",
2375 => "100000000000000000000000",
2376 => "100000000000000000000000",
2377 => "100000000000000000000000",
2378 => "100000000000000000000000",
2379 => "100000000000000000000000",
2380 => "100000000000000000000010",
2381 => "100000000000000000000000",
2382 => "100000000000000000000000",
2383 => "100000000000000000000000",
2384 => "100000000000000000000100",
2385 => "100000000000000000000010",
2386 => "100000000000000000000000",
2387 => "100000000000000000000000",
2388 => "100000000000000000000011",
2389 => "100000000000000000000010",
2390 => "100000000000000000000000",
2391 => "100000000000000000000000",
2392 => "100000000000000000000000",
2393 => "100000000000000000000010",
2394 => "100000000000000000000010",
2395 => "100000000000000000000000",
2396 => "100000000000000000000000",
2397 => "100000000000000000000100",
2398 => "100000000000000000000000",
2399 => "100000000000000000000000",
2400 => "100000000000000000000010",
2401 => "100000000000000000000000",
2402 => "100000000000000000000000",
2403 => "100000000000000000000010",
2404 => "100000000000000000000100",
2405 => "011111111111111111111101",
2406 => "011111111111111111111100",
2407 => "011111111111111111111111",
2408 => "011111111111111111111111",
2409 => "011111111111111111111111",
2410 => "011111111111111111111110",
2411 => "011111111111111111111111",
2412 => "011111111111111111111111",
2413 => "011111111111111111111111",
2414 => "011111111111111111111111",
2415 => "011111111111111111111111",
2416 => "011111111111111111111111",
2417 => "011111111111111111111111",
2418 => "011111111111111111111111",
2419 => "011111111111111111111111",
2420 => "011111111111111111111111",
2421 => "011111111111111111111111",
2422 => "011111111111111111111100",
2423 => "011111111111111111111111",
2424 => "011111111111111111111111",
2425 => "011111111111111111111110",
2426 => "011111111111111111111100",
2427 => "011111111111111111111111",
2428 => "011111111111111111111111",
2429 => "011111111111111111111110",
2430 => "011111111111111111111111",
2431 => "011111111111111111111111",
2432 => "011111111111111111111111",
2433 => "011111111111111111111111",
2434 => "011111111111111111111111",
2435 => "011111111111111111111110",
2436 => "011111111111111111111110",
2437 => "011111111111111111111111",
2438 => "011111111111111111111111",
2439 => "011111111111111111111110",
2440 => "011111111111111111111100",
2441 => "011111111111111111111111",
2442 => "011111111111111111111111",
2443 => "011111111111111111111111",
2444 => "011111111111111111111101",
2445 => "011111111111111111111111",
2446 => "011111111111111111111111",
2447 => "011111111111111111111111",
2448 => "011111111111111111111111",
2449 => "011111111111111111111111",
2450 => "011111111111111111111100",
2451 => "011111111111111111111110",
2452 => "011111111111111111111111",
2453 => "011111111111111111111111",
2454 => "011111111111111111111010",
2455 => "011111111111111111111111",
2456 => "011111111111111111111111",
2457 => "011111111111111111111111",
2458 => "011111111111111111111100",
2459 => "011111111111111111111111",
2460 => "011111111111111111111111",
2461 => "011111111111111111111110",
2462 => "011111111111111111111110",
2463 => "011111111111111111111111",
2464 => "011111111111111111111111",
2465 => "011111111111111111111110",
2466 => "011111111111111111111111",
2467 => "011111111111111111111111",
2468 => "011111111111111111111110",
2469 => "011111111111111111111101",
2470 => "011111111111111111111111",
2471 => "011111111111111111111111",
2472 => "011111111111111111111110",
2473 => "011111111111111111111100",
2474 => "011111111111111111111111",
2475 => "011111111111111111111111",
2476 => "011111111111111111111111",
2477 => "011111111111111111111111",
2478 => "011111111111111111111110",
2479 => "011111111111111111111110",
2480 => "011111111111111111111111",
2481 => "011111111111111111111111",
2482 => "011111111111111111111110",
2483 => "011111111111111111111111",
2484 => "011111111111111111111111",
2485 => "011111111111111111111101",
2486 => "011111111111111111111111",
2487 => "011111111111111111111111",
2488 => "011111111111111111111101",
2489 => "011111111111111111111100",
2490 => "011111111111111111111111",
2491 => "011111111111111111111111",
2492 => "011111111111111111111100",
2493 => "011111111111111111111110",
2494 => "011111111111111111111111",
2495 => "011111111111111111111111",
2496 => "011111111111111111111111",
2497 => "011111111111111111111111",
2498 => "011111111111111111111111",
2499 => "011111111111111111111111",
2500 => "011111111111111111111111",
2501 => "011111111111111111111111",
2502 => "011111111111111111111110",
2503 => "011111111111111111111111",
2504 => "011111111111111111111111",
2505 => "100000000000000000000000",
2506 => "100000000000000000000000",
2507 => "100000000000000000000000",
2508 => "100000000000000000000000",
2509 => "100000000000000000000000",
2510 => "100000000000000000000010",
2511 => "100000000000000000000000",
2512 => "100000000000000000000000",
2513 => "100000000000000000000000",
2514 => "100000000000000000000100",
2515 => "100000000000000000000010",
2516 => "100000000000000000000000",
2517 => "100000000000000000000000",
2518 => "100000000000000000000011",
2519 => "100000000000000000000011",
2520 => "100000000000000000000000",
2521 => "100000000000000000000000",
2522 => "100000000000000000000001",
2523 => "100000000000000000000010",
2524 => "100000000000000000000000",
2525 => "100000000000000000000000",
2526 => "100000000000000000000001",
2527 => "100000000000000000000000",
2528 => "100000000000000000000000",
2529 => "100000000000000000000000",
2530 => "100000000000000000000010",
2531 => "100000000000000000000000",
2532 => "100000000000000000000000",
2533 => "100000000000000000000000",
2534 => "100000000000000000000001",
2535 => "100000000000000000000000",
2536 => "100000000000000000000000",
2537 => "100000000000000000000000",
2538 => "100000000000000000000011",
2539 => "100000000000000000000010",
2540 => "100000000000000000000000",
2541 => "100000000000000000000000",
2542 => "100000000000000000000000",
2543 => "100000000000000000000010",
2544 => "100000000000000000000000",
2545 => "100000000000000000000000",
2546 => "100000000000000000000000",
2547 => "100000000000000000000000",
2548 => "100000000000000000000001",
2549 => "100000000000000000000010",
2550 => "100000000000000000000000",
2551 => "100000000000000000000000",
2552 => "100000000000000000000001",
2553 => "100000000000000000000010",
2554 => "100000000000000000000000",
2555 => "100000000000000000000000",
2556 => "100000000000000000000010",
2557 => "100000000000000000000010",
2558 => "100000000000000000000000",
2559 => "100000000000000000000000",
2560 => "100000000000000000000000",
2561 => "100000000000000000000001",
2562 => "100000000000000000000010",
2563 => "100000000000000000000000",
2564 => "100000000000000000000000",
2565 => "100000000000000000000000",
2566 => "100000000000000000000100",
2567 => "100000000000000000000000",
2568 => "100000000000000000000000",
2569 => "100000000000000000000000",
2570 => "100000000000000000000011",
2571 => "100000000000000000000000",
2572 => "100000000000000000000000",
2573 => "100000000000000000000000",
2574 => "100000000000000000000010",
2575 => "100000000000000000000000",
2576 => "100000000000000000000000",
2577 => "100000000000000000000010",
2578 => "100000000000000000000000",
2579 => "100000000000000000000000",
2580 => "100000000000000000000000",
2581 => "100000000000000000000010",
2582 => "100000000000000000000000",
2583 => "100000000000000000000000",
2584 => "100000000000000000000000",
2585 => "100000000000000000000000",
2586 => "100000000000000000000010",
2587 => "100000000000000000000001",
2588 => "100000000000000000000000",
2589 => "100000000000000000000000",
2590 => "100000000000000000000011",
2591 => "100000000000000000000001",
2592 => "100000000000000000000000",
2593 => "100000000000000000000000",
2594 => "100000000000000000000010",
2595 => "100000000000000000000000",
2596 => "100000000000000000000000",
2597 => "100000000000000000000000",
2598 => "100000000000000000000000",
2599 => "100000000000000000000001",
2600 => "100000000000000000000000",
2601 => "100000000000000000000000",
2602 => "100000000000000000000000",
2603 => "100000000000000000000000",
2604 => "100000000000000000000000",
2605 => "011111111111111111111111",
2606 => "011111111111111111111111",
2607 => "011111111111111111111111",
2608 => "011111111111111111111110",
2609 => "011111111111111111111111",
2610 => "011111111111111111111111",
2611 => "011111111111111111111111",
2612 => "011111111111111111111110",
2613 => "011111111111111111111111",
2614 => "011111111111111111111111",
2615 => "011111111111111111111100",
2616 => "011111111111111111111111",
2617 => "011111111111111111111111",
2618 => "011111111111111111111111",
2619 => "011111111111111111111010",
2620 => "011111111111111111111100",
2621 => "011111111111111111111111",
2622 => "011111111111111111111111",
2623 => "011111111111111111111111",
2624 => "011111111111111111111100",
2625 => "011111111111111111111111",
2626 => "011111111111111111111111",
2627 => "011111111111111111111111",
2628 => "011111111111111111111110",
2629 => "011111111111111111111111",
2630 => "011111111111111111111111",
2631 => "011111111111111111111101",
2632 => "011111111111111111111111",
2633 => "011111111111111111111111",
2634 => "011111111111111111111110",
2635 => "011111111111111111111110",
2636 => "011111111111111111111111",
2637 => "011111111111111111111111",
2638 => "011111111111111111111111",
2639 => "011111111111111111111110",
2640 => "011111111111111111111110",
2641 => "011111111111111111111111",
2642 => "011111111111111111111111",
2643 => "011111111111111111111101",
2644 => "011111111111111111111100",
2645 => "011111111111111111111111",
2646 => "011111111111111111111111",
2647 => "011111111111111111111111",
2648 => "011111111111111111111111",
2649 => "011111111111111111111111",
2650 => "011111111111111111111111",
2651 => "011111111111111111111111",
2652 => "011111111111111111111111",
2653 => "011111111111111111111111",
2654 => "011111111111111111111111",
2655 => "011111111111111111111111",
2656 => "011111111111111111111110",
2657 => "011111111111111111111111",
2658 => "011111111111111111111111",
2659 => "011111111111111111111110",
2660 => "011111111111111111111100",
2661 => "011111111111111111111111",
2662 => "011111111111111111111111",
2663 => "011111111111111111111111",
2664 => "011111111111111111111110",
2665 => "011111111111111111111110",
2666 => "011111111111111111111111",
2667 => "011111111111111111111111",
2668 => "011111111111111111111111",
2669 => "011111111111111111111101",
2670 => "011111111111111111111111",
2671 => "011111111111111111111111",
2672 => "011111111111111111111111",
2673 => "011111111111111111111110",
2674 => "011111111111111111111111",
2675 => "011111111111111111111111",
2676 => "011111111111111111111111",
2677 => "011111111111111111111111",
2678 => "011111111111111111111111",
2679 => "011111111111111111111110",
2680 => "011111111111111111111111",
2681 => "011111111111111111111111",
2682 => "011111111111111111111111",
2683 => "011111111111111111111110",
2684 => "011111111111111111111111",
2685 => "011111111111111111111111",
2686 => "011111111111111111111111",
2687 => "011111111111111111111110",
2688 => "011111111111111111111111",
2689 => "011111111111111111111111",
2690 => "011111111111111111111111",
2691 => "011111111111111111111101",
2692 => "011111111111111111111111",
2693 => "011111111111111111111111",
2694 => "011111111111111111111111",
2695 => "011111111111111111111110",
2696 => "011111111111111111111111",
2697 => "011111111111111111111111",
2698 => "011111111111111111111111",
2699 => "011111111111111111111111",
2700 => "011111111111111111111111",
2701 => "011111111111111111111111",
2702 => "011111111111111111111110",
2703 => "011111111111111111111111",
2704 => "011111111111111111111111",
2705 => "011111111111111111111111",
2706 => "011111111111111111111111",
2707 => "100000000000000000000000",
2708 => "100000000000000000000000",
2709 => "100000000000000000000000",
2710 => "100000000000000000000011",
2711 => "100000000000000000000000",
2712 => "100000000000000000000000",
2713 => "100000000000000000000000",
2714 => "100000000000000000000010",
2715 => "100000000000000000000000",
2716 => "100000000000000000000000",
2717 => "100000000000000000000000",
2718 => "100000000000000000000000",
2719 => "100000000000000000000000",
2720 => "100000000000000000000010",
2721 => "100000000000000000000000",
2722 => "100000000000000000000000",
2723 => "100000000000000000000010",
2724 => "100000000000000000000001",
2725 => "100000000000000000000000",
2726 => "100000000000000000000000",
2727 => "100000000000000000000010",
2728 => "100000000000000000000000",
2729 => "100000000000000000000000",
2730 => "100000000000000000000001",
2731 => "100000000000000000000000",
2732 => "100000000000000000000000",
2733 => "100000000000000000000010",
2734 => "100000000000000000000001",
2735 => "100000000000000000000000",
2736 => "100000000000000000000000",
2737 => "100000000000000000000011",
2738 => "100000000000000000000010",
2739 => "100000000000000000000000",
2740 => "100000000000000000000000",
2741 => "100000000000000000000010",
2742 => "100000000000000000000010",
2743 => "100000000000000000000000",
2744 => "100000000000000000000000",
2745 => "100000000000000000000000",
2746 => "100000000000000000000010",
2747 => "100000000000000000000010",
2748 => "100000000000000000000000",
2749 => "100000000000000000000000",
2750 => "100000000000000000000001",
2751 => "100000000000000000000000",
2752 => "100000000000000000000000",
2753 => "100000000000000000000011",
2754 => "100000000000000000000001",
2755 => "100000000000000000000000",
2756 => "100000000000000000000000",
2757 => "100000000000000000000010",
2758 => "100000000000000000000000",
2759 => "100000000000000000000000",
2760 => "100000000000000000000000",
2761 => "100000000000000000000000",
2762 => "100000000000000000000000",
2763 => "100000000000000000000100",
2764 => "100000000000000000000000",
2765 => "100000000000000000000000",
2766 => "100000000000000000000000",
2767 => "100000000000000000000001",
2768 => "100000000000000000000010",
2769 => "100000000000000000000000",
2770 => "100000000000000000000000",
2771 => "100000000000000000000010",
2772 => "100000000000000000000010",
2773 => "100000000000000000000000",
2774 => "100000000000000000000000",
2775 => "100000000000000000000010",
2776 => "100000000000000000000000",
2777 => "100000000000000000000000",
2778 => "100000000000000000000001",
2779 => "100000000000000000000000",
2780 => "100000000000000000000000",
2781 => "100000000000000000000001",
2782 => "100000000000000000000001",
2783 => "100000000000000000000000",
2784 => "100000000000000000000000",
2785 => "100000000000000000000010",
2786 => "100000000000000000000000",
2787 => "100000000000000000000000",
2788 => "100000000000000000000010",
2789 => "100000000000000000000010",
2790 => "100000000000000000000000",
2791 => "100000000000000000000000",
2792 => "100000000000000000000011",
2793 => "100000000000000000000000",
2794 => "100000000000000000000000",
2795 => "100000000000000000000001",
2796 => "100000000000000000000100",
2797 => "100000000000000000000000",
2798 => "100000000000000000000000",
2799 => "100000000000000000000000",
2800 => "100000000000000000000010",
2801 => "100000000000000000000010",
2802 => "100000000000000000000000",
2803 => "100000000000000000000000",
2804 => "100000000000000000000000",
2805 => "100000000000000000000011",
2806 => "100000000000000000000001",
2807 => "011111111111111111111110",
2808 => "011111111111111111111111",
2809 => "011111111111111111111111",
2810 => "011111111111111111111111",
2811 => "011111111111111111111101",
2812 => "011111111111111111111111",
2813 => "011111111111111111111111",
2814 => "011111111111111111111111",
2815 => "011111111111111111111111",
2816 => "011111111111111111111110",
2817 => "011111111111111111111111",
2818 => "011111111111111111111111",
2819 => "011111111111111111111111",
2820 => "011111111111111111111100",
2821 => "011111111111111111111111",
2822 => "011111111111111111111111",
2823 => "011111111111111111111111",
2824 => "011111111111111111111110",
2825 => "011111111111111111111111",
2826 => "011111111111111111111111",
2827 => "011111111111111111111111",
2828 => "011111111111111111111111",
2829 => "011111111111111111111111",
2830 => "011111111111111111111101",
2831 => "011111111111111111111111",
2832 => "011111111111111111111111",
2833 => "011111111111111111111100",
2834 => "011111111111111111111100",
2835 => "011111111111111111111111",
2836 => "011111111111111111111111",
2837 => "011111111111111111111100",
2838 => "011111111111111111111101",
2839 => "011111111111111111111111",
2840 => "011111111111111111111111",
2841 => "011111111111111111111100",
2842 => "011111111111111111111100",
2843 => "011111111111111111111111",
2844 => "011111111111111111111111",
2845 => "011111111111111111111101",
2846 => "011111111111111111111110",
2847 => "011111111111111111111111",
2848 => "011111111111111111111111",
2849 => "011111111111111111111110",
2850 => "011111111111111111111111",
2851 => "011111111111111111111111",
2852 => "011111111111111111111110",
2853 => "011111111111111111111111",
2854 => "011111111111111111111111",
2855 => "011111111111111111111111",
2856 => "011111111111111111111110",
2857 => "011111111111111111111111",
2858 => "011111111111111111111111",
2859 => "011111111111111111111111",
2860 => "011111111111111111111111",
2861 => "011111111111111111111111",
2862 => "011111111111111111111110",
2863 => "011111111111111111111111",
2864 => "011111111111111111111111",
2865 => "011111111111111111111111",
2866 => "011111111111111111111111",
2867 => "011111111111111111111111",
2868 => "011111111111111111111111",
2869 => "011111111111111111111111",
2870 => "011111111111111111111111",
2871 => "011111111111111111111111",
2872 => "011111111111111111111111",
2873 => "011111111111111111111111",
2874 => "011111111111111111111111",
2875 => "011111111111111111111110",
2876 => "011111111111111111111111",
2877 => "011111111111111111111111",
2878 => "011111111111111111111111",
2879 => "011111111111111111111110",
2880 => "011111111111111111111110",
2881 => "011111111111111111111111",
2882 => "011111111111111111111111",
2883 => "011111111111111111111111",
2884 => "011111111111111111111110",
2885 => "011111111111111111111111",
2886 => "011111111111111111111111",
2887 => "011111111111111111111111",
2888 => "011111111111111111111111",
2889 => "011111111111111111111111",
2890 => "011111111111111111111110",
2891 => "011111111111111111111110",
2892 => "011111111111111111111111",
2893 => "011111111111111111111111",
2894 => "011111111111111111111100",
2895 => "011111111111111111111100",
2896 => "011111111111111111111111",
2897 => "011111111111111111111111",
2898 => "011111111111111111111100",
2899 => "011111111111111111111110",
2900 => "011111111111111111111111",
2901 => "011111111111111111111111",
2902 => "011111111111111111111110",
2903 => "011111111111111111111110",
2904 => "011111111111111111111111",
2905 => "011111111111111111111111",
2906 => "011111111111111111111110",
2907 => "100000000000000000000000",
2908 => "100000000000000000000010",
2909 => "100000000000000000000001",
2910 => "100000000000000000000000",
2911 => "100000000000000000000001",
2912 => "100000000000000000000010",
2913 => "100000000000000000000000",
2914 => "100000000000000000000000",
2915 => "100000000000000000000010",
2916 => "100000000000000000000000",
2917 => "100000000000000000000000",
2918 => "100000000000000000000001",
2919 => "100000000000000000000000",
2920 => "100000000000000000000000",
2921 => "100000000000000000000010",
2922 => "100000000000000000000010",
2923 => "100000000000000000000000",
2924 => "100000000000000000000000",
2925 => "100000000000000000000110",
2926 => "100000000000000000000001",
2927 => "100000000000000000000000",
2928 => "100000000000000000000000",
2929 => "100000000000000000000110",
2930 => "100000000000000000000000",
2931 => "100000000000000000000000",
2932 => "100000000000000000000001",
2933 => "100000000000000000000100",
2934 => "100000000000000000000000",
2935 => "100000000000000000000000",
2936 => "100000000000000000000000",
2937 => "100000000000000000000010",
2938 => "100000000000000000000010",
2939 => "100000000000000000000000",
2940 => "100000000000000000000000",
2941 => "100000000000000000000001",
2942 => "100000000000000000000010",
2943 => "100000000000000000000000",
2944 => "100000000000000000000000",
2945 => "100000000000000000000000",
2946 => "100000000000000000000001",
2947 => "100000000000000000000000",
2948 => "100000000000000000000000",
2949 => "100000000000000000000000",
2950 => "100000000000000000000001",
2951 => "100000000000000000000000",
2952 => "100000000000000000000000",
2953 => "100000000000000000000000",
2954 => "100000000000000000000000",
2955 => "100000000000000000000000",
2956 => "100000000000000000000000",
2957 => "100000000000000000000000",
2958 => "100000000000000000000000",
2959 => "100000000000000000000000",
2960 => "100000000000000000000000",
2961 => "100000000000000000000000",
2962 => "100000000000000000000010",
2963 => "100000000000000000000010",
2964 => "100000000000000000000000",
2965 => "100000000000000000000000",
2966 => "100000000000000000000010",
2967 => "100000000000000000000010",
2968 => "100000000000000000000000",
2969 => "100000000000000000000000",
2970 => "100000000000000000000000",
2971 => "100000000000000000000000",
2972 => "100000000000000000000001",
2973 => "100000000000000000000000",
2974 => "100000000000000000000000",
2975 => "100000000000000000000000",
2976 => "100000000000000000000000",
2977 => "100000000000000000000001",
2978 => "100000000000000000000010",
2979 => "100000000000000000000000",
2980 => "100000000000000000000000",
2981 => "100000000000000000000000",
2982 => "100000000000000000000001",
2983 => "100000000000000000000000",
2984 => "100000000000000000000000",
2985 => "100000000000000000000000",
2986 => "100000000000000000000000",
2987 => "100000000000000000000010",
2988 => "100000000000000000000000",
2989 => "100000000000000000000000",
2990 => "100000000000000000000001",
2991 => "100000000000000000000000",
2992 => "100000000000000000000000",
2993 => "100000000000000000000010",
2994 => "100000000000000000000000",
2995 => "100000000000000000000000",
2996 => "100000000000000000000000",
2997 => "100000000000000000000100",
2998 => "100000000000000000000000",
2999 => "100000000000000000000000",
3000 => "100000000000000000000010",
3001 => "100000000000000000000010",
3002 => "100000000000000000000000",
3003 => "100000000000000000000000",
3004 => "100000000000000000000010",
3005 => "100000000000000000000000",
3006 => "100000000000000000000000",
3007 => "011111111111111111111111",
3008 => "011111111111111111111111",
3009 => "011111111111111111111111",
3010 => "011111111111111111111100",
3011 => "011111111111111111111111",
3012 => "011111111111111111111111",
3013 => "011111111111111111111111",
3014 => "011111111111111111111110",
3015 => "011111111111111111111111",
3016 => "011111111111111111111111",
3017 => "011111111111111111111111",
3018 => "011111111111111111111111",
3019 => "011111111111111111111111",
3020 => "011111111111111111111111",
3021 => "011111111111111111111111",
3022 => "011111111111111111111111",
3023 => "011111111111111111111110",
3024 => "011111111111111111111111",
3025 => "011111111111111111111111",
3026 => "011111111111111111111111",
3027 => "011111111111111111111100",
3028 => "011111111111111111111111",
3029 => "011111111111111111111111",
3030 => "011111111111111111111110",
3031 => "011111111111111111111111",
3032 => "011111111111111111111111",
3033 => "011111111111111111111111",
3034 => "011111111111111111111110",
3035 => "011111111111111111111111",
3036 => "011111111111111111111111",
3037 => "011111111111111111111110",
3038 => "011111111111111111111110",
3039 => "011111111111111111111111",
3040 => "011111111111111111111111",
3041 => "011111111111111111111110",
3042 => "011111111111111111111111",
3043 => "011111111111111111111111",
3044 => "011111111111111111111111",
3045 => "011111111111111111111100",
3046 => "011111111111111111111111",
3047 => "011111111111111111111111",
3048 => "011111111111111111111111",
3049 => "011111111111111111111110",
3050 => "011111111111111111111111",
3051 => "011111111111111111111111",
3052 => "011111111111111111111111",
3053 => "011111111111111111111111",
3054 => "011111111111111111111111",
3055 => "011111111111111111111111",
3056 => "011111111111111111111111",
3057 => "011111111111111111111110",
3058 => "011111111111111111111111",
3059 => "011111111111111111111111",
3060 => "011111111111111111111110",
3061 => "011111111111111111111010",
3062 => "011111111111111111111111",
3063 => "011111111111111111111111",
3064 => "011111111111111111111110",
3065 => "011111111111111111111010",
3066 => "011111111111111111111111",
3067 => "011111111111111111111111",
3068 => "011111111111111111111111",
3069 => "011111111111111111111111",
3070 => "011111111111111111111110",
3071 => "011111111111111111111111",
3072 => "011111111111111111111111",
3073 => "011111111111111111111111",
3074 => "011111111111111111111100",
3075 => "011111111111111111111111",
3076 => "011111111111111111111111",
3077 => "011111111111111111111111",
3078 => "011111111111111111111110",
3079 => "011111111111111111111110",
3080 => "011111111111111111111111",
3081 => "011111111111111111111111",
3082 => "011111111111111111111111",
3083 => "011111111111111111111100",
3084 => "011111111111111111111110",
3085 => "011111111111111111111111",
3086 => "011111111111111111111111",
3087 => "011111111111111111111110",
3088 => "011111111111111111111111",
3089 => "011111111111111111111111",
3090 => "011111111111111111111111",
3091 => "011111111111111111111110",
3092 => "011111111111111111111111",
3093 => "011111111111111111111111",
3094 => "011111111111111111111110",
3095 => "011111111111111111111110",
3096 => "011111111111111111111111",
3097 => "011111111111111111111111",
3098 => "011111111111111111111111",
3099 => "011111111111111111111111",
3100 => "011111111111111111111110",
3101 => "011111111111111111111111",
3102 => "011111111111111111111111",
3103 => "011111111111111111111111",
3104 => "011111111111111111111011",
3105 => "011111111111111111111111",
3106 => "011111111111111111111111",
3107 => "100000000000000000000000",
3108 => "100000000000000000000000",
3109 => "100000000000000000000100",
3110 => "100000000000000000000000",
3111 => "100000000000000000000000",
3112 => "100000000000000000000010",
3113 => "100000000000000000000100",
3114 => "100000000000000000000000",
3115 => "100000000000000000000000",
3116 => "100000000000000000000010",
3117 => "100000000000000000000001",
3118 => "100000000000000000000000",
3119 => "100000000000000000000000",
3120 => "100000000000000000000100",
3121 => "100000000000000000000000",
3122 => "100000000000000000000000",
3123 => "100000000000000000000001",
3124 => "100000000000000000000011",
3125 => "100000000000000000000000",
3126 => "100000000000000000000000",
3127 => "100000000000000000000001",
3128 => "100000000000000000000001",
3129 => "100000000000000000000000",
3130 => "100000000000000000000000",
3131 => "100000000000000000000000",
3132 => "100000000000000000000000",
3133 => "100000000000000000000001",
3134 => "100000000000000000000000",
3135 => "100000000000000000000000",
3136 => "100000000000000000000001",
3137 => "100000000000000000000010",
3138 => "100000000000000000000000",
3139 => "100000000000000000000000",
3140 => "100000000000000000000010",
3141 => "100000000000000000000010",
3142 => "100000000000000000000000",
3143 => "100000000000000000000000",
3144 => "100000000000000000000011",
3145 => "100000000000000000000001",
3146 => "100000000000000000000000",
3147 => "100000000000000000000000",
3148 => "100000000000000000000100",
3149 => "100000000000000000000000",
3150 => "100000000000000000000000",
3151 => "100000000000000000000000",
3152 => "100000000000000000000100",
3153 => "100000000000000000000000",
3154 => "100000000000000000000000",
3155 => "100000000000000000000000",
3156 => "100000000000000000000100",
3157 => "100000000000000000000000",
3158 => "100000000000000000000000",
3159 => "100000000000000000000010",
3160 => "100000000000000000000100",
3161 => "100000000000000000000000",
3162 => "100000000000000000000000",
3163 => "100000000000000000000010",
3164 => "100000000000000000000010",
3165 => "100000000000000000000000",
3166 => "100000000000000000000000",
3167 => "100000000000000000000000",
3168 => "100000000000000000000010",
3169 => "100000000000000000000000",
3170 => "100000000000000000000000",
3171 => "100000000000000000000000",
3172 => "100000000000000000000100",
3173 => "100000000000000000000001",
3174 => "100000000000000000000000",
3175 => "100000000000000000000000",
3176 => "100000000000000000000100",
3177 => "100000000000000000000000",
3178 => "100000000000000000000000",
3179 => "100000000000000000000000",
3180 => "100000000000000000000100",
3181 => "100000000000000000000000",
3182 => "100000000000000000000000",
3183 => "100000000000000000000001",
3184 => "100000000000000000000011",
3185 => "100000000000000000000000",
3186 => "100000000000000000000000",
3187 => "100000000000000000000001",
3188 => "100000000000000000000010",
3189 => "100000000000000000000000",
3190 => "100000000000000000000000",
3191 => "100000000000000000000001",
3192 => "100000000000000000000001",
3193 => "100000000000000000000000",
3194 => "100000000000000000000000",
3195 => "100000000000000000000010",
3196 => "100000000000000000000000",
3197 => "100000000000000000000000",
3198 => "100000000000000000000010",
3199 => "100000000000000000000010",
3200 => "100000000000000000000000",
3201 => "100000000000000000000000",
3202 => "100000000000000000000001",
3203 => "100000000000000000000010",
3204 => "100000000000000000000001",
3205 => "100000000000000000000000",
3206 => "100000000000000000000000",
3207 => "011111111111111111111111",
3208 => "011111111111111111111111",
3209 => "011111111111111111111111",
3210 => "011111111111111111111111",
3211 => "011111111111111111111111",
3212 => "011111111111111111111100",
3213 => "011111111111111111111111",
3214 => "011111111111111111111111",
3215 => "011111111111111111111111",
3216 => "011111111111111111111011",
3217 => "011111111111111111111111",
3218 => "011111111111111111111111",
3219 => "011111111111111111111110",
3220 => "011111111111111111111101",
3221 => "011111111111111111111111",
3222 => "011111111111111111111111",
3223 => "011111111111111111111110",
3224 => "011111111111111111111110",
3225 => "011111111111111111111111",
3226 => "011111111111111111111111",
3227 => "011111111111111111111111",
3228 => "011111111111111111111111",
3229 => "011111111111111111111111",
3230 => "011111111111111111111110",
3231 => "011111111111111111111111",
3232 => "011111111111111111111111",
3233 => "011111111111111111111111",
3234 => "011111111111111111111110",
3235 => "011111111111111111111111",
3236 => "011111111111111111111111",
3237 => "011111111111111111111111",
3238 => "011111111111111111111110",
3239 => "011111111111111111111110",
3240 => "011111111111111111111111",
3241 => "011111111111111111111111",
3242 => "011111111111111111111100",
3243 => "011111111111111111111111",
3244 => "011111111111111111111111",
3245 => "011111111111111111111111",
3246 => "011111111111111111111110",
3247 => "011111111111111111111111",
3248 => "011111111111111111111111",
3249 => "011111111111111111111111",
3250 => "011111111111111111111111",
3251 => "011111111111111111111111",
3252 => "011111111111111111111111",
3253 => "011111111111111111111111",
3254 => "011111111111111111111111",
3255 => "011111111111111111111111",
3256 => "011111111111111111111111",
3257 => "011111111111111111111110",
3258 => "011111111111111111111111",
3259 => "011111111111111111111111",
3260 => "011111111111111111111111",
3261 => "011111111111111111111110",
3262 => "011111111111111111111111",
3263 => "011111111111111111111111",
3264 => "011111111111111111111110",
3265 => "011111111111111111111111",
3266 => "011111111111111111111111",
3267 => "011111111111111111111111",
3268 => "011111111111111111111110",
3269 => "011111111111111111111111",
3270 => "011111111111111111111111",
3271 => "011111111111111111111111",
3272 => "011111111111111111111111",
3273 => "011111111111111111111111",
3274 => "011111111111111111111111",
3275 => "011111111111111111111111",
3276 => "011111111111111111111110",
3277 => "011111111111111111111111",
3278 => "011111111111111111111111",
3279 => "011111111111111111111111",
3280 => "011111111111111111111110",
3281 => "011111111111111111111111",
3282 => "011111111111111111111111",
3283 => "011111111111111111111110",
3284 => "011111111111111111111111",
3285 => "011111111111111111111111",
3286 => "011111111111111111111110",
3287 => "011111111111111111111100",
3288 => "011111111111111111111111",
3289 => "011111111111111111111111",
3290 => "011111111111111111111111",
3291 => "011111111111111111111110",
3292 => "011111111111111111111111",
3293 => "011111111111111111111111",
3294 => "011111111111111111111111",
3295 => "011111111111111111111111",
3296 => "011111111111111111111111",
3297 => "011111111111111111111110",
3298 => "011111111111111111111111",
3299 => "011111111111111111111111",
3300 => "011111111111111111111111",
3301 => "011111111111111111111110",
3302 => "011111111111111111111111",
3303 => "011111111111111111111111",
3304 => "011111111111111111111110",
3305 => "011111111111111111111111",
3306 => "011111111111111111111111",
3307 => "100000000000000000000000",
3308 => "100000000000000000000000",
3309 => "100000000000000000000000",
3310 => "100000000000000000000110",
3311 => "100000000000000000000001",
3312 => "100000000000000000000000",
3313 => "100000000000000000000000",
3314 => "100000000000000000000100",
3315 => "100000000000000000000001",
3316 => "100000000000000000000000",
3317 => "100000000000000000000000",
3318 => "100000000000000000000101",
3319 => "100000000000000000000000",
3320 => "100000000000000000000000",
3321 => "100000000000000000000100",
3322 => "100000000000000000000110",
3323 => "100000000000000000000000",
3324 => "100000000000000000000000",
3325 => "100000000000000000000110",
3326 => "100000000000000000000010",
3327 => "100000000000000000000000",
3328 => "100000000000000000000000",
3329 => "100000000000000000000100",
3330 => "100000000000000000000000",
3331 => "100000000000000000000000",
3332 => "100000000000000000000000",
3333 => "100000000000000000000010",
3334 => "100000000000000000000001",
3335 => "100000000000000000000000",
3336 => "100000000000000000000000",
3337 => "100000000000000000000010",
3338 => "100000000000000000000010",
3339 => "100000000000000000000000",
3340 => "100000000000000000000000",
3341 => "100000000000000000000001",
3342 => "100000000000000000000100",
3343 => "100000000000000000000000",
3344 => "100000000000000000000000",
3345 => "100000000000000000000000",
3346 => "100000000000000000000010",
3347 => "100000000000000000000000",
3348 => "100000000000000000000000",
3349 => "100000000000000000000000",
3350 => "100000000000000000000000",
3351 => "100000000000000000000000",
3352 => "100000000000000000000010",
3353 => "100000000000000000000000",
3354 => "100000000000000000000000",
3355 => "100000000000000000000000",
3356 => "100000000000000000000001",
3357 => "100000000000000000000000",
3358 => "100000000000000000000000",
3359 => "100000000000000000000010",
3360 => "100000000000000000000000",
3361 => "100000000000000000000000",
3362 => "100000000000000000000000",
3363 => "100000000000000000000010",
3364 => "100000000000000000000000",
3365 => "100000000000000000000000",
3366 => "100000000000000000000010",
3367 => "100000000000000000000001",
3368 => "100000000000000000000000",
3369 => "100000000000000000000000",
3370 => "100000000000000000000100",
3371 => "100000000000000000000001",
3372 => "100000000000000000000000",
3373 => "100000000000000000000000",
3374 => "100000000000000000000010",
3375 => "100000000000000000000001",
3376 => "100000000000000000000000",
3377 => "100000000000000000000000",
3378 => "100000000000000000000000",
3379 => "100000000000000000000000",
3380 => "100000000000000000000010",
3381 => "100000000000000000000001",
3382 => "100000000000000000000000",
3383 => "100000000000000000000000",
3384 => "100000000000000000000010",
3385 => "100000000000000000000010",
3386 => "100000000000000000000000",
3387 => "100000000000000000000000",
3388 => "100000000000000000000010",
3389 => "100000000000000000000100",
3390 => "100000000000000000000000",
3391 => "100000000000000000000000",
3392 => "100000000000000000000001",
3393 => "100000000000000000000100",
3394 => "100000000000000000000000",
3395 => "100000000000000000000000",
3396 => "100000000000000000000001",
3397 => "100000000000000000000100",
3398 => "100000000000000000000000",
3399 => "100000000000000000000000",
3400 => "100000000000000000000100",
3401 => "100000000000000000000010",
3402 => "100000000000000000000000",
3403 => "100000000000000000000000",
3404 => "100000000000000000000110",
3405 => "100000000000000000000000",
3406 => "100000000000000000000000",
3407 => "011111111111111111111111",
3408 => "011111111111111111111111",
3409 => "011111111111111111111111",
3410 => "011111111111111111111110",
3411 => "011111111111111111111110",
3412 => "011111111111111111111111",
3413 => "011111111111111111111111",
3414 => "011111111111111111111110",
3415 => "011111111111111111111110",
3416 => "011111111111111111111111",
3417 => "011111111111111111111111",
3418 => "011111111111111111111100",
3419 => "011111111111111111111111",
3420 => "011111111111111111111111",
3421 => "011111111111111111111111",
3422 => "011111111111111111111110",
3423 => "011111111111111111111111",
3424 => "011111111111111111111111",
3425 => "011111111111111111111111",
3426 => "011111111111111111111111",
3427 => "011111111111111111111111",
3428 => "011111111111111111111110",
3429 => "011111111111111111111110",
3430 => "011111111111111111111111",
3431 => "011111111111111111111111",
3432 => "011111111111111111111110",
3433 => "011111111111111111111100",
3434 => "011111111111111111111111",
3435 => "011111111111111111111111",
3436 => "011111111111111111111110",
3437 => "011111111111111111111110",
3438 => "011111111111111111111111",
3439 => "011111111111111111111111",
3440 => "011111111111111111111111",
3441 => "011111111111111111111111",
3442 => "011111111111111111111111",
3443 => "011111111111111111111111",
3444 => "011111111111111111111111",
3445 => "011111111111111111111111",
3446 => "011111111111111111111111",
3447 => "011111111111111111111110",
3448 => "011111111111111111111111",
3449 => "011111111111111111111111",
3450 => "011111111111111111111111",
3451 => "011111111111111111111110",
3452 => "011111111111111111111111",
3453 => "011111111111111111111111",
3454 => "011111111111111111111111",
3455 => "011111111111111111111111",
3456 => "011111111111111111111111",
3457 => "011111111111111111111111",
3458 => "011111111111111111111111",
3459 => "011111111111111111111111",
3460 => "011111111111111111111111",
3461 => "011111111111111111111111",
3462 => "011111111111111111111110",
3463 => "011111111111111111111111",
3464 => "011111111111111111111111",
3465 => "011111111111111111111111",
3466 => "011111111111111111111111",
3467 => "011111111111111111111111",
3468 => "011111111111111111111110",
3469 => "011111111111111111111111",
3470 => "011111111111111111111111",
3471 => "011111111111111111111111",
3472 => "011111111111111111111100",
3473 => "011111111111111111111111",
3474 => "011111111111111111111111",
3475 => "011111111111111111111111",
3476 => "011111111111111111111110",
3477 => "011111111111111111111111",
3478 => "011111111111111111111111",
3479 => "011111111111111111111111",
3480 => "011111111111111111111111",
3481 => "011111111111111111111111",
3482 => "011111111111111111111111",
3483 => "011111111111111111111111",
3484 => "011111111111111111111111",
3485 => "011111111111111111111111",
3486 => "011111111111111111111111",
3487 => "011111111111111111111111",
3488 => "011111111111111111111100",
3489 => "011111111111111111111111",
3490 => "011111111111111111111111",
3491 => "011111111111111111111111",
3492 => "011111111111111111111101",
3493 => "011111111111111111111111",
3494 => "011111111111111111111111",
3495 => "011111111111111111111111",
3496 => "011111111111111111111110",
3497 => "011111111111111111111111",
3498 => "011111111111111111111111",
3499 => "011111111111111111111111",
3500 => "011111111111111111111110",
3501 => "011111111111111111111111",
3502 => "011111111111111111111111",
3503 => "011111111111111111111111",
3504 => "011111111111111111111100",
3505 => "011111111111111111111111",
3506 => "011111111111111111111111",
3507 => "100000000000000000000000",
3508 => "100000000000000000000000",
3509 => "100000000000000000000000",
3510 => "100000000000000000000010",
3511 => "100000000000000000000000",
3512 => "100000000000000000000000",
3513 => "100000000000000000000010",
3514 => "100000000000000000000000",
3515 => "100000000000000000000000",
3516 => "100000000000000000000000",
3517 => "100000000000000000000010",
3518 => "100000000000000000000001",
3519 => "100000000000000000000000",
3520 => "100000000000000000000000",
3521 => "100000000000000000000001",
3522 => "100000000000000000000000",
3523 => "100000000000000000000000",
3524 => "100000000000000000000000",
3525 => "100000000000000000000010",
3526 => "100000000000000000000000",
3527 => "100000000000000000000000",
3528 => "100000000000000000000010",
3529 => "100000000000000000000000",
3530 => "100000000000000000000000",
3531 => "100000000000000000000001",
3532 => "100000000000000000000010",
3533 => "100000000000000000000000",
3534 => "100000000000000000000000",
3535 => "100000000000000000000010",
3536 => "100000000000000000000011",
3537 => "100000000000000000000000",
3538 => "100000000000000000000000",
3539 => "100000000000000000000010",
3540 => "100000000000000000000010",
3541 => "100000000000000000000000",
3542 => "100000000000000000000000",
3543 => "100000000000000000000100",
3544 => "100000000000000000000000",
3545 => "100000000000000000000000",
3546 => "100000000000000000000001",
3547 => "100000000000000000000010",
3548 => "100000000000000000000000",
3549 => "100000000000000000000000",
3550 => "100000000000000000000010",
3551 => "100000000000000000000000",
3552 => "100000000000000000000000",
3553 => "100000000000000000000100",
3554 => "100000000000000000000010",
3555 => "100000000000000000000000",
3556 => "100000000000000000000000",
3557 => "100000000000000000000010",
3558 => "100000000000000000000100",
3559 => "100000000000000000000000",
3560 => "100000000000000000000000",
3561 => "100000000000000000000000",
3562 => "100000000000000000000011",
3563 => "100000000000000000000000",
3564 => "100000000000000000000000",
3565 => "100000000000000000000010",
3566 => "100000000000000000000000",
3567 => "100000000000000000000000",
3568 => "100000000000000000000001",
3569 => "100000000000000000000100",
3570 => "100000000000000000000000",
3571 => "100000000000000000000000",
3572 => "100000000000000000000010",
3573 => "100000000000000000000010",
3574 => "100000000000000000000000",
3575 => "100000000000000000000000",
3576 => "100000000000000000000100",
3577 => "100000000000000000000000",
3578 => "100000000000000000000000",
3579 => "100000000000000000000000",
3580 => "100000000000000000000011",
3581 => "100000000000000000000000",
3582 => "100000000000000000000000",
3583 => "100000000000000000000000",
3584 => "100000000000000000000000",
3585 => "100000000000000000000000",
3586 => "100000000000000000000010",
3587 => "100000000000000000000000",
3588 => "100000000000000000000000",
3589 => "100000000000000000000000",
3590 => "100000000000000000000100",
3591 => "100000000000000000000000",
3592 => "100000000000000000000000",
3593 => "100000000000000000000000",
3594 => "100000000000000000000101",
3595 => "100000000000000000000000",
3596 => "100000000000000000000000",
3597 => "100000000000000000000001",
3598 => "100000000000000000000001",
3599 => "100000000000000000000000",
3600 => "100000000000000000000000",
3601 => "100000000000000000000010",
3602 => "100000000000000000000000",
3603 => "100000000000000000000000",
3604 => "100000000000000000000011",
3605 => "100000000000000000000010",
3606 => "100000000000000000000000",
3607 => "100000000000000000000000",
3608 => "100000000000000000000010",
3609 => "011111111111111111111111",
3610 => "011111111111111111111110",
3611 => "011111111111111111111111",
3612 => "011111111111111111111111",
3613 => "011111111111111111111111",
3614 => "011111111111111111111111",
3615 => "011111111111111111111111",
3616 => "011111111111111111111110",
3617 => "011111111111111111111110",
3618 => "011111111111111111111111",
3619 => "011111111111111111111111",
3620 => "011111111111111111111111",
3621 => "011111111111111111111111",
3622 => "011111111111111111111110",
3623 => "011111111111111111111111",
3624 => "011111111111111111111111",
3625 => "011111111111111111111111",
3626 => "011111111111111111111110",
3627 => "011111111111111111111111",
3628 => "011111111111111111111111",
3629 => "011111111111111111111111",
3630 => "011111111111111111111110",
3631 => "011111111111111111111111",
3632 => "011111111111111111111111",
3633 => "011111111111111111111110",
3634 => "011111111111111111111110",
3635 => "011111111111111111111111",
3636 => "011111111111111111111111",
3637 => "011111111111111111111101",
3638 => "011111111111111111111110",
3639 => "011111111111111111111111",
3640 => "011111111111111111111111",
3641 => "011111111111111111111110",
3642 => "011111111111111111111111",
3643 => "011111111111111111111111",
3644 => "011111111111111111111111",
3645 => "011111111111111111111110",
3646 => "011111111111111111111111",
3647 => "011111111111111111111111",
3648 => "011111111111111111111111",
3649 => "011111111111111111111110",
3650 => "011111111111111111111111",
3651 => "011111111111111111111111",
3652 => "011111111111111111111111",
3653 => "011111111111111111111110",
3654 => "011111111111111111111111",
3655 => "011111111111111111111111",
3656 => "011111111111111111111111",
3657 => "011111111111111111111110",
3658 => "011111111111111111111111",
3659 => "011111111111111111111111",
3660 => "011111111111111111111111",
3661 => "011111111111111111111111",
3662 => "011111111111111111111101",
3663 => "011111111111111111111100",
3664 => "011111111111111111111111",
3665 => "011111111111111111111111",
3666 => "011111111111111111111101",
3667 => "011111111111111111111100",
3668 => "011111111111111111111111",
3669 => "011111111111111111111111",
3670 => "011111111111111111111111",
3671 => "011111111111111111111111",
3672 => "011111111111111111111111",
3673 => "011111111111111111111111",
3674 => "011111111111111111111111",
3675 => "011111111111111111111111",
3676 => "011111111111111111111111",
3677 => "011111111111111111111111",
3678 => "011111111111111111111111",
3679 => "011111111111111111111111",
3680 => "011111111111111111111111",
3681 => "011111111111111111111111",
3682 => "011111111111111111111110",
3683 => "011111111111111111111111",
3684 => "011111111111111111111111",
3685 => "011111111111111111111110",
3686 => "011111111111111111111010",
3687 => "011111111111111111111111",
3688 => "011111111111111111111111",
3689 => "011111111111111111111011",
3690 => "011111111111111111111100",
3691 => "011111111111111111111111",
3692 => "011111111111111111111111",
3693 => "011111111111111111111110",
3694 => "011111111111111111111110",
3695 => "011111111111111111111111",
3696 => "011111111111111111111111",
3697 => "011111111111111111111111",
3698 => "011111111111111111111110",
3699 => "011111111111111111111110",
3700 => "011111111111111111111111",
3701 => "011111111111111111111111",
3702 => "011111111111111111111111",
3703 => "011111111111111111111111",
3704 => "011111111111111111111111",
3705 => "011111111111111111111111",
3706 => "011111111111111111111110",
3707 => "011111111111111111111111",
3708 => "011111111111111111111111",
3709 => "100000000000000000000010",
3710 => "100000000000000000000000",
3711 => "100000000000000000000000",
3712 => "100000000000000000000100",
3713 => "100000000000000000000001",
3714 => "100000000000000000000000",
3715 => "100000000000000000000000",
3716 => "100000000000000000000010",
3717 => "100000000000000000000000",
3718 => "100000000000000000000000",
3719 => "100000000000000000000000",
3720 => "100000000000000000000001",
3721 => "100000000000000000000001",
3722 => "100000000000000000000000",
3723 => "100000000000000000000000",
3724 => "100000000000000000000100",
3725 => "100000000000000000000010",
3726 => "100000000000000000000000",
3727 => "100000000000000000000000",
3728 => "100000000000000000000011",
3729 => "100000000000000000000000",
3730 => "100000000000000000000000",
3731 => "100000000000000000000000",
3732 => "100000000000000000000000",
3733 => "100000000000000000000001",
3734 => "100000000000000000000010",
3735 => "100000000000000000000000",
3736 => "100000000000000000000000",
3737 => "100000000000000000000010",
3738 => "100000000000000000000001",
3739 => "100000000000000000000000",
3740 => "100000000000000000000000",
3741 => "100000000000000000000010",
3742 => "100000000000000000000000",
3743 => "100000000000000000000000",
3744 => "100000000000000000000000",
3745 => "100000000000000000000011",
3746 => "100000000000000000000000",
3747 => "100000000000000000000000",
3748 => "100000000000000000000000",
3749 => "100000000000000000000010",
3750 => "100000000000000000000000",
3751 => "100000000000000000000000",
3752 => "100000000000000000000001",
3753 => "100000000000000000000000",
3754 => "100000000000000000000000",
3755 => "100000000000000000000000",
3756 => "100000000000000000000010",
3757 => "100000000000000000000000",
3758 => "100000000000000000000000",
3759 => "100000000000000000000000",
3760 => "100000000000000000000000",
3761 => "100000000000000000000001",
3762 => "100000000000000000000000",
3763 => "100000000000000000000000",
3764 => "100000000000000000000000",
3765 => "100000000000000000000000",
3766 => "100000000000000000000001",
3767 => "100000000000000000000001",
3768 => "100000000000000000000000",
3769 => "100000000000000000000000",
3770 => "100000000000000000000010",
3771 => "100000000000000000000010",
3772 => "100000000000000000000000",
3773 => "100000000000000000000000",
3774 => "100000000000000000000001",
3775 => "100000000000000000000001",
3776 => "100000000000000000000000",
3777 => "100000000000000000000001",
3778 => "100000000000000000000000",
3779 => "100000000000000000000000",
3780 => "100000000000000000000000",
3781 => "100000000000000000000010",
3782 => "100000000000000000000000",
3783 => "100000000000000000000000",
3784 => "100000000000000000000000",
3785 => "100000000000000000000001",
3786 => "100000000000000000000000",
3787 => "100000000000000000000000",
3788 => "100000000000000000000010",
3789 => "100000000000000000000000",
3790 => "100000000000000000000000",
3791 => "100000000000000000000000",
3792 => "100000000000000000000011",
3793 => "100000000000000000000000",
3794 => "100000000000000000000000",
3795 => "100000000000000000000000",
3796 => "100000000000000000000010",
3797 => "100000000000000000000000",
3798 => "100000000000000000000000",
3799 => "100000000000000000000010",
3800 => "100000000000000000000000",
3801 => "100000000000000000000000",
3802 => "100000000000000000000000",
3803 => "100000000000000000000011",
3804 => "100000000000000000000000",
3805 => "100000000000000000000000",
3806 => "100000000000000000000000",
3807 => "100000000000000000000010",
3808 => "100000000000000000000000",
3809 => "011111111111111111111111",
3810 => "011111111111111111111111",
3811 => "011111111111111111111111",
3812 => "011111111111111111111110",
3813 => "011111111111111111111111",
3814 => "011111111111111111111111",
3815 => "011111111111111111111101",
3816 => "011111111111111111111110",
3817 => "011111111111111111111111",
3818 => "011111111111111111111111",
3819 => "011111111111111111111110",
3820 => "011111111111111111111110",
3821 => "011111111111111111111111",
3822 => "011111111111111111111111",
3823 => "011111111111111111111111",
3824 => "011111111111111111111111",
3825 => "011111111111111111111111",
3826 => "011111111111111111111110",
3827 => "011111111111111111111111",
3828 => "011111111111111111111111",
3829 => "011111111111111111111111",
3830 => "011111111111111111111110",
3831 => "011111111111111111111111",
3832 => "011111111111111111111111",
3833 => "011111111111111111111111",
3834 => "011111111111111111111111",
3835 => "011111111111111111111111",
3836 => "011111111111111111111110",
3837 => "011111111111111111111111",
3838 => "011111111111111111111111",
3839 => "011111111111111111111101",
3840 => "011111111111111111111110",
3841 => "011111111111111111111111",
3842 => "011111111111111111111111",
3843 => "011111111111111111111111",
3844 => "011111111111111111111111",
3845 => "011111111111111111111111",
3846 => "011111111111111111111110",
3847 => "011111111111111111111111",
3848 => "011111111111111111111111",
3849 => "011111111111111111111111",
3850 => "011111111111111111111100",
3851 => "011111111111111111111111",
3852 => "011111111111111111111111",
3853 => "011111111111111111111111",
3854 => "011111111111111111111101",
3855 => "011111111111111111111111",
3856 => "011111111111111111111111",
3857 => "011111111111111111111111",
3858 => "011111111111111111111110",
3859 => "011111111111111111111110",
3860 => "011111111111111111111111",
3861 => "011111111111111111111111",
3862 => "011111111111111111111111",
3863 => "011111111111111111111111",
3864 => "011111111111111111111111",
3865 => "011111111111111111111110",
3866 => "011111111111111111111111",
3867 => "011111111111111111111111",
3868 => "011111111111111111111110",
3869 => "011111111111111111111100",
3870 => "011111111111111111111111",
3871 => "011111111111111111111111",
3872 => "011111111111111111111111",
3873 => "011111111111111111111111",
3874 => "011111111111111111111111",
3875 => "011111111111111111111110",
3876 => "011111111111111111111110",
3877 => "011111111111111111111111",
3878 => "011111111111111111111111",
3879 => "011111111111111111111111",
3880 => "011111111111111111111110",
3881 => "011111111111111111111110",
3882 => "011111111111111111111111",
3883 => "011111111111111111111111",
3884 => "011111111111111111111111",
3885 => "011111111111111111111100",
3886 => "011111111111111111111110",
3887 => "011111111111111111111111",
3888 => "011111111111111111111111",
3889 => "011111111111111111111110",
3890 => "011111111111111111111101",
3891 => "011111111111111111111111",
3892 => "011111111111111111111111",
3893 => "011111111111111111111110",
3894 => "011111111111111111111110",
3895 => "011111111111111111111111",
3896 => "011111111111111111111111",
3897 => "011111111111111111111110",
3898 => "011111111111111111111111",
3899 => "011111111111111111111111",
3900 => "011111111111111111111111",
3901 => "011111111111111111111110",
3902 => "011111111111111111111111",
3903 => "011111111111111111111111",
3904 => "011111111111111111111111",
3905 => "011111111111111111111111",
3906 => "011111111111111111111111",
3907 => "011111111111111111111111",
3908 => "011111111111111111111111",
3909 => "100000000000000000000000",
3910 => "100000000000000000000001",
3911 => "100000000000000000000000",
3912 => "100000000000000000000000",
3913 => "100000000000000000000000",
3914 => "100000000000000000000010",
3915 => "100000000000000000000001",
3916 => "100000000000000000000000",
3917 => "100000000000000000000000",
3918 => "100000000000000000000010",
3919 => "100000000000000000000001",
3920 => "100000000000000000000000",
3921 => "100000000000000000000000",
3922 => "100000000000000000000010",
3923 => "100000000000000000000000",
3924 => "100000000000000000000000",
3925 => "100000000000000000000010",
3926 => "100000000000000000000011",
3927 => "100000000000000000000000",
3928 => "100000000000000000000000",
3929 => "100000000000000000000011",
3930 => "100000000000000000000001",
3931 => "100000000000000000000000",
3932 => "100000000000000000000000",
3933 => "100000000000000000000010",
3934 => "100000000000000000000000",
3935 => "100000000000000000000000",
3936 => "100000000000000000000000",
3937 => "100000000000000000000000",
3938 => "100000000000000000000010",
3939 => "100000000000000000000010",
3940 => "100000000000000000000000",
3941 => "100000000000000000000000",
3942 => "100000000000000000000100",
3943 => "100000000000000000000100",
3944 => "100000000000000000000000",
3945 => "100000000000000000000000",
3946 => "100000000000000000000100",
3947 => "100000000000000000000100",
3948 => "100000000000000000000000",
3949 => "100000000000000000000000",
3950 => "100000000000000000000010",
3951 => "100000000000000000000100",
3952 => "100000000000000000000000",
3953 => "100000000000000000000000",
3954 => "100000000000000000000000",
3955 => "100000000000000000000010",
3956 => "100000000000000000000010",
3957 => "100000000000000000000000",
3958 => "100000000000000000000000",
3959 => "100000000000000000000000",
3960 => "100000000000000000000001",
3961 => "100000000000000000000011",
3962 => "100000000000000000000000",
3963 => "100000000000000000000000",
3964 => "100000000000000000000000",
3965 => "100000000000000000000000",
3966 => "100000000000000000000001",
3967 => "100000000000000000000100",
3968 => "100000000000000000000000",
3969 => "100000000000000000000000",
3970 => "100000000000000000000000",
3971 => "100000000000000000000010",
3972 => "100000000000000000000000",
3973 => "100000000000000000000000",
3974 => "100000000000000000000000",
3975 => "100000000000000000000000",
3976 => "100000000000000000000010",
3977 => "100000000000000000000011",
3978 => "100000000000000000000000",
3979 => "100000000000000000000000",
3980 => "100000000000000000000100",
3981 => "100000000000000000000010",
3982 => "100000000000000000000000",
3983 => "100000000000000000000000",
3984 => "100000000000000000000000",
3985 => "100000000000000000000010",
3986 => "100000000000000000000010",
3987 => "100000000000000000000000",
3988 => "100000000000000000000000",
3989 => "100000000000000000000001",
3990 => "100000000000000000000100",
3991 => "100000000000000000000000",
3992 => "100000000000000000000000",
3993 => "100000000000000000000000",
3994 => "100000000000000000000010",
3995 => "100000000000000000000000",
3996 => "100000000000000000000000",
3997 => "100000000000000000000000",
3998 => "100000000000000000000010",
3999 => "100000000000000000000000",
4000 => "100000000000000000000000",
4001 => "100000000000000000000000",
4002 => "100000000000000000000010",
4003 => "100000000000000000000010",
4004 => "100000000000000000000000",
4005 => "100000000000000000000000",
4006 => "100000000000000000000010",
4007 => "100000000000000000000000",
4008 => "100000000000000000000000",
4009 => "011111111111111111111111",
4010 => "011111111111111111111111",
4011 => "011111111111111111111110",
4012 => "011111111111111111111111",
4013 => "011111111111111111111111",
4014 => "011111111111111111111111",
4015 => "011111111111111111111100",
4016 => "011111111111111111111110",
4017 => "011111111111111111111111",
4018 => "011111111111111111111111",
4019 => "011111111111111111111101",
4020 => "011111111111111111111110",
4021 => "011111111111111111111111",
4022 => "011111111111111111111111",
4023 => "011111111111111111111110",
4024 => "011111111111111111111111",
4025 => "011111111111111111111111",
4026 => "011111111111111111111111",
4027 => "011111111111111111111110",
4028 => "011111111111111111111111",
4029 => "011111111111111111111111",
4030 => "011111111111111111111111",
4031 => "011111111111111111111111",
4032 => "011111111111111111111111",
4033 => "011111111111111111111110",
4034 => "011111111111111111111111",
4035 => "011111111111111111111111",
4036 => "011111111111111111111110",
4037 => "011111111111111111111111",
4038 => "011111111111111111111111",
4039 => "011111111111111111111111",
4040 => "011111111111111111111111",
4041 => "011111111111111111111111",
4042 => "011111111111111111111111",
4043 => "011111111111111111111110",
4044 => "011111111111111111111111",
4045 => "011111111111111111111111",
4046 => "011111111111111111111111",
4047 => "011111111111111111111111",
4048 => "011111111111111111111101",
4049 => "011111111111111111111111",
4050 => "011111111111111111111111",
4051 => "011111111111111111111111",
4052 => "011111111111111111111110",
4053 => "011111111111111111111110",
4054 => "011111111111111111111111",
4055 => "011111111111111111111111",
4056 => "011111111111111111111111",
4057 => "011111111111111111111100",
4058 => "011111111111111111111110",
4059 => "011111111111111111111111",
4060 => "011111111111111111111111",
4061 => "011111111111111111111011",
4062 => "011111111111111111111111",
4063 => "011111111111111111111111",
4064 => "011111111111111111111110",
4065 => "011111111111111111111111",
4066 => "011111111111111111111111",
4067 => "011111111111111111111110",
4068 => "011111111111111111111100",
4069 => "011111111111111111111111",
4070 => "011111111111111111111111",
4071 => "011111111111111111111100",
4072 => "011111111111111111111110",
4073 => "011111111111111111111111",
4074 => "011111111111111111111111",
4075 => "011111111111111111111111",
4076 => "011111111111111111111111",
4077 => "011111111111111111111111",
4078 => "011111111111111111111111",
4079 => "011111111111111111111110",
4080 => "011111111111111111111111",
4081 => "011111111111111111111111",
4082 => "011111111111111111111111",
4083 => "011111111111111111111101",
4084 => "011111111111111111111111",
4085 => "011111111111111111111111",
4086 => "011111111111111111111111",
4087 => "011111111111111111111111",
4088 => "011111111111111111111111",
4089 => "011111111111111111111111",
4090 => "011111111111111111111111",
4091 => "011111111111111111111111",
4092 => "011111111111111111111111",
4093 => "011111111111111111111111",
4094 => "011111111111111111111110",
4095 => "011111111111111111111111",
4096 => "011111111111111111111111",
4097 => "011111111111111111111111",
4098 => "011111111111111111111110",
4099 => "011111111111111111111111",
4100 => "011111111111111111111111",
4101 => "011111111111111111111111",
4102 => "011111111111111111111111",
4103 => "011111111111111111111111",
4104 => "011111111111111111111110",
4105 => "011111111111111111111111",
4106 => "011111111111111111111111",
4107 => "011111111111111111111111",
4108 => "011111111111111111111101",
4109 => "100000000000000000000010",
4110 => "100000000000000000000010",
4111 => "100000000000000000000000",
4112 => "100000000000000000000000",
4113 => "100000000000000000000001",
4114 => "100000000000000000000000",
4115 => "100000000000000000000000",
4116 => "100000000000000000000010",
4117 => "100000000000000000000000",
4118 => "100000000000000000000000",
4119 => "100000000000000000000010",
4120 => "100000000000000000000000",
4121 => "100000000000000000000000",
4122 => "100000000000000000000001",
4123 => "100000000000000000000011",
4124 => "100000000000000000000000",
4125 => "100000000000000000000000",
4126 => "100000000000000000000000",
4127 => "100000000000000000000010",
4128 => "100000000000000000000000",
4129 => "100000000000000000000000",
4130 => "100000000000000000000000",
4131 => "100000000000000000000010",
4132 => "100000000000000000000000",
4133 => "100000000000000000000000",
4134 => "100000000000000000000000",
4135 => "100000000000000000000011",
4136 => "100000000000000000000001",
4137 => "100000000000000000000000",
4138 => "100000000000000000000000",
4139 => "100000000000000000000100",
4140 => "100000000000000000000011",
4141 => "100000000000000000000000",
4142 => "100000000000000000000000",
4143 => "100000000000000000000100",
4144 => "100000000000000000000010",
4145 => "100000000000000000000000",
4146 => "100000000000000000000000",
4147 => "100000000000000000000011",
4148 => "100000000000000000000000",
4149 => "100000000000000000000000",
4150 => "100000000000000000000000",
4151 => "100000000000000000000000",
4152 => "100000000000000000000000",
4153 => "100000000000000000000010",
4154 => "100000000000000000000000",
4155 => "100000000000000000000000",
4156 => "100000000000000000000000",
4157 => "100000000000000000000010",
4158 => "100000000000000000000000",
4159 => "100000000000000000000000",
4160 => "100000000000000000000000",
4161 => "100000000000000000000000",
4162 => "100000000000000000000000",
4163 => "100000000000000000000000",
4164 => "100000000000000000000001",
4165 => "100000000000000000000000",
4166 => "100000000000000000000000",
4167 => "100000000000000000000000",
4168 => "100000000000000000000000",
4169 => "100000000000000000000000",
4170 => "100000000000000000000000",
4171 => "100000000000000000000001",
4172 => "100000000000000000000001",
4173 => "100000000000000000000000",
4174 => "100000000000000000000000",
4175 => "100000000000000000000000",
4176 => "100000000000000000000001",
4177 => "100000000000000000000001",
4178 => "100000000000000000000000",
4179 => "100000000000000000000000",
4180 => "100000000000000000000001",
4181 => "100000000000000000000000",
4182 => "100000000000000000000000",
4183 => "100000000000000000000000",
4184 => "100000000000000000000001",
4185 => "100000000000000000000000",
4186 => "100000000000000000000000",
4187 => "100000000000000000000000",
4188 => "100000000000000000000000",
4189 => "100000000000000000000000",
4190 => "100000000000000000000000",
4191 => "100000000000000000000001",
4192 => "100000000000000000000000",
4193 => "100000000000000000000000",
4194 => "100000000000000000000000",
4195 => "100000000000000000000000",
4196 => "100000000000000000000000",
4197 => "100000000000000000000010",
4198 => "100000000000000000000000",
4199 => "100000000000000000000000",
4200 => "100000000000000000000000",
4201 => "100000000000000000000100",
4202 => "100000000000000000000000",
4203 => "100000000000000000000000",
4204 => "100000000000000000000000",
4205 => "100000000000000000000100",
4206 => "100000000000000000000000",
4207 => "100000000000000000000000",
4208 => "100000000000000000000000",
4209 => "011111111111111111111111",
4210 => "011111111111111111111111",
4211 => "011111111111111111111110",
4212 => "011111111111111111111111",
4213 => "011111111111111111111111",
4214 => "011111111111111111111111",
4215 => "011111111111111111111110",
4216 => "011111111111111111111110",
4217 => "011111111111111111111111",
4218 => "011111111111111111111111",
4219 => "011111111111111111111110",
4220 => "011111111111111111111110",
4221 => "011111111111111111111111",
4222 => "011111111111111111111111",
4223 => "011111111111111111111111",
4224 => "011111111111111111111111",
4225 => "011111111111111111111100",
4226 => "011111111111111111111111",
4227 => "011111111111111111111111",
4228 => "011111111111111111111111",
4229 => "011111111111111111111100",
4230 => "011111111111111111111111",
4231 => "011111111111111111111111",
4232 => "011111111111111111111111",
4233 => "011111111111111111111110",
4234 => "011111111111111111111111",
4235 => "011111111111111111111111",
4236 => "011111111111111111111111",
4237 => "011111111111111111111111",
4238 => "011111111111111111111111",
4239 => "011111111111111111111111",
4240 => "011111111111111111111111",
4241 => "011111111111111111111111",
4242 => "011111111111111111111111",
4243 => "011111111111111111111111",
4244 => "011111111111111111111111",
4245 => "011111111111111111111101",
4246 => "011111111111111111111111",
4247 => "011111111111111111111111",
4248 => "011111111111111111111111",
4249 => "011111111111111111111110",
4250 => "011111111111111111111111",
4251 => "011111111111111111111111",
4252 => "011111111111111111111111",
4253 => "011111111111111111111111",
4254 => "011111111111111111111111",
4255 => "011111111111111111111111",
4256 => "011111111111111111111111",
4257 => "011111111111111111111111",
4258 => "011111111111111111111111",
4259 => "011111111111111111111111",
4260 => "011111111111111111111111",
4261 => "011111111111111111111110",
4262 => "011111111111111111111111",
4263 => "011111111111111111111111",
4264 => "011111111111111111111111",
4265 => "011111111111111111111111",
4266 => "011111111111111111111111",
4267 => "011111111111111111111111",
4268 => "011111111111111111111111",
4269 => "011111111111111111111111",
4270 => "011111111111111111111111",
4271 => "011111111111111111111110",
4272 => "011111111111111111111111",
4273 => "011111111111111111111111",
4274 => "011111111111111111111111",
4275 => "011111111111111111111110",
4276 => "011111111111111111111111",
4277 => "011111111111111111111111",
4278 => "011111111111111111111111",
4279 => "011111111111111111111111",
4280 => "011111111111111111111110",
4281 => "011111111111111111111111",
4282 => "011111111111111111111111",
4283 => "011111111111111111111111",
4284 => "011111111111111111111110",
4285 => "011111111111111111111111",
4286 => "011111111111111111111111",
4287 => "011111111111111111111111",
4288 => "011111111111111111111111",
4289 => "011111111111111111111111",
4290 => "011111111111111111111110",
4291 => "011111111111111111111111",
4292 => "011111111111111111111111",
4293 => "011111111111111111111111",
4294 => "011111111111111111111101",
4295 => "011111111111111111111111",
4296 => "011111111111111111111111",
4297 => "011111111111111111111110",
4298 => "011111111111111111111110",
4299 => "011111111111111111111111",
4300 => "011111111111111111111111",
4301 => "011111111111111111111101",
4302 => "011111111111111111111111",
4303 => "011111111111111111111111",
4304 => "011111111111111111111111",
4305 => "011111111111111111111110",
4306 => "011111111111111111111111",
4307 => "011111111111111111111111",
4308 => "011111111111111111111111",
4309 => "100000000000000000000000",
4310 => "100000000000000000000000",
4311 => "100000000000000000000001",
4312 => "100000000000000000000000",
4313 => "100000000000000000000000",
4314 => "100000000000000000000000",
4315 => "100000000000000000000010",
4316 => "100000000000000000000000",
4317 => "100000000000000000000000",
4318 => "100000000000000000000000",
4319 => "100000000000000000000010",
4320 => "100000000000000000000000",
4321 => "100000000000000000000000",
4322 => "100000000000000000000010",
4323 => "100000000000000000000000",
4324 => "100000000000000000000000",
4325 => "100000000000000000000010",
4326 => "100000000000000000000010",
4327 => "100000000000000000000000",
4328 => "100000000000000000000000",
4329 => "100000000000000000000011",
4330 => "100000000000000000000000",
4331 => "100000000000000000000000",
4332 => "100000000000000000000000",
4333 => "100000000000000000000001",
4334 => "100000000000000000000001",
4335 => "100000000000000000000000",
4336 => "100000000000000000000000",
4337 => "100000000000000000000000",
4338 => "100000000000000000000000",
4339 => "100000000000000000000000",
4340 => "100000000000000000000000",
4341 => "100000000000000000000000",
4342 => "100000000000000000000000",
4343 => "100000000000000000000000",
4344 => "100000000000000000000000",
4345 => "100000000000000000000000",
4346 => "100000000000000000000010",
4347 => "100000000000000000000000",
4348 => "100000000000000000000000",
4349 => "100000000000000000000000",
4350 => "100000000000000000000100",
4351 => "100000000000000000000001",
4352 => "100000000000000000000000",
4353 => "100000000000000000000000",
4354 => "100000000000000000000010",
4355 => "100000000000000000000010",
4356 => "100000000000000000000000",
4357 => "100000000000000000000000",
4358 => "100000000000000000000000",
4359 => "100000000000000000000010",
4360 => "100000000000000000000000",
4361 => "100000000000000000000000",
4362 => "100000000000000000000010",
4363 => "100000000000000000000010",
4364 => "100000000000000000000000",
4365 => "100000000000000000000000",
4366 => "100000000000000000000110",
4367 => "100000000000000000000010",
4368 => "100000000000000000000000",
4369 => "100000000000000000000000",
4370 => "100000000000000000000110",
4371 => "100000000000000000000010",
4372 => "100000000000000000000000",
4373 => "100000000000000000000000",
4374 => "100000000000000000000011",
4375 => "100000000000000000000010",
4376 => "100000000000000000000000",
4377 => "100000000000000000000000",
4378 => "100000000000000000000001",
4379 => "100000000000000000000001",
4380 => "100000000000000000000000",
4381 => "100000000000000000000000",
4382 => "100000000000000000000000",
4383 => "100000000000000000000000",
4384 => "100000000000000000000000",
4385 => "100000000000000000000000",
4386 => "100000000000000000000000",
4387 => "100000000000000000000010",
4388 => "100000000000000000000000",
4389 => "100000000000000000000000",
4390 => "100000000000000000000001",
4391 => "100000000000000000000010",
4392 => "100000000000000000000000",
4393 => "100000000000000000000000",
4394 => "100000000000000000000000",
4395 => "100000000000000000000000",
4396 => "100000000000000000000010",
4397 => "100000000000000000000100",
4398 => "100000000000000000000000",
4399 => "100000000000000000000000",
4400 => "100000000000000000000100",
4401 => "100000000000000000000101",
4402 => "100000000000000000000000",
4403 => "100000000000000000000000",
4404 => "100000000000000000000010",
4405 => "100000000000000000000110",
4406 => "100000000000000000000000",
4407 => "100000000000000000000000",
4408 => "100000000000000000000010");
signal count : std_logic_vector(13 -1 downto 0) := (others => '0');
begin
	getRomData: process (count)
	begin
		case count is
		when "0000000000000" => data_out <= rom_array(0);
		when "0000000000001" => data_out <= rom_array(1);
		when "0000000000010" => data_out <= rom_array(2);
		when "0000000000011" => data_out <= rom_array(3);
		when "0000000000100" => data_out <= rom_array(4);
		when "0000000000101" => data_out <= rom_array(5);
		when "0000000000110" => data_out <= rom_array(6);
		when "0000000000111" => data_out <= rom_array(7);
		when "0000000001000" => data_out <= rom_array(8);
		when "0000000001001" => data_out <= rom_array(9);
		when "0000000001010" => data_out <= rom_array(10);
		when "0000000001011" => data_out <= rom_array(11);
		when "0000000001100" => data_out <= rom_array(12);
		when "0000000001101" => data_out <= rom_array(13);
		when "0000000001110" => data_out <= rom_array(14);
		when "0000000001111" => data_out <= rom_array(15);
		when "0000000010000" => data_out <= rom_array(16);
		when "0000000010001" => data_out <= rom_array(17);
		when "0000000010010" => data_out <= rom_array(18);
		when "0000000010011" => data_out <= rom_array(19);
		when "0000000010100" => data_out <= rom_array(20);
		when "0000000010101" => data_out <= rom_array(21);
		when "0000000010110" => data_out <= rom_array(22);
		when "0000000010111" => data_out <= rom_array(23);
		when "0000000011000" => data_out <= rom_array(24);
		when "0000000011001" => data_out <= rom_array(25);
		when "0000000011010" => data_out <= rom_array(26);
		when "0000000011011" => data_out <= rom_array(27);
		when "0000000011100" => data_out <= rom_array(28);
		when "0000000011101" => data_out <= rom_array(29);
		when "0000000011110" => data_out <= rom_array(30);
		when "0000000011111" => data_out <= rom_array(31);
		when "0000000100000" => data_out <= rom_array(32);
		when "0000000100001" => data_out <= rom_array(33);
		when "0000000100010" => data_out <= rom_array(34);
		when "0000000100011" => data_out <= rom_array(35);
		when "0000000100100" => data_out <= rom_array(36);
		when "0000000100101" => data_out <= rom_array(37);
		when "0000000100110" => data_out <= rom_array(38);
		when "0000000100111" => data_out <= rom_array(39);
		when "0000000101000" => data_out <= rom_array(40);
		when "0000000101001" => data_out <= rom_array(41);
		when "0000000101010" => data_out <= rom_array(42);
		when "0000000101011" => data_out <= rom_array(43);
		when "0000000101100" => data_out <= rom_array(44);
		when "0000000101101" => data_out <= rom_array(45);
		when "0000000101110" => data_out <= rom_array(46);
		when "0000000101111" => data_out <= rom_array(47);
		when "0000000110000" => data_out <= rom_array(48);
		when "0000000110001" => data_out <= rom_array(49);
		when "0000000110010" => data_out <= rom_array(50);
		when "0000000110011" => data_out <= rom_array(51);
		when "0000000110100" => data_out <= rom_array(52);
		when "0000000110101" => data_out <= rom_array(53);
		when "0000000110110" => data_out <= rom_array(54);
		when "0000000110111" => data_out <= rom_array(55);
		when "0000000111000" => data_out <= rom_array(56);
		when "0000000111001" => data_out <= rom_array(57);
		when "0000000111010" => data_out <= rom_array(58);
		when "0000000111011" => data_out <= rom_array(59);
		when "0000000111100" => data_out <= rom_array(60);
		when "0000000111101" => data_out <= rom_array(61);
		when "0000000111110" => data_out <= rom_array(62);
		when "0000000111111" => data_out <= rom_array(63);
		when "0000001000000" => data_out <= rom_array(64);
		when "0000001000001" => data_out <= rom_array(65);
		when "0000001000010" => data_out <= rom_array(66);
		when "0000001000011" => data_out <= rom_array(67);
		when "0000001000100" => data_out <= rom_array(68);
		when "0000001000101" => data_out <= rom_array(69);
		when "0000001000110" => data_out <= rom_array(70);
		when "0000001000111" => data_out <= rom_array(71);
		when "0000001001000" => data_out <= rom_array(72);
		when "0000001001001" => data_out <= rom_array(73);
		when "0000001001010" => data_out <= rom_array(74);
		when "0000001001011" => data_out <= rom_array(75);
		when "0000001001100" => data_out <= rom_array(76);
		when "0000001001101" => data_out <= rom_array(77);
		when "0000001001110" => data_out <= rom_array(78);
		when "0000001001111" => data_out <= rom_array(79);
		when "0000001010000" => data_out <= rom_array(80);
		when "0000001010001" => data_out <= rom_array(81);
		when "0000001010010" => data_out <= rom_array(82);
		when "0000001010011" => data_out <= rom_array(83);
		when "0000001010100" => data_out <= rom_array(84);
		when "0000001010101" => data_out <= rom_array(85);
		when "0000001010110" => data_out <= rom_array(86);
		when "0000001010111" => data_out <= rom_array(87);
		when "0000001011000" => data_out <= rom_array(88);
		when "0000001011001" => data_out <= rom_array(89);
		when "0000001011010" => data_out <= rom_array(90);
		when "0000001011011" => data_out <= rom_array(91);
		when "0000001011100" => data_out <= rom_array(92);
		when "0000001011101" => data_out <= rom_array(93);
		when "0000001011110" => data_out <= rom_array(94);
		when "0000001011111" => data_out <= rom_array(95);
		when "0000001100000" => data_out <= rom_array(96);
		when "0000001100001" => data_out <= rom_array(97);
		when "0000001100010" => data_out <= rom_array(98);
		when "0000001100011" => data_out <= rom_array(99);
		when "0000001100100" => data_out <= rom_array(100);
		when "0000001100101" => data_out <= rom_array(101);
		when "0000001100110" => data_out <= rom_array(102);
		when "0000001100111" => data_out <= rom_array(103);
		when "0000001101000" => data_out <= rom_array(104);
		when "0000001101001" => data_out <= rom_array(105);
		when "0000001101010" => data_out <= rom_array(106);
		when "0000001101011" => data_out <= rom_array(107);
		when "0000001101100" => data_out <= rom_array(108);
		when "0000001101101" => data_out <= rom_array(109);
		when "0000001101110" => data_out <= rom_array(110);
		when "0000001101111" => data_out <= rom_array(111);
		when "0000001110000" => data_out <= rom_array(112);
		when "0000001110001" => data_out <= rom_array(113);
		when "0000001110010" => data_out <= rom_array(114);
		when "0000001110011" => data_out <= rom_array(115);
		when "0000001110100" => data_out <= rom_array(116);
		when "0000001110101" => data_out <= rom_array(117);
		when "0000001110110" => data_out <= rom_array(118);
		when "0000001110111" => data_out <= rom_array(119);
		when "0000001111000" => data_out <= rom_array(120);
		when "0000001111001" => data_out <= rom_array(121);
		when "0000001111010" => data_out <= rom_array(122);
		when "0000001111011" => data_out <= rom_array(123);
		when "0000001111100" => data_out <= rom_array(124);
		when "0000001111101" => data_out <= rom_array(125);
		when "0000001111110" => data_out <= rom_array(126);
		when "0000001111111" => data_out <= rom_array(127);
		when "0000010000000" => data_out <= rom_array(128);
		when "0000010000001" => data_out <= rom_array(129);
		when "0000010000010" => data_out <= rom_array(130);
		when "0000010000011" => data_out <= rom_array(131);
		when "0000010000100" => data_out <= rom_array(132);
		when "0000010000101" => data_out <= rom_array(133);
		when "0000010000110" => data_out <= rom_array(134);
		when "0000010000111" => data_out <= rom_array(135);
		when "0000010001000" => data_out <= rom_array(136);
		when "0000010001001" => data_out <= rom_array(137);
		when "0000010001010" => data_out <= rom_array(138);
		when "0000010001011" => data_out <= rom_array(139);
		when "0000010001100" => data_out <= rom_array(140);
		when "0000010001101" => data_out <= rom_array(141);
		when "0000010001110" => data_out <= rom_array(142);
		when "0000010001111" => data_out <= rom_array(143);
		when "0000010010000" => data_out <= rom_array(144);
		when "0000010010001" => data_out <= rom_array(145);
		when "0000010010010" => data_out <= rom_array(146);
		when "0000010010011" => data_out <= rom_array(147);
		when "0000010010100" => data_out <= rom_array(148);
		when "0000010010101" => data_out <= rom_array(149);
		when "0000010010110" => data_out <= rom_array(150);
		when "0000010010111" => data_out <= rom_array(151);
		when "0000010011000" => data_out <= rom_array(152);
		when "0000010011001" => data_out <= rom_array(153);
		when "0000010011010" => data_out <= rom_array(154);
		when "0000010011011" => data_out <= rom_array(155);
		when "0000010011100" => data_out <= rom_array(156);
		when "0000010011101" => data_out <= rom_array(157);
		when "0000010011110" => data_out <= rom_array(158);
		when "0000010011111" => data_out <= rom_array(159);
		when "0000010100000" => data_out <= rom_array(160);
		when "0000010100001" => data_out <= rom_array(161);
		when "0000010100010" => data_out <= rom_array(162);
		when "0000010100011" => data_out <= rom_array(163);
		when "0000010100100" => data_out <= rom_array(164);
		when "0000010100101" => data_out <= rom_array(165);
		when "0000010100110" => data_out <= rom_array(166);
		when "0000010100111" => data_out <= rom_array(167);
		when "0000010101000" => data_out <= rom_array(168);
		when "0000010101001" => data_out <= rom_array(169);
		when "0000010101010" => data_out <= rom_array(170);
		when "0000010101011" => data_out <= rom_array(171);
		when "0000010101100" => data_out <= rom_array(172);
		when "0000010101101" => data_out <= rom_array(173);
		when "0000010101110" => data_out <= rom_array(174);
		when "0000010101111" => data_out <= rom_array(175);
		when "0000010110000" => data_out <= rom_array(176);
		when "0000010110001" => data_out <= rom_array(177);
		when "0000010110010" => data_out <= rom_array(178);
		when "0000010110011" => data_out <= rom_array(179);
		when "0000010110100" => data_out <= rom_array(180);
		when "0000010110101" => data_out <= rom_array(181);
		when "0000010110110" => data_out <= rom_array(182);
		when "0000010110111" => data_out <= rom_array(183);
		when "0000010111000" => data_out <= rom_array(184);
		when "0000010111001" => data_out <= rom_array(185);
		when "0000010111010" => data_out <= rom_array(186);
		when "0000010111011" => data_out <= rom_array(187);
		when "0000010111100" => data_out <= rom_array(188);
		when "0000010111101" => data_out <= rom_array(189);
		when "0000010111110" => data_out <= rom_array(190);
		when "0000010111111" => data_out <= rom_array(191);
		when "0000011000000" => data_out <= rom_array(192);
		when "0000011000001" => data_out <= rom_array(193);
		when "0000011000010" => data_out <= rom_array(194);
		when "0000011000011" => data_out <= rom_array(195);
		when "0000011000100" => data_out <= rom_array(196);
		when "0000011000101" => data_out <= rom_array(197);
		when "0000011000110" => data_out <= rom_array(198);
		when "0000011000111" => data_out <= rom_array(199);
		when "0000011001000" => data_out <= rom_array(200);
		when "0000011001001" => data_out <= rom_array(201);
		when "0000011001010" => data_out <= rom_array(202);
		when "0000011001011" => data_out <= rom_array(203);
		when "0000011001100" => data_out <= rom_array(204);
		when "0000011001101" => data_out <= rom_array(205);
		when "0000011001110" => data_out <= rom_array(206);
		when "0000011001111" => data_out <= rom_array(207);
		when "0000011010000" => data_out <= rom_array(208);
		when "0000011010001" => data_out <= rom_array(209);
		when "0000011010010" => data_out <= rom_array(210);
		when "0000011010011" => data_out <= rom_array(211);
		when "0000011010100" => data_out <= rom_array(212);
		when "0000011010101" => data_out <= rom_array(213);
		when "0000011010110" => data_out <= rom_array(214);
		when "0000011010111" => data_out <= rom_array(215);
		when "0000011011000" => data_out <= rom_array(216);
		when "0000011011001" => data_out <= rom_array(217);
		when "0000011011010" => data_out <= rom_array(218);
		when "0000011011011" => data_out <= rom_array(219);
		when "0000011011100" => data_out <= rom_array(220);
		when "0000011011101" => data_out <= rom_array(221);
		when "0000011011110" => data_out <= rom_array(222);
		when "0000011011111" => data_out <= rom_array(223);
		when "0000011100000" => data_out <= rom_array(224);
		when "0000011100001" => data_out <= rom_array(225);
		when "0000011100010" => data_out <= rom_array(226);
		when "0000011100011" => data_out <= rom_array(227);
		when "0000011100100" => data_out <= rom_array(228);
		when "0000011100101" => data_out <= rom_array(229);
		when "0000011100110" => data_out <= rom_array(230);
		when "0000011100111" => data_out <= rom_array(231);
		when "0000011101000" => data_out <= rom_array(232);
		when "0000011101001" => data_out <= rom_array(233);
		when "0000011101010" => data_out <= rom_array(234);
		when "0000011101011" => data_out <= rom_array(235);
		when "0000011101100" => data_out <= rom_array(236);
		when "0000011101101" => data_out <= rom_array(237);
		when "0000011101110" => data_out <= rom_array(238);
		when "0000011101111" => data_out <= rom_array(239);
		when "0000011110000" => data_out <= rom_array(240);
		when "0000011110001" => data_out <= rom_array(241);
		when "0000011110010" => data_out <= rom_array(242);
		when "0000011110011" => data_out <= rom_array(243);
		when "0000011110100" => data_out <= rom_array(244);
		when "0000011110101" => data_out <= rom_array(245);
		when "0000011110110" => data_out <= rom_array(246);
		when "0000011110111" => data_out <= rom_array(247);
		when "0000011111000" => data_out <= rom_array(248);
		when "0000011111001" => data_out <= rom_array(249);
		when "0000011111010" => data_out <= rom_array(250);
		when "0000011111011" => data_out <= rom_array(251);
		when "0000011111100" => data_out <= rom_array(252);
		when "0000011111101" => data_out <= rom_array(253);
		when "0000011111110" => data_out <= rom_array(254);
		when "0000011111111" => data_out <= rom_array(255);
		when "0000100000000" => data_out <= rom_array(256);
		when "0000100000001" => data_out <= rom_array(257);
		when "0000100000010" => data_out <= rom_array(258);
		when "0000100000011" => data_out <= rom_array(259);
		when "0000100000100" => data_out <= rom_array(260);
		when "0000100000101" => data_out <= rom_array(261);
		when "0000100000110" => data_out <= rom_array(262);
		when "0000100000111" => data_out <= rom_array(263);
		when "0000100001000" => data_out <= rom_array(264);
		when "0000100001001" => data_out <= rom_array(265);
		when "0000100001010" => data_out <= rom_array(266);
		when "0000100001011" => data_out <= rom_array(267);
		when "0000100001100" => data_out <= rom_array(268);
		when "0000100001101" => data_out <= rom_array(269);
		when "0000100001110" => data_out <= rom_array(270);
		when "0000100001111" => data_out <= rom_array(271);
		when "0000100010000" => data_out <= rom_array(272);
		when "0000100010001" => data_out <= rom_array(273);
		when "0000100010010" => data_out <= rom_array(274);
		when "0000100010011" => data_out <= rom_array(275);
		when "0000100010100" => data_out <= rom_array(276);
		when "0000100010101" => data_out <= rom_array(277);
		when "0000100010110" => data_out <= rom_array(278);
		when "0000100010111" => data_out <= rom_array(279);
		when "0000100011000" => data_out <= rom_array(280);
		when "0000100011001" => data_out <= rom_array(281);
		when "0000100011010" => data_out <= rom_array(282);
		when "0000100011011" => data_out <= rom_array(283);
		when "0000100011100" => data_out <= rom_array(284);
		when "0000100011101" => data_out <= rom_array(285);
		when "0000100011110" => data_out <= rom_array(286);
		when "0000100011111" => data_out <= rom_array(287);
		when "0000100100000" => data_out <= rom_array(288);
		when "0000100100001" => data_out <= rom_array(289);
		when "0000100100010" => data_out <= rom_array(290);
		when "0000100100011" => data_out <= rom_array(291);
		when "0000100100100" => data_out <= rom_array(292);
		when "0000100100101" => data_out <= rom_array(293);
		when "0000100100110" => data_out <= rom_array(294);
		when "0000100100111" => data_out <= rom_array(295);
		when "0000100101000" => data_out <= rom_array(296);
		when "0000100101001" => data_out <= rom_array(297);
		when "0000100101010" => data_out <= rom_array(298);
		when "0000100101011" => data_out <= rom_array(299);
		when "0000100101100" => data_out <= rom_array(300);
		when "0000100101101" => data_out <= rom_array(301);
		when "0000100101110" => data_out <= rom_array(302);
		when "0000100101111" => data_out <= rom_array(303);
		when "0000100110000" => data_out <= rom_array(304);
		when "0000100110001" => data_out <= rom_array(305);
		when "0000100110010" => data_out <= rom_array(306);
		when "0000100110011" => data_out <= rom_array(307);
		when "0000100110100" => data_out <= rom_array(308);
		when "0000100110101" => data_out <= rom_array(309);
		when "0000100110110" => data_out <= rom_array(310);
		when "0000100110111" => data_out <= rom_array(311);
		when "0000100111000" => data_out <= rom_array(312);
		when "0000100111001" => data_out <= rom_array(313);
		when "0000100111010" => data_out <= rom_array(314);
		when "0000100111011" => data_out <= rom_array(315);
		when "0000100111100" => data_out <= rom_array(316);
		when "0000100111101" => data_out <= rom_array(317);
		when "0000100111110" => data_out <= rom_array(318);
		when "0000100111111" => data_out <= rom_array(319);
		when "0000101000000" => data_out <= rom_array(320);
		when "0000101000001" => data_out <= rom_array(321);
		when "0000101000010" => data_out <= rom_array(322);
		when "0000101000011" => data_out <= rom_array(323);
		when "0000101000100" => data_out <= rom_array(324);
		when "0000101000101" => data_out <= rom_array(325);
		when "0000101000110" => data_out <= rom_array(326);
		when "0000101000111" => data_out <= rom_array(327);
		when "0000101001000" => data_out <= rom_array(328);
		when "0000101001001" => data_out <= rom_array(329);
		when "0000101001010" => data_out <= rom_array(330);
		when "0000101001011" => data_out <= rom_array(331);
		when "0000101001100" => data_out <= rom_array(332);
		when "0000101001101" => data_out <= rom_array(333);
		when "0000101001110" => data_out <= rom_array(334);
		when "0000101001111" => data_out <= rom_array(335);
		when "0000101010000" => data_out <= rom_array(336);
		when "0000101010001" => data_out <= rom_array(337);
		when "0000101010010" => data_out <= rom_array(338);
		when "0000101010011" => data_out <= rom_array(339);
		when "0000101010100" => data_out <= rom_array(340);
		when "0000101010101" => data_out <= rom_array(341);
		when "0000101010110" => data_out <= rom_array(342);
		when "0000101010111" => data_out <= rom_array(343);
		when "0000101011000" => data_out <= rom_array(344);
		when "0000101011001" => data_out <= rom_array(345);
		when "0000101011010" => data_out <= rom_array(346);
		when "0000101011011" => data_out <= rom_array(347);
		when "0000101011100" => data_out <= rom_array(348);
		when "0000101011101" => data_out <= rom_array(349);
		when "0000101011110" => data_out <= rom_array(350);
		when "0000101011111" => data_out <= rom_array(351);
		when "0000101100000" => data_out <= rom_array(352);
		when "0000101100001" => data_out <= rom_array(353);
		when "0000101100010" => data_out <= rom_array(354);
		when "0000101100011" => data_out <= rom_array(355);
		when "0000101100100" => data_out <= rom_array(356);
		when "0000101100101" => data_out <= rom_array(357);
		when "0000101100110" => data_out <= rom_array(358);
		when "0000101100111" => data_out <= rom_array(359);
		when "0000101101000" => data_out <= rom_array(360);
		when "0000101101001" => data_out <= rom_array(361);
		when "0000101101010" => data_out <= rom_array(362);
		when "0000101101011" => data_out <= rom_array(363);
		when "0000101101100" => data_out <= rom_array(364);
		when "0000101101101" => data_out <= rom_array(365);
		when "0000101101110" => data_out <= rom_array(366);
		when "0000101101111" => data_out <= rom_array(367);
		when "0000101110000" => data_out <= rom_array(368);
		when "0000101110001" => data_out <= rom_array(369);
		when "0000101110010" => data_out <= rom_array(370);
		when "0000101110011" => data_out <= rom_array(371);
		when "0000101110100" => data_out <= rom_array(372);
		when "0000101110101" => data_out <= rom_array(373);
		when "0000101110110" => data_out <= rom_array(374);
		when "0000101110111" => data_out <= rom_array(375);
		when "0000101111000" => data_out <= rom_array(376);
		when "0000101111001" => data_out <= rom_array(377);
		when "0000101111010" => data_out <= rom_array(378);
		when "0000101111011" => data_out <= rom_array(379);
		when "0000101111100" => data_out <= rom_array(380);
		when "0000101111101" => data_out <= rom_array(381);
		when "0000101111110" => data_out <= rom_array(382);
		when "0000101111111" => data_out <= rom_array(383);
		when "0000110000000" => data_out <= rom_array(384);
		when "0000110000001" => data_out <= rom_array(385);
		when "0000110000010" => data_out <= rom_array(386);
		when "0000110000011" => data_out <= rom_array(387);
		when "0000110000100" => data_out <= rom_array(388);
		when "0000110000101" => data_out <= rom_array(389);
		when "0000110000110" => data_out <= rom_array(390);
		when "0000110000111" => data_out <= rom_array(391);
		when "0000110001000" => data_out <= rom_array(392);
		when "0000110001001" => data_out <= rom_array(393);
		when "0000110001010" => data_out <= rom_array(394);
		when "0000110001011" => data_out <= rom_array(395);
		when "0000110001100" => data_out <= rom_array(396);
		when "0000110001101" => data_out <= rom_array(397);
		when "0000110001110" => data_out <= rom_array(398);
		when "0000110001111" => data_out <= rom_array(399);
		when "0000110010000" => data_out <= rom_array(400);
		when "0000110010001" => data_out <= rom_array(401);
		when "0000110010010" => data_out <= rom_array(402);
		when "0000110010011" => data_out <= rom_array(403);
		when "0000110010100" => data_out <= rom_array(404);
		when "0000110010101" => data_out <= rom_array(405);
		when "0000110010110" => data_out <= rom_array(406);
		when "0000110010111" => data_out <= rom_array(407);
		when "0000110011000" => data_out <= rom_array(408);
		when "0000110011001" => data_out <= rom_array(409);
		when "0000110011010" => data_out <= rom_array(410);
		when "0000110011011" => data_out <= rom_array(411);
		when "0000110011100" => data_out <= rom_array(412);
		when "0000110011101" => data_out <= rom_array(413);
		when "0000110011110" => data_out <= rom_array(414);
		when "0000110011111" => data_out <= rom_array(415);
		when "0000110100000" => data_out <= rom_array(416);
		when "0000110100001" => data_out <= rom_array(417);
		when "0000110100010" => data_out <= rom_array(418);
		when "0000110100011" => data_out <= rom_array(419);
		when "0000110100100" => data_out <= rom_array(420);
		when "0000110100101" => data_out <= rom_array(421);
		when "0000110100110" => data_out <= rom_array(422);
		when "0000110100111" => data_out <= rom_array(423);
		when "0000110101000" => data_out <= rom_array(424);
		when "0000110101001" => data_out <= rom_array(425);
		when "0000110101010" => data_out <= rom_array(426);
		when "0000110101011" => data_out <= rom_array(427);
		when "0000110101100" => data_out <= rom_array(428);
		when "0000110101101" => data_out <= rom_array(429);
		when "0000110101110" => data_out <= rom_array(430);
		when "0000110101111" => data_out <= rom_array(431);
		when "0000110110000" => data_out <= rom_array(432);
		when "0000110110001" => data_out <= rom_array(433);
		when "0000110110010" => data_out <= rom_array(434);
		when "0000110110011" => data_out <= rom_array(435);
		when "0000110110100" => data_out <= rom_array(436);
		when "0000110110101" => data_out <= rom_array(437);
		when "0000110110110" => data_out <= rom_array(438);
		when "0000110110111" => data_out <= rom_array(439);
		when "0000110111000" => data_out <= rom_array(440);
		when "0000110111001" => data_out <= rom_array(441);
		when "0000110111010" => data_out <= rom_array(442);
		when "0000110111011" => data_out <= rom_array(443);
		when "0000110111100" => data_out <= rom_array(444);
		when "0000110111101" => data_out <= rom_array(445);
		when "0000110111110" => data_out <= rom_array(446);
		when "0000110111111" => data_out <= rom_array(447);
		when "0000111000000" => data_out <= rom_array(448);
		when "0000111000001" => data_out <= rom_array(449);
		when "0000111000010" => data_out <= rom_array(450);
		when "0000111000011" => data_out <= rom_array(451);
		when "0000111000100" => data_out <= rom_array(452);
		when "0000111000101" => data_out <= rom_array(453);
		when "0000111000110" => data_out <= rom_array(454);
		when "0000111000111" => data_out <= rom_array(455);
		when "0000111001000" => data_out <= rom_array(456);
		when "0000111001001" => data_out <= rom_array(457);
		when "0000111001010" => data_out <= rom_array(458);
		when "0000111001011" => data_out <= rom_array(459);
		when "0000111001100" => data_out <= rom_array(460);
		when "0000111001101" => data_out <= rom_array(461);
		when "0000111001110" => data_out <= rom_array(462);
		when "0000111001111" => data_out <= rom_array(463);
		when "0000111010000" => data_out <= rom_array(464);
		when "0000111010001" => data_out <= rom_array(465);
		when "0000111010010" => data_out <= rom_array(466);
		when "0000111010011" => data_out <= rom_array(467);
		when "0000111010100" => data_out <= rom_array(468);
		when "0000111010101" => data_out <= rom_array(469);
		when "0000111010110" => data_out <= rom_array(470);
		when "0000111010111" => data_out <= rom_array(471);
		when "0000111011000" => data_out <= rom_array(472);
		when "0000111011001" => data_out <= rom_array(473);
		when "0000111011010" => data_out <= rom_array(474);
		when "0000111011011" => data_out <= rom_array(475);
		when "0000111011100" => data_out <= rom_array(476);
		when "0000111011101" => data_out <= rom_array(477);
		when "0000111011110" => data_out <= rom_array(478);
		when "0000111011111" => data_out <= rom_array(479);
		when "0000111100000" => data_out <= rom_array(480);
		when "0000111100001" => data_out <= rom_array(481);
		when "0000111100010" => data_out <= rom_array(482);
		when "0000111100011" => data_out <= rom_array(483);
		when "0000111100100" => data_out <= rom_array(484);
		when "0000111100101" => data_out <= rom_array(485);
		when "0000111100110" => data_out <= rom_array(486);
		when "0000111100111" => data_out <= rom_array(487);
		when "0000111101000" => data_out <= rom_array(488);
		when "0000111101001" => data_out <= rom_array(489);
		when "0000111101010" => data_out <= rom_array(490);
		when "0000111101011" => data_out <= rom_array(491);
		when "0000111101100" => data_out <= rom_array(492);
		when "0000111101101" => data_out <= rom_array(493);
		when "0000111101110" => data_out <= rom_array(494);
		when "0000111101111" => data_out <= rom_array(495);
		when "0000111110000" => data_out <= rom_array(496);
		when "0000111110001" => data_out <= rom_array(497);
		when "0000111110010" => data_out <= rom_array(498);
		when "0000111110011" => data_out <= rom_array(499);
		when "0000111110100" => data_out <= rom_array(500);
		when "0000111110101" => data_out <= rom_array(501);
		when "0000111110110" => data_out <= rom_array(502);
		when "0000111110111" => data_out <= rom_array(503);
		when "0000111111000" => data_out <= rom_array(504);
		when "0000111111001" => data_out <= rom_array(505);
		when "0000111111010" => data_out <= rom_array(506);
		when "0000111111011" => data_out <= rom_array(507);
		when "0000111111100" => data_out <= rom_array(508);
		when "0000111111101" => data_out <= rom_array(509);
		when "0000111111110" => data_out <= rom_array(510);
		when "0000111111111" => data_out <= rom_array(511);
		when "0001000000000" => data_out <= rom_array(512);
		when "0001000000001" => data_out <= rom_array(513);
		when "0001000000010" => data_out <= rom_array(514);
		when "0001000000011" => data_out <= rom_array(515);
		when "0001000000100" => data_out <= rom_array(516);
		when "0001000000101" => data_out <= rom_array(517);
		when "0001000000110" => data_out <= rom_array(518);
		when "0001000000111" => data_out <= rom_array(519);
		when "0001000001000" => data_out <= rom_array(520);
		when "0001000001001" => data_out <= rom_array(521);
		when "0001000001010" => data_out <= rom_array(522);
		when "0001000001011" => data_out <= rom_array(523);
		when "0001000001100" => data_out <= rom_array(524);
		when "0001000001101" => data_out <= rom_array(525);
		when "0001000001110" => data_out <= rom_array(526);
		when "0001000001111" => data_out <= rom_array(527);
		when "0001000010000" => data_out <= rom_array(528);
		when "0001000010001" => data_out <= rom_array(529);
		when "0001000010010" => data_out <= rom_array(530);
		when "0001000010011" => data_out <= rom_array(531);
		when "0001000010100" => data_out <= rom_array(532);
		when "0001000010101" => data_out <= rom_array(533);
		when "0001000010110" => data_out <= rom_array(534);
		when "0001000010111" => data_out <= rom_array(535);
		when "0001000011000" => data_out <= rom_array(536);
		when "0001000011001" => data_out <= rom_array(537);
		when "0001000011010" => data_out <= rom_array(538);
		when "0001000011011" => data_out <= rom_array(539);
		when "0001000011100" => data_out <= rom_array(540);
		when "0001000011101" => data_out <= rom_array(541);
		when "0001000011110" => data_out <= rom_array(542);
		when "0001000011111" => data_out <= rom_array(543);
		when "0001000100000" => data_out <= rom_array(544);
		when "0001000100001" => data_out <= rom_array(545);
		when "0001000100010" => data_out <= rom_array(546);
		when "0001000100011" => data_out <= rom_array(547);
		when "0001000100100" => data_out <= rom_array(548);
		when "0001000100101" => data_out <= rom_array(549);
		when "0001000100110" => data_out <= rom_array(550);
		when "0001000100111" => data_out <= rom_array(551);
		when "0001000101000" => data_out <= rom_array(552);
		when "0001000101001" => data_out <= rom_array(553);
		when "0001000101010" => data_out <= rom_array(554);
		when "0001000101011" => data_out <= rom_array(555);
		when "0001000101100" => data_out <= rom_array(556);
		when "0001000101101" => data_out <= rom_array(557);
		when "0001000101110" => data_out <= rom_array(558);
		when "0001000101111" => data_out <= rom_array(559);
		when "0001000110000" => data_out <= rom_array(560);
		when "0001000110001" => data_out <= rom_array(561);
		when "0001000110010" => data_out <= rom_array(562);
		when "0001000110011" => data_out <= rom_array(563);
		when "0001000110100" => data_out <= rom_array(564);
		when "0001000110101" => data_out <= rom_array(565);
		when "0001000110110" => data_out <= rom_array(566);
		when "0001000110111" => data_out <= rom_array(567);
		when "0001000111000" => data_out <= rom_array(568);
		when "0001000111001" => data_out <= rom_array(569);
		when "0001000111010" => data_out <= rom_array(570);
		when "0001000111011" => data_out <= rom_array(571);
		when "0001000111100" => data_out <= rom_array(572);
		when "0001000111101" => data_out <= rom_array(573);
		when "0001000111110" => data_out <= rom_array(574);
		when "0001000111111" => data_out <= rom_array(575);
		when "0001001000000" => data_out <= rom_array(576);
		when "0001001000001" => data_out <= rom_array(577);
		when "0001001000010" => data_out <= rom_array(578);
		when "0001001000011" => data_out <= rom_array(579);
		when "0001001000100" => data_out <= rom_array(580);
		when "0001001000101" => data_out <= rom_array(581);
		when "0001001000110" => data_out <= rom_array(582);
		when "0001001000111" => data_out <= rom_array(583);
		when "0001001001000" => data_out <= rom_array(584);
		when "0001001001001" => data_out <= rom_array(585);
		when "0001001001010" => data_out <= rom_array(586);
		when "0001001001011" => data_out <= rom_array(587);
		when "0001001001100" => data_out <= rom_array(588);
		when "0001001001101" => data_out <= rom_array(589);
		when "0001001001110" => data_out <= rom_array(590);
		when "0001001001111" => data_out <= rom_array(591);
		when "0001001010000" => data_out <= rom_array(592);
		when "0001001010001" => data_out <= rom_array(593);
		when "0001001010010" => data_out <= rom_array(594);
		when "0001001010011" => data_out <= rom_array(595);
		when "0001001010100" => data_out <= rom_array(596);
		when "0001001010101" => data_out <= rom_array(597);
		when "0001001010110" => data_out <= rom_array(598);
		when "0001001010111" => data_out <= rom_array(599);
		when "0001001011000" => data_out <= rom_array(600);
		when "0001001011001" => data_out <= rom_array(601);
		when "0001001011010" => data_out <= rom_array(602);
		when "0001001011011" => data_out <= rom_array(603);
		when "0001001011100" => data_out <= rom_array(604);
		when "0001001011101" => data_out <= rom_array(605);
		when "0001001011110" => data_out <= rom_array(606);
		when "0001001011111" => data_out <= rom_array(607);
		when "0001001100000" => data_out <= rom_array(608);
		when "0001001100001" => data_out <= rom_array(609);
		when "0001001100010" => data_out <= rom_array(610);
		when "0001001100011" => data_out <= rom_array(611);
		when "0001001100100" => data_out <= rom_array(612);
		when "0001001100101" => data_out <= rom_array(613);
		when "0001001100110" => data_out <= rom_array(614);
		when "0001001100111" => data_out <= rom_array(615);
		when "0001001101000" => data_out <= rom_array(616);
		when "0001001101001" => data_out <= rom_array(617);
		when "0001001101010" => data_out <= rom_array(618);
		when "0001001101011" => data_out <= rom_array(619);
		when "0001001101100" => data_out <= rom_array(620);
		when "0001001101101" => data_out <= rom_array(621);
		when "0001001101110" => data_out <= rom_array(622);
		when "0001001101111" => data_out <= rom_array(623);
		when "0001001110000" => data_out <= rom_array(624);
		when "0001001110001" => data_out <= rom_array(625);
		when "0001001110010" => data_out <= rom_array(626);
		when "0001001110011" => data_out <= rom_array(627);
		when "0001001110100" => data_out <= rom_array(628);
		when "0001001110101" => data_out <= rom_array(629);
		when "0001001110110" => data_out <= rom_array(630);
		when "0001001110111" => data_out <= rom_array(631);
		when "0001001111000" => data_out <= rom_array(632);
		when "0001001111001" => data_out <= rom_array(633);
		when "0001001111010" => data_out <= rom_array(634);
		when "0001001111011" => data_out <= rom_array(635);
		when "0001001111100" => data_out <= rom_array(636);
		when "0001001111101" => data_out <= rom_array(637);
		when "0001001111110" => data_out <= rom_array(638);
		when "0001001111111" => data_out <= rom_array(639);
		when "0001010000000" => data_out <= rom_array(640);
		when "0001010000001" => data_out <= rom_array(641);
		when "0001010000010" => data_out <= rom_array(642);
		when "0001010000011" => data_out <= rom_array(643);
		when "0001010000100" => data_out <= rom_array(644);
		when "0001010000101" => data_out <= rom_array(645);
		when "0001010000110" => data_out <= rom_array(646);
		when "0001010000111" => data_out <= rom_array(647);
		when "0001010001000" => data_out <= rom_array(648);
		when "0001010001001" => data_out <= rom_array(649);
		when "0001010001010" => data_out <= rom_array(650);
		when "0001010001011" => data_out <= rom_array(651);
		when "0001010001100" => data_out <= rom_array(652);
		when "0001010001101" => data_out <= rom_array(653);
		when "0001010001110" => data_out <= rom_array(654);
		when "0001010001111" => data_out <= rom_array(655);
		when "0001010010000" => data_out <= rom_array(656);
		when "0001010010001" => data_out <= rom_array(657);
		when "0001010010010" => data_out <= rom_array(658);
		when "0001010010011" => data_out <= rom_array(659);
		when "0001010010100" => data_out <= rom_array(660);
		when "0001010010101" => data_out <= rom_array(661);
		when "0001010010110" => data_out <= rom_array(662);
		when "0001010010111" => data_out <= rom_array(663);
		when "0001010011000" => data_out <= rom_array(664);
		when "0001010011001" => data_out <= rom_array(665);
		when "0001010011010" => data_out <= rom_array(666);
		when "0001010011011" => data_out <= rom_array(667);
		when "0001010011100" => data_out <= rom_array(668);
		when "0001010011101" => data_out <= rom_array(669);
		when "0001010011110" => data_out <= rom_array(670);
		when "0001010011111" => data_out <= rom_array(671);
		when "0001010100000" => data_out <= rom_array(672);
		when "0001010100001" => data_out <= rom_array(673);
		when "0001010100010" => data_out <= rom_array(674);
		when "0001010100011" => data_out <= rom_array(675);
		when "0001010100100" => data_out <= rom_array(676);
		when "0001010100101" => data_out <= rom_array(677);
		when "0001010100110" => data_out <= rom_array(678);
		when "0001010100111" => data_out <= rom_array(679);
		when "0001010101000" => data_out <= rom_array(680);
		when "0001010101001" => data_out <= rom_array(681);
		when "0001010101010" => data_out <= rom_array(682);
		when "0001010101011" => data_out <= rom_array(683);
		when "0001010101100" => data_out <= rom_array(684);
		when "0001010101101" => data_out <= rom_array(685);
		when "0001010101110" => data_out <= rom_array(686);
		when "0001010101111" => data_out <= rom_array(687);
		when "0001010110000" => data_out <= rom_array(688);
		when "0001010110001" => data_out <= rom_array(689);
		when "0001010110010" => data_out <= rom_array(690);
		when "0001010110011" => data_out <= rom_array(691);
		when "0001010110100" => data_out <= rom_array(692);
		when "0001010110101" => data_out <= rom_array(693);
		when "0001010110110" => data_out <= rom_array(694);
		when "0001010110111" => data_out <= rom_array(695);
		when "0001010111000" => data_out <= rom_array(696);
		when "0001010111001" => data_out <= rom_array(697);
		when "0001010111010" => data_out <= rom_array(698);
		when "0001010111011" => data_out <= rom_array(699);
		when "0001010111100" => data_out <= rom_array(700);
		when "0001010111101" => data_out <= rom_array(701);
		when "0001010111110" => data_out <= rom_array(702);
		when "0001010111111" => data_out <= rom_array(703);
		when "0001011000000" => data_out <= rom_array(704);
		when "0001011000001" => data_out <= rom_array(705);
		when "0001011000010" => data_out <= rom_array(706);
		when "0001011000011" => data_out <= rom_array(707);
		when "0001011000100" => data_out <= rom_array(708);
		when "0001011000101" => data_out <= rom_array(709);
		when "0001011000110" => data_out <= rom_array(710);
		when "0001011000111" => data_out <= rom_array(711);
		when "0001011001000" => data_out <= rom_array(712);
		when "0001011001001" => data_out <= rom_array(713);
		when "0001011001010" => data_out <= rom_array(714);
		when "0001011001011" => data_out <= rom_array(715);
		when "0001011001100" => data_out <= rom_array(716);
		when "0001011001101" => data_out <= rom_array(717);
		when "0001011001110" => data_out <= rom_array(718);
		when "0001011001111" => data_out <= rom_array(719);
		when "0001011010000" => data_out <= rom_array(720);
		when "0001011010001" => data_out <= rom_array(721);
		when "0001011010010" => data_out <= rom_array(722);
		when "0001011010011" => data_out <= rom_array(723);
		when "0001011010100" => data_out <= rom_array(724);
		when "0001011010101" => data_out <= rom_array(725);
		when "0001011010110" => data_out <= rom_array(726);
		when "0001011010111" => data_out <= rom_array(727);
		when "0001011011000" => data_out <= rom_array(728);
		when "0001011011001" => data_out <= rom_array(729);
		when "0001011011010" => data_out <= rom_array(730);
		when "0001011011011" => data_out <= rom_array(731);
		when "0001011011100" => data_out <= rom_array(732);
		when "0001011011101" => data_out <= rom_array(733);
		when "0001011011110" => data_out <= rom_array(734);
		when "0001011011111" => data_out <= rom_array(735);
		when "0001011100000" => data_out <= rom_array(736);
		when "0001011100001" => data_out <= rom_array(737);
		when "0001011100010" => data_out <= rom_array(738);
		when "0001011100011" => data_out <= rom_array(739);
		when "0001011100100" => data_out <= rom_array(740);
		when "0001011100101" => data_out <= rom_array(741);
		when "0001011100110" => data_out <= rom_array(742);
		when "0001011100111" => data_out <= rom_array(743);
		when "0001011101000" => data_out <= rom_array(744);
		when "0001011101001" => data_out <= rom_array(745);
		when "0001011101010" => data_out <= rom_array(746);
		when "0001011101011" => data_out <= rom_array(747);
		when "0001011101100" => data_out <= rom_array(748);
		when "0001011101101" => data_out <= rom_array(749);
		when "0001011101110" => data_out <= rom_array(750);
		when "0001011101111" => data_out <= rom_array(751);
		when "0001011110000" => data_out <= rom_array(752);
		when "0001011110001" => data_out <= rom_array(753);
		when "0001011110010" => data_out <= rom_array(754);
		when "0001011110011" => data_out <= rom_array(755);
		when "0001011110100" => data_out <= rom_array(756);
		when "0001011110101" => data_out <= rom_array(757);
		when "0001011110110" => data_out <= rom_array(758);
		when "0001011110111" => data_out <= rom_array(759);
		when "0001011111000" => data_out <= rom_array(760);
		when "0001011111001" => data_out <= rom_array(761);
		when "0001011111010" => data_out <= rom_array(762);
		when "0001011111011" => data_out <= rom_array(763);
		when "0001011111100" => data_out <= rom_array(764);
		when "0001011111101" => data_out <= rom_array(765);
		when "0001011111110" => data_out <= rom_array(766);
		when "0001011111111" => data_out <= rom_array(767);
		when "0001100000000" => data_out <= rom_array(768);
		when "0001100000001" => data_out <= rom_array(769);
		when "0001100000010" => data_out <= rom_array(770);
		when "0001100000011" => data_out <= rom_array(771);
		when "0001100000100" => data_out <= rom_array(772);
		when "0001100000101" => data_out <= rom_array(773);
		when "0001100000110" => data_out <= rom_array(774);
		when "0001100000111" => data_out <= rom_array(775);
		when "0001100001000" => data_out <= rom_array(776);
		when "0001100001001" => data_out <= rom_array(777);
		when "0001100001010" => data_out <= rom_array(778);
		when "0001100001011" => data_out <= rom_array(779);
		when "0001100001100" => data_out <= rom_array(780);
		when "0001100001101" => data_out <= rom_array(781);
		when "0001100001110" => data_out <= rom_array(782);
		when "0001100001111" => data_out <= rom_array(783);
		when "0001100010000" => data_out <= rom_array(784);
		when "0001100010001" => data_out <= rom_array(785);
		when "0001100010010" => data_out <= rom_array(786);
		when "0001100010011" => data_out <= rom_array(787);
		when "0001100010100" => data_out <= rom_array(788);
		when "0001100010101" => data_out <= rom_array(789);
		when "0001100010110" => data_out <= rom_array(790);
		when "0001100010111" => data_out <= rom_array(791);
		when "0001100011000" => data_out <= rom_array(792);
		when "0001100011001" => data_out <= rom_array(793);
		when "0001100011010" => data_out <= rom_array(794);
		when "0001100011011" => data_out <= rom_array(795);
		when "0001100011100" => data_out <= rom_array(796);
		when "0001100011101" => data_out <= rom_array(797);
		when "0001100011110" => data_out <= rom_array(798);
		when "0001100011111" => data_out <= rom_array(799);
		when "0001100100000" => data_out <= rom_array(800);
		when "0001100100001" => data_out <= rom_array(801);
		when "0001100100010" => data_out <= rom_array(802);
		when "0001100100011" => data_out <= rom_array(803);
		when "0001100100100" => data_out <= rom_array(804);
		when "0001100100101" => data_out <= rom_array(805);
		when "0001100100110" => data_out <= rom_array(806);
		when "0001100100111" => data_out <= rom_array(807);
		when "0001100101000" => data_out <= rom_array(808);
		when "0001100101001" => data_out <= rom_array(809);
		when "0001100101010" => data_out <= rom_array(810);
		when "0001100101011" => data_out <= rom_array(811);
		when "0001100101100" => data_out <= rom_array(812);
		when "0001100101101" => data_out <= rom_array(813);
		when "0001100101110" => data_out <= rom_array(814);
		when "0001100101111" => data_out <= rom_array(815);
		when "0001100110000" => data_out <= rom_array(816);
		when "0001100110001" => data_out <= rom_array(817);
		when "0001100110010" => data_out <= rom_array(818);
		when "0001100110011" => data_out <= rom_array(819);
		when "0001100110100" => data_out <= rom_array(820);
		when "0001100110101" => data_out <= rom_array(821);
		when "0001100110110" => data_out <= rom_array(822);
		when "0001100110111" => data_out <= rom_array(823);
		when "0001100111000" => data_out <= rom_array(824);
		when "0001100111001" => data_out <= rom_array(825);
		when "0001100111010" => data_out <= rom_array(826);
		when "0001100111011" => data_out <= rom_array(827);
		when "0001100111100" => data_out <= rom_array(828);
		when "0001100111101" => data_out <= rom_array(829);
		when "0001100111110" => data_out <= rom_array(830);
		when "0001100111111" => data_out <= rom_array(831);
		when "0001101000000" => data_out <= rom_array(832);
		when "0001101000001" => data_out <= rom_array(833);
		when "0001101000010" => data_out <= rom_array(834);
		when "0001101000011" => data_out <= rom_array(835);
		when "0001101000100" => data_out <= rom_array(836);
		when "0001101000101" => data_out <= rom_array(837);
		when "0001101000110" => data_out <= rom_array(838);
		when "0001101000111" => data_out <= rom_array(839);
		when "0001101001000" => data_out <= rom_array(840);
		when "0001101001001" => data_out <= rom_array(841);
		when "0001101001010" => data_out <= rom_array(842);
		when "0001101001011" => data_out <= rom_array(843);
		when "0001101001100" => data_out <= rom_array(844);
		when "0001101001101" => data_out <= rom_array(845);
		when "0001101001110" => data_out <= rom_array(846);
		when "0001101001111" => data_out <= rom_array(847);
		when "0001101010000" => data_out <= rom_array(848);
		when "0001101010001" => data_out <= rom_array(849);
		when "0001101010010" => data_out <= rom_array(850);
		when "0001101010011" => data_out <= rom_array(851);
		when "0001101010100" => data_out <= rom_array(852);
		when "0001101010101" => data_out <= rom_array(853);
		when "0001101010110" => data_out <= rom_array(854);
		when "0001101010111" => data_out <= rom_array(855);
		when "0001101011000" => data_out <= rom_array(856);
		when "0001101011001" => data_out <= rom_array(857);
		when "0001101011010" => data_out <= rom_array(858);
		when "0001101011011" => data_out <= rom_array(859);
		when "0001101011100" => data_out <= rom_array(860);
		when "0001101011101" => data_out <= rom_array(861);
		when "0001101011110" => data_out <= rom_array(862);
		when "0001101011111" => data_out <= rom_array(863);
		when "0001101100000" => data_out <= rom_array(864);
		when "0001101100001" => data_out <= rom_array(865);
		when "0001101100010" => data_out <= rom_array(866);
		when "0001101100011" => data_out <= rom_array(867);
		when "0001101100100" => data_out <= rom_array(868);
		when "0001101100101" => data_out <= rom_array(869);
		when "0001101100110" => data_out <= rom_array(870);
		when "0001101100111" => data_out <= rom_array(871);
		when "0001101101000" => data_out <= rom_array(872);
		when "0001101101001" => data_out <= rom_array(873);
		when "0001101101010" => data_out <= rom_array(874);
		when "0001101101011" => data_out <= rom_array(875);
		when "0001101101100" => data_out <= rom_array(876);
		when "0001101101101" => data_out <= rom_array(877);
		when "0001101101110" => data_out <= rom_array(878);
		when "0001101101111" => data_out <= rom_array(879);
		when "0001101110000" => data_out <= rom_array(880);
		when "0001101110001" => data_out <= rom_array(881);
		when "0001101110010" => data_out <= rom_array(882);
		when "0001101110011" => data_out <= rom_array(883);
		when "0001101110100" => data_out <= rom_array(884);
		when "0001101110101" => data_out <= rom_array(885);
		when "0001101110110" => data_out <= rom_array(886);
		when "0001101110111" => data_out <= rom_array(887);
		when "0001101111000" => data_out <= rom_array(888);
		when "0001101111001" => data_out <= rom_array(889);
		when "0001101111010" => data_out <= rom_array(890);
		when "0001101111011" => data_out <= rom_array(891);
		when "0001101111100" => data_out <= rom_array(892);
		when "0001101111101" => data_out <= rom_array(893);
		when "0001101111110" => data_out <= rom_array(894);
		when "0001101111111" => data_out <= rom_array(895);
		when "0001110000000" => data_out <= rom_array(896);
		when "0001110000001" => data_out <= rom_array(897);
		when "0001110000010" => data_out <= rom_array(898);
		when "0001110000011" => data_out <= rom_array(899);
		when "0001110000100" => data_out <= rom_array(900);
		when "0001110000101" => data_out <= rom_array(901);
		when "0001110000110" => data_out <= rom_array(902);
		when "0001110000111" => data_out <= rom_array(903);
		when "0001110001000" => data_out <= rom_array(904);
		when "0001110001001" => data_out <= rom_array(905);
		when "0001110001010" => data_out <= rom_array(906);
		when "0001110001011" => data_out <= rom_array(907);
		when "0001110001100" => data_out <= rom_array(908);
		when "0001110001101" => data_out <= rom_array(909);
		when "0001110001110" => data_out <= rom_array(910);
		when "0001110001111" => data_out <= rom_array(911);
		when "0001110010000" => data_out <= rom_array(912);
		when "0001110010001" => data_out <= rom_array(913);
		when "0001110010010" => data_out <= rom_array(914);
		when "0001110010011" => data_out <= rom_array(915);
		when "0001110010100" => data_out <= rom_array(916);
		when "0001110010101" => data_out <= rom_array(917);
		when "0001110010110" => data_out <= rom_array(918);
		when "0001110010111" => data_out <= rom_array(919);
		when "0001110011000" => data_out <= rom_array(920);
		when "0001110011001" => data_out <= rom_array(921);
		when "0001110011010" => data_out <= rom_array(922);
		when "0001110011011" => data_out <= rom_array(923);
		when "0001110011100" => data_out <= rom_array(924);
		when "0001110011101" => data_out <= rom_array(925);
		when "0001110011110" => data_out <= rom_array(926);
		when "0001110011111" => data_out <= rom_array(927);
		when "0001110100000" => data_out <= rom_array(928);
		when "0001110100001" => data_out <= rom_array(929);
		when "0001110100010" => data_out <= rom_array(930);
		when "0001110100011" => data_out <= rom_array(931);
		when "0001110100100" => data_out <= rom_array(932);
		when "0001110100101" => data_out <= rom_array(933);
		when "0001110100110" => data_out <= rom_array(934);
		when "0001110100111" => data_out <= rom_array(935);
		when "0001110101000" => data_out <= rom_array(936);
		when "0001110101001" => data_out <= rom_array(937);
		when "0001110101010" => data_out <= rom_array(938);
		when "0001110101011" => data_out <= rom_array(939);
		when "0001110101100" => data_out <= rom_array(940);
		when "0001110101101" => data_out <= rom_array(941);
		when "0001110101110" => data_out <= rom_array(942);
		when "0001110101111" => data_out <= rom_array(943);
		when "0001110110000" => data_out <= rom_array(944);
		when "0001110110001" => data_out <= rom_array(945);
		when "0001110110010" => data_out <= rom_array(946);
		when "0001110110011" => data_out <= rom_array(947);
		when "0001110110100" => data_out <= rom_array(948);
		when "0001110110101" => data_out <= rom_array(949);
		when "0001110110110" => data_out <= rom_array(950);
		when "0001110110111" => data_out <= rom_array(951);
		when "0001110111000" => data_out <= rom_array(952);
		when "0001110111001" => data_out <= rom_array(953);
		when "0001110111010" => data_out <= rom_array(954);
		when "0001110111011" => data_out <= rom_array(955);
		when "0001110111100" => data_out <= rom_array(956);
		when "0001110111101" => data_out <= rom_array(957);
		when "0001110111110" => data_out <= rom_array(958);
		when "0001110111111" => data_out <= rom_array(959);
		when "0001111000000" => data_out <= rom_array(960);
		when "0001111000001" => data_out <= rom_array(961);
		when "0001111000010" => data_out <= rom_array(962);
		when "0001111000011" => data_out <= rom_array(963);
		when "0001111000100" => data_out <= rom_array(964);
		when "0001111000101" => data_out <= rom_array(965);
		when "0001111000110" => data_out <= rom_array(966);
		when "0001111000111" => data_out <= rom_array(967);
		when "0001111001000" => data_out <= rom_array(968);
		when "0001111001001" => data_out <= rom_array(969);
		when "0001111001010" => data_out <= rom_array(970);
		when "0001111001011" => data_out <= rom_array(971);
		when "0001111001100" => data_out <= rom_array(972);
		when "0001111001101" => data_out <= rom_array(973);
		when "0001111001110" => data_out <= rom_array(974);
		when "0001111001111" => data_out <= rom_array(975);
		when "0001111010000" => data_out <= rom_array(976);
		when "0001111010001" => data_out <= rom_array(977);
		when "0001111010010" => data_out <= rom_array(978);
		when "0001111010011" => data_out <= rom_array(979);
		when "0001111010100" => data_out <= rom_array(980);
		when "0001111010101" => data_out <= rom_array(981);
		when "0001111010110" => data_out <= rom_array(982);
		when "0001111010111" => data_out <= rom_array(983);
		when "0001111011000" => data_out <= rom_array(984);
		when "0001111011001" => data_out <= rom_array(985);
		when "0001111011010" => data_out <= rom_array(986);
		when "0001111011011" => data_out <= rom_array(987);
		when "0001111011100" => data_out <= rom_array(988);
		when "0001111011101" => data_out <= rom_array(989);
		when "0001111011110" => data_out <= rom_array(990);
		when "0001111011111" => data_out <= rom_array(991);
		when "0001111100000" => data_out <= rom_array(992);
		when "0001111100001" => data_out <= rom_array(993);
		when "0001111100010" => data_out <= rom_array(994);
		when "0001111100011" => data_out <= rom_array(995);
		when "0001111100100" => data_out <= rom_array(996);
		when "0001111100101" => data_out <= rom_array(997);
		when "0001111100110" => data_out <= rom_array(998);
		when "0001111100111" => data_out <= rom_array(999);
		when "0001111101000" => data_out <= rom_array(1000);
		when "0001111101001" => data_out <= rom_array(1001);
		when "0001111101010" => data_out <= rom_array(1002);
		when "0001111101011" => data_out <= rom_array(1003);
		when "0001111101100" => data_out <= rom_array(1004);
		when "0001111101101" => data_out <= rom_array(1005);
		when "0001111101110" => data_out <= rom_array(1006);
		when "0001111101111" => data_out <= rom_array(1007);
		when "0001111110000" => data_out <= rom_array(1008);
		when "0001111110001" => data_out <= rom_array(1009);
		when "0001111110010" => data_out <= rom_array(1010);
		when "0001111110011" => data_out <= rom_array(1011);
		when "0001111110100" => data_out <= rom_array(1012);
		when "0001111110101" => data_out <= rom_array(1013);
		when "0001111110110" => data_out <= rom_array(1014);
		when "0001111110111" => data_out <= rom_array(1015);
		when "0001111111000" => data_out <= rom_array(1016);
		when "0001111111001" => data_out <= rom_array(1017);
		when "0001111111010" => data_out <= rom_array(1018);
		when "0001111111011" => data_out <= rom_array(1019);
		when "0001111111100" => data_out <= rom_array(1020);
		when "0001111111101" => data_out <= rom_array(1021);
		when "0001111111110" => data_out <= rom_array(1022);
		when "0001111111111" => data_out <= rom_array(1023);
		when "0010000000000" => data_out <= rom_array(1024);
		when "0010000000001" => data_out <= rom_array(1025);
		when "0010000000010" => data_out <= rom_array(1026);
		when "0010000000011" => data_out <= rom_array(1027);
		when "0010000000100" => data_out <= rom_array(1028);
		when "0010000000101" => data_out <= rom_array(1029);
		when "0010000000110" => data_out <= rom_array(1030);
		when "0010000000111" => data_out <= rom_array(1031);
		when "0010000001000" => data_out <= rom_array(1032);
		when "0010000001001" => data_out <= rom_array(1033);
		when "0010000001010" => data_out <= rom_array(1034);
		when "0010000001011" => data_out <= rom_array(1035);
		when "0010000001100" => data_out <= rom_array(1036);
		when "0010000001101" => data_out <= rom_array(1037);
		when "0010000001110" => data_out <= rom_array(1038);
		when "0010000001111" => data_out <= rom_array(1039);
		when "0010000010000" => data_out <= rom_array(1040);
		when "0010000010001" => data_out <= rom_array(1041);
		when "0010000010010" => data_out <= rom_array(1042);
		when "0010000010011" => data_out <= rom_array(1043);
		when "0010000010100" => data_out <= rom_array(1044);
		when "0010000010101" => data_out <= rom_array(1045);
		when "0010000010110" => data_out <= rom_array(1046);
		when "0010000010111" => data_out <= rom_array(1047);
		when "0010000011000" => data_out <= rom_array(1048);
		when "0010000011001" => data_out <= rom_array(1049);
		when "0010000011010" => data_out <= rom_array(1050);
		when "0010000011011" => data_out <= rom_array(1051);
		when "0010000011100" => data_out <= rom_array(1052);
		when "0010000011101" => data_out <= rom_array(1053);
		when "0010000011110" => data_out <= rom_array(1054);
		when "0010000011111" => data_out <= rom_array(1055);
		when "0010000100000" => data_out <= rom_array(1056);
		when "0010000100001" => data_out <= rom_array(1057);
		when "0010000100010" => data_out <= rom_array(1058);
		when "0010000100011" => data_out <= rom_array(1059);
		when "0010000100100" => data_out <= rom_array(1060);
		when "0010000100101" => data_out <= rom_array(1061);
		when "0010000100110" => data_out <= rom_array(1062);
		when "0010000100111" => data_out <= rom_array(1063);
		when "0010000101000" => data_out <= rom_array(1064);
		when "0010000101001" => data_out <= rom_array(1065);
		when "0010000101010" => data_out <= rom_array(1066);
		when "0010000101011" => data_out <= rom_array(1067);
		when "0010000101100" => data_out <= rom_array(1068);
		when "0010000101101" => data_out <= rom_array(1069);
		when "0010000101110" => data_out <= rom_array(1070);
		when "0010000101111" => data_out <= rom_array(1071);
		when "0010000110000" => data_out <= rom_array(1072);
		when "0010000110001" => data_out <= rom_array(1073);
		when "0010000110010" => data_out <= rom_array(1074);
		when "0010000110011" => data_out <= rom_array(1075);
		when "0010000110100" => data_out <= rom_array(1076);
		when "0010000110101" => data_out <= rom_array(1077);
		when "0010000110110" => data_out <= rom_array(1078);
		when "0010000110111" => data_out <= rom_array(1079);
		when "0010000111000" => data_out <= rom_array(1080);
		when "0010000111001" => data_out <= rom_array(1081);
		when "0010000111010" => data_out <= rom_array(1082);
		when "0010000111011" => data_out <= rom_array(1083);
		when "0010000111100" => data_out <= rom_array(1084);
		when "0010000111101" => data_out <= rom_array(1085);
		when "0010000111110" => data_out <= rom_array(1086);
		when "0010000111111" => data_out <= rom_array(1087);
		when "0010001000000" => data_out <= rom_array(1088);
		when "0010001000001" => data_out <= rom_array(1089);
		when "0010001000010" => data_out <= rom_array(1090);
		when "0010001000011" => data_out <= rom_array(1091);
		when "0010001000100" => data_out <= rom_array(1092);
		when "0010001000101" => data_out <= rom_array(1093);
		when "0010001000110" => data_out <= rom_array(1094);
		when "0010001000111" => data_out <= rom_array(1095);
		when "0010001001000" => data_out <= rom_array(1096);
		when "0010001001001" => data_out <= rom_array(1097);
		when "0010001001010" => data_out <= rom_array(1098);
		when "0010001001011" => data_out <= rom_array(1099);
		when "0010001001100" => data_out <= rom_array(1100);
		when "0010001001101" => data_out <= rom_array(1101);
		when "0010001001110" => data_out <= rom_array(1102);
		when "0010001001111" => data_out <= rom_array(1103);
		when "0010001010000" => data_out <= rom_array(1104);
		when "0010001010001" => data_out <= rom_array(1105);
		when "0010001010010" => data_out <= rom_array(1106);
		when "0010001010011" => data_out <= rom_array(1107);
		when "0010001010100" => data_out <= rom_array(1108);
		when "0010001010101" => data_out <= rom_array(1109);
		when "0010001010110" => data_out <= rom_array(1110);
		when "0010001010111" => data_out <= rom_array(1111);
		when "0010001011000" => data_out <= rom_array(1112);
		when "0010001011001" => data_out <= rom_array(1113);
		when "0010001011010" => data_out <= rom_array(1114);
		when "0010001011011" => data_out <= rom_array(1115);
		when "0010001011100" => data_out <= rom_array(1116);
		when "0010001011101" => data_out <= rom_array(1117);
		when "0010001011110" => data_out <= rom_array(1118);
		when "0010001011111" => data_out <= rom_array(1119);
		when "0010001100000" => data_out <= rom_array(1120);
		when "0010001100001" => data_out <= rom_array(1121);
		when "0010001100010" => data_out <= rom_array(1122);
		when "0010001100011" => data_out <= rom_array(1123);
		when "0010001100100" => data_out <= rom_array(1124);
		when "0010001100101" => data_out <= rom_array(1125);
		when "0010001100110" => data_out <= rom_array(1126);
		when "0010001100111" => data_out <= rom_array(1127);
		when "0010001101000" => data_out <= rom_array(1128);
		when "0010001101001" => data_out <= rom_array(1129);
		when "0010001101010" => data_out <= rom_array(1130);
		when "0010001101011" => data_out <= rom_array(1131);
		when "0010001101100" => data_out <= rom_array(1132);
		when "0010001101101" => data_out <= rom_array(1133);
		when "0010001101110" => data_out <= rom_array(1134);
		when "0010001101111" => data_out <= rom_array(1135);
		when "0010001110000" => data_out <= rom_array(1136);
		when "0010001110001" => data_out <= rom_array(1137);
		when "0010001110010" => data_out <= rom_array(1138);
		when "0010001110011" => data_out <= rom_array(1139);
		when "0010001110100" => data_out <= rom_array(1140);
		when "0010001110101" => data_out <= rom_array(1141);
		when "0010001110110" => data_out <= rom_array(1142);
		when "0010001110111" => data_out <= rom_array(1143);
		when "0010001111000" => data_out <= rom_array(1144);
		when "0010001111001" => data_out <= rom_array(1145);
		when "0010001111010" => data_out <= rom_array(1146);
		when "0010001111011" => data_out <= rom_array(1147);
		when "0010001111100" => data_out <= rom_array(1148);
		when "0010001111101" => data_out <= rom_array(1149);
		when "0010001111110" => data_out <= rom_array(1150);
		when "0010001111111" => data_out <= rom_array(1151);
		when "0010010000000" => data_out <= rom_array(1152);
		when "0010010000001" => data_out <= rom_array(1153);
		when "0010010000010" => data_out <= rom_array(1154);
		when "0010010000011" => data_out <= rom_array(1155);
		when "0010010000100" => data_out <= rom_array(1156);
		when "0010010000101" => data_out <= rom_array(1157);
		when "0010010000110" => data_out <= rom_array(1158);
		when "0010010000111" => data_out <= rom_array(1159);
		when "0010010001000" => data_out <= rom_array(1160);
		when "0010010001001" => data_out <= rom_array(1161);
		when "0010010001010" => data_out <= rom_array(1162);
		when "0010010001011" => data_out <= rom_array(1163);
		when "0010010001100" => data_out <= rom_array(1164);
		when "0010010001101" => data_out <= rom_array(1165);
		when "0010010001110" => data_out <= rom_array(1166);
		when "0010010001111" => data_out <= rom_array(1167);
		when "0010010010000" => data_out <= rom_array(1168);
		when "0010010010001" => data_out <= rom_array(1169);
		when "0010010010010" => data_out <= rom_array(1170);
		when "0010010010011" => data_out <= rom_array(1171);
		when "0010010010100" => data_out <= rom_array(1172);
		when "0010010010101" => data_out <= rom_array(1173);
		when "0010010010110" => data_out <= rom_array(1174);
		when "0010010010111" => data_out <= rom_array(1175);
		when "0010010011000" => data_out <= rom_array(1176);
		when "0010010011001" => data_out <= rom_array(1177);
		when "0010010011010" => data_out <= rom_array(1178);
		when "0010010011011" => data_out <= rom_array(1179);
		when "0010010011100" => data_out <= rom_array(1180);
		when "0010010011101" => data_out <= rom_array(1181);
		when "0010010011110" => data_out <= rom_array(1182);
		when "0010010011111" => data_out <= rom_array(1183);
		when "0010010100000" => data_out <= rom_array(1184);
		when "0010010100001" => data_out <= rom_array(1185);
		when "0010010100010" => data_out <= rom_array(1186);
		when "0010010100011" => data_out <= rom_array(1187);
		when "0010010100100" => data_out <= rom_array(1188);
		when "0010010100101" => data_out <= rom_array(1189);
		when "0010010100110" => data_out <= rom_array(1190);
		when "0010010100111" => data_out <= rom_array(1191);
		when "0010010101000" => data_out <= rom_array(1192);
		when "0010010101001" => data_out <= rom_array(1193);
		when "0010010101010" => data_out <= rom_array(1194);
		when "0010010101011" => data_out <= rom_array(1195);
		when "0010010101100" => data_out <= rom_array(1196);
		when "0010010101101" => data_out <= rom_array(1197);
		when "0010010101110" => data_out <= rom_array(1198);
		when "0010010101111" => data_out <= rom_array(1199);
		when "0010010110000" => data_out <= rom_array(1200);
		when "0010010110001" => data_out <= rom_array(1201);
		when "0010010110010" => data_out <= rom_array(1202);
		when "0010010110011" => data_out <= rom_array(1203);
		when "0010010110100" => data_out <= rom_array(1204);
		when "0010010110101" => data_out <= rom_array(1205);
		when "0010010110110" => data_out <= rom_array(1206);
		when "0010010110111" => data_out <= rom_array(1207);
		when "0010010111000" => data_out <= rom_array(1208);
		when "0010010111001" => data_out <= rom_array(1209);
		when "0010010111010" => data_out <= rom_array(1210);
		when "0010010111011" => data_out <= rom_array(1211);
		when "0010010111100" => data_out <= rom_array(1212);
		when "0010010111101" => data_out <= rom_array(1213);
		when "0010010111110" => data_out <= rom_array(1214);
		when "0010010111111" => data_out <= rom_array(1215);
		when "0010011000000" => data_out <= rom_array(1216);
		when "0010011000001" => data_out <= rom_array(1217);
		when "0010011000010" => data_out <= rom_array(1218);
		when "0010011000011" => data_out <= rom_array(1219);
		when "0010011000100" => data_out <= rom_array(1220);
		when "0010011000101" => data_out <= rom_array(1221);
		when "0010011000110" => data_out <= rom_array(1222);
		when "0010011000111" => data_out <= rom_array(1223);
		when "0010011001000" => data_out <= rom_array(1224);
		when "0010011001001" => data_out <= rom_array(1225);
		when "0010011001010" => data_out <= rom_array(1226);
		when "0010011001011" => data_out <= rom_array(1227);
		when "0010011001100" => data_out <= rom_array(1228);
		when "0010011001101" => data_out <= rom_array(1229);
		when "0010011001110" => data_out <= rom_array(1230);
		when "0010011001111" => data_out <= rom_array(1231);
		when "0010011010000" => data_out <= rom_array(1232);
		when "0010011010001" => data_out <= rom_array(1233);
		when "0010011010010" => data_out <= rom_array(1234);
		when "0010011010011" => data_out <= rom_array(1235);
		when "0010011010100" => data_out <= rom_array(1236);
		when "0010011010101" => data_out <= rom_array(1237);
		when "0010011010110" => data_out <= rom_array(1238);
		when "0010011010111" => data_out <= rom_array(1239);
		when "0010011011000" => data_out <= rom_array(1240);
		when "0010011011001" => data_out <= rom_array(1241);
		when "0010011011010" => data_out <= rom_array(1242);
		when "0010011011011" => data_out <= rom_array(1243);
		when "0010011011100" => data_out <= rom_array(1244);
		when "0010011011101" => data_out <= rom_array(1245);
		when "0010011011110" => data_out <= rom_array(1246);
		when "0010011011111" => data_out <= rom_array(1247);
		when "0010011100000" => data_out <= rom_array(1248);
		when "0010011100001" => data_out <= rom_array(1249);
		when "0010011100010" => data_out <= rom_array(1250);
		when "0010011100011" => data_out <= rom_array(1251);
		when "0010011100100" => data_out <= rom_array(1252);
		when "0010011100101" => data_out <= rom_array(1253);
		when "0010011100110" => data_out <= rom_array(1254);
		when "0010011100111" => data_out <= rom_array(1255);
		when "0010011101000" => data_out <= rom_array(1256);
		when "0010011101001" => data_out <= rom_array(1257);
		when "0010011101010" => data_out <= rom_array(1258);
		when "0010011101011" => data_out <= rom_array(1259);
		when "0010011101100" => data_out <= rom_array(1260);
		when "0010011101101" => data_out <= rom_array(1261);
		when "0010011101110" => data_out <= rom_array(1262);
		when "0010011101111" => data_out <= rom_array(1263);
		when "0010011110000" => data_out <= rom_array(1264);
		when "0010011110001" => data_out <= rom_array(1265);
		when "0010011110010" => data_out <= rom_array(1266);
		when "0010011110011" => data_out <= rom_array(1267);
		when "0010011110100" => data_out <= rom_array(1268);
		when "0010011110101" => data_out <= rom_array(1269);
		when "0010011110110" => data_out <= rom_array(1270);
		when "0010011110111" => data_out <= rom_array(1271);
		when "0010011111000" => data_out <= rom_array(1272);
		when "0010011111001" => data_out <= rom_array(1273);
		when "0010011111010" => data_out <= rom_array(1274);
		when "0010011111011" => data_out <= rom_array(1275);
		when "0010011111100" => data_out <= rom_array(1276);
		when "0010011111101" => data_out <= rom_array(1277);
		when "0010011111110" => data_out <= rom_array(1278);
		when "0010011111111" => data_out <= rom_array(1279);
		when "0010100000000" => data_out <= rom_array(1280);
		when "0010100000001" => data_out <= rom_array(1281);
		when "0010100000010" => data_out <= rom_array(1282);
		when "0010100000011" => data_out <= rom_array(1283);
		when "0010100000100" => data_out <= rom_array(1284);
		when "0010100000101" => data_out <= rom_array(1285);
		when "0010100000110" => data_out <= rom_array(1286);
		when "0010100000111" => data_out <= rom_array(1287);
		when "0010100001000" => data_out <= rom_array(1288);
		when "0010100001001" => data_out <= rom_array(1289);
		when "0010100001010" => data_out <= rom_array(1290);
		when "0010100001011" => data_out <= rom_array(1291);
		when "0010100001100" => data_out <= rom_array(1292);
		when "0010100001101" => data_out <= rom_array(1293);
		when "0010100001110" => data_out <= rom_array(1294);
		when "0010100001111" => data_out <= rom_array(1295);
		when "0010100010000" => data_out <= rom_array(1296);
		when "0010100010001" => data_out <= rom_array(1297);
		when "0010100010010" => data_out <= rom_array(1298);
		when "0010100010011" => data_out <= rom_array(1299);
		when "0010100010100" => data_out <= rom_array(1300);
		when "0010100010101" => data_out <= rom_array(1301);
		when "0010100010110" => data_out <= rom_array(1302);
		when "0010100010111" => data_out <= rom_array(1303);
		when "0010100011000" => data_out <= rom_array(1304);
		when "0010100011001" => data_out <= rom_array(1305);
		when "0010100011010" => data_out <= rom_array(1306);
		when "0010100011011" => data_out <= rom_array(1307);
		when "0010100011100" => data_out <= rom_array(1308);
		when "0010100011101" => data_out <= rom_array(1309);
		when "0010100011110" => data_out <= rom_array(1310);
		when "0010100011111" => data_out <= rom_array(1311);
		when "0010100100000" => data_out <= rom_array(1312);
		when "0010100100001" => data_out <= rom_array(1313);
		when "0010100100010" => data_out <= rom_array(1314);
		when "0010100100011" => data_out <= rom_array(1315);
		when "0010100100100" => data_out <= rom_array(1316);
		when "0010100100101" => data_out <= rom_array(1317);
		when "0010100100110" => data_out <= rom_array(1318);
		when "0010100100111" => data_out <= rom_array(1319);
		when "0010100101000" => data_out <= rom_array(1320);
		when "0010100101001" => data_out <= rom_array(1321);
		when "0010100101010" => data_out <= rom_array(1322);
		when "0010100101011" => data_out <= rom_array(1323);
		when "0010100101100" => data_out <= rom_array(1324);
		when "0010100101101" => data_out <= rom_array(1325);
		when "0010100101110" => data_out <= rom_array(1326);
		when "0010100101111" => data_out <= rom_array(1327);
		when "0010100110000" => data_out <= rom_array(1328);
		when "0010100110001" => data_out <= rom_array(1329);
		when "0010100110010" => data_out <= rom_array(1330);
		when "0010100110011" => data_out <= rom_array(1331);
		when "0010100110100" => data_out <= rom_array(1332);
		when "0010100110101" => data_out <= rom_array(1333);
		when "0010100110110" => data_out <= rom_array(1334);
		when "0010100110111" => data_out <= rom_array(1335);
		when "0010100111000" => data_out <= rom_array(1336);
		when "0010100111001" => data_out <= rom_array(1337);
		when "0010100111010" => data_out <= rom_array(1338);
		when "0010100111011" => data_out <= rom_array(1339);
		when "0010100111100" => data_out <= rom_array(1340);
		when "0010100111101" => data_out <= rom_array(1341);
		when "0010100111110" => data_out <= rom_array(1342);
		when "0010100111111" => data_out <= rom_array(1343);
		when "0010101000000" => data_out <= rom_array(1344);
		when "0010101000001" => data_out <= rom_array(1345);
		when "0010101000010" => data_out <= rom_array(1346);
		when "0010101000011" => data_out <= rom_array(1347);
		when "0010101000100" => data_out <= rom_array(1348);
		when "0010101000101" => data_out <= rom_array(1349);
		when "0010101000110" => data_out <= rom_array(1350);
		when "0010101000111" => data_out <= rom_array(1351);
		when "0010101001000" => data_out <= rom_array(1352);
		when "0010101001001" => data_out <= rom_array(1353);
		when "0010101001010" => data_out <= rom_array(1354);
		when "0010101001011" => data_out <= rom_array(1355);
		when "0010101001100" => data_out <= rom_array(1356);
		when "0010101001101" => data_out <= rom_array(1357);
		when "0010101001110" => data_out <= rom_array(1358);
		when "0010101001111" => data_out <= rom_array(1359);
		when "0010101010000" => data_out <= rom_array(1360);
		when "0010101010001" => data_out <= rom_array(1361);
		when "0010101010010" => data_out <= rom_array(1362);
		when "0010101010011" => data_out <= rom_array(1363);
		when "0010101010100" => data_out <= rom_array(1364);
		when "0010101010101" => data_out <= rom_array(1365);
		when "0010101010110" => data_out <= rom_array(1366);
		when "0010101010111" => data_out <= rom_array(1367);
		when "0010101011000" => data_out <= rom_array(1368);
		when "0010101011001" => data_out <= rom_array(1369);
		when "0010101011010" => data_out <= rom_array(1370);
		when "0010101011011" => data_out <= rom_array(1371);
		when "0010101011100" => data_out <= rom_array(1372);
		when "0010101011101" => data_out <= rom_array(1373);
		when "0010101011110" => data_out <= rom_array(1374);
		when "0010101011111" => data_out <= rom_array(1375);
		when "0010101100000" => data_out <= rom_array(1376);
		when "0010101100001" => data_out <= rom_array(1377);
		when "0010101100010" => data_out <= rom_array(1378);
		when "0010101100011" => data_out <= rom_array(1379);
		when "0010101100100" => data_out <= rom_array(1380);
		when "0010101100101" => data_out <= rom_array(1381);
		when "0010101100110" => data_out <= rom_array(1382);
		when "0010101100111" => data_out <= rom_array(1383);
		when "0010101101000" => data_out <= rom_array(1384);
		when "0010101101001" => data_out <= rom_array(1385);
		when "0010101101010" => data_out <= rom_array(1386);
		when "0010101101011" => data_out <= rom_array(1387);
		when "0010101101100" => data_out <= rom_array(1388);
		when "0010101101101" => data_out <= rom_array(1389);
		when "0010101101110" => data_out <= rom_array(1390);
		when "0010101101111" => data_out <= rom_array(1391);
		when "0010101110000" => data_out <= rom_array(1392);
		when "0010101110001" => data_out <= rom_array(1393);
		when "0010101110010" => data_out <= rom_array(1394);
		when "0010101110011" => data_out <= rom_array(1395);
		when "0010101110100" => data_out <= rom_array(1396);
		when "0010101110101" => data_out <= rom_array(1397);
		when "0010101110110" => data_out <= rom_array(1398);
		when "0010101110111" => data_out <= rom_array(1399);
		when "0010101111000" => data_out <= rom_array(1400);
		when "0010101111001" => data_out <= rom_array(1401);
		when "0010101111010" => data_out <= rom_array(1402);
		when "0010101111011" => data_out <= rom_array(1403);
		when "0010101111100" => data_out <= rom_array(1404);
		when "0010101111101" => data_out <= rom_array(1405);
		when "0010101111110" => data_out <= rom_array(1406);
		when "0010101111111" => data_out <= rom_array(1407);
		when "0010110000000" => data_out <= rom_array(1408);
		when "0010110000001" => data_out <= rom_array(1409);
		when "0010110000010" => data_out <= rom_array(1410);
		when "0010110000011" => data_out <= rom_array(1411);
		when "0010110000100" => data_out <= rom_array(1412);
		when "0010110000101" => data_out <= rom_array(1413);
		when "0010110000110" => data_out <= rom_array(1414);
		when "0010110000111" => data_out <= rom_array(1415);
		when "0010110001000" => data_out <= rom_array(1416);
		when "0010110001001" => data_out <= rom_array(1417);
		when "0010110001010" => data_out <= rom_array(1418);
		when "0010110001011" => data_out <= rom_array(1419);
		when "0010110001100" => data_out <= rom_array(1420);
		when "0010110001101" => data_out <= rom_array(1421);
		when "0010110001110" => data_out <= rom_array(1422);
		when "0010110001111" => data_out <= rom_array(1423);
		when "0010110010000" => data_out <= rom_array(1424);
		when "0010110010001" => data_out <= rom_array(1425);
		when "0010110010010" => data_out <= rom_array(1426);
		when "0010110010011" => data_out <= rom_array(1427);
		when "0010110010100" => data_out <= rom_array(1428);
		when "0010110010101" => data_out <= rom_array(1429);
		when "0010110010110" => data_out <= rom_array(1430);
		when "0010110010111" => data_out <= rom_array(1431);
		when "0010110011000" => data_out <= rom_array(1432);
		when "0010110011001" => data_out <= rom_array(1433);
		when "0010110011010" => data_out <= rom_array(1434);
		when "0010110011011" => data_out <= rom_array(1435);
		when "0010110011100" => data_out <= rom_array(1436);
		when "0010110011101" => data_out <= rom_array(1437);
		when "0010110011110" => data_out <= rom_array(1438);
		when "0010110011111" => data_out <= rom_array(1439);
		when "0010110100000" => data_out <= rom_array(1440);
		when "0010110100001" => data_out <= rom_array(1441);
		when "0010110100010" => data_out <= rom_array(1442);
		when "0010110100011" => data_out <= rom_array(1443);
		when "0010110100100" => data_out <= rom_array(1444);
		when "0010110100101" => data_out <= rom_array(1445);
		when "0010110100110" => data_out <= rom_array(1446);
		when "0010110100111" => data_out <= rom_array(1447);
		when "0010110101000" => data_out <= rom_array(1448);
		when "0010110101001" => data_out <= rom_array(1449);
		when "0010110101010" => data_out <= rom_array(1450);
		when "0010110101011" => data_out <= rom_array(1451);
		when "0010110101100" => data_out <= rom_array(1452);
		when "0010110101101" => data_out <= rom_array(1453);
		when "0010110101110" => data_out <= rom_array(1454);
		when "0010110101111" => data_out <= rom_array(1455);
		when "0010110110000" => data_out <= rom_array(1456);
		when "0010110110001" => data_out <= rom_array(1457);
		when "0010110110010" => data_out <= rom_array(1458);
		when "0010110110011" => data_out <= rom_array(1459);
		when "0010110110100" => data_out <= rom_array(1460);
		when "0010110110101" => data_out <= rom_array(1461);
		when "0010110110110" => data_out <= rom_array(1462);
		when "0010110110111" => data_out <= rom_array(1463);
		when "0010110111000" => data_out <= rom_array(1464);
		when "0010110111001" => data_out <= rom_array(1465);
		when "0010110111010" => data_out <= rom_array(1466);
		when "0010110111011" => data_out <= rom_array(1467);
		when "0010110111100" => data_out <= rom_array(1468);
		when "0010110111101" => data_out <= rom_array(1469);
		when "0010110111110" => data_out <= rom_array(1470);
		when "0010110111111" => data_out <= rom_array(1471);
		when "0010111000000" => data_out <= rom_array(1472);
		when "0010111000001" => data_out <= rom_array(1473);
		when "0010111000010" => data_out <= rom_array(1474);
		when "0010111000011" => data_out <= rom_array(1475);
		when "0010111000100" => data_out <= rom_array(1476);
		when "0010111000101" => data_out <= rom_array(1477);
		when "0010111000110" => data_out <= rom_array(1478);
		when "0010111000111" => data_out <= rom_array(1479);
		when "0010111001000" => data_out <= rom_array(1480);
		when "0010111001001" => data_out <= rom_array(1481);
		when "0010111001010" => data_out <= rom_array(1482);
		when "0010111001011" => data_out <= rom_array(1483);
		when "0010111001100" => data_out <= rom_array(1484);
		when "0010111001101" => data_out <= rom_array(1485);
		when "0010111001110" => data_out <= rom_array(1486);
		when "0010111001111" => data_out <= rom_array(1487);
		when "0010111010000" => data_out <= rom_array(1488);
		when "0010111010001" => data_out <= rom_array(1489);
		when "0010111010010" => data_out <= rom_array(1490);
		when "0010111010011" => data_out <= rom_array(1491);
		when "0010111010100" => data_out <= rom_array(1492);
		when "0010111010101" => data_out <= rom_array(1493);
		when "0010111010110" => data_out <= rom_array(1494);
		when "0010111010111" => data_out <= rom_array(1495);
		when "0010111011000" => data_out <= rom_array(1496);
		when "0010111011001" => data_out <= rom_array(1497);
		when "0010111011010" => data_out <= rom_array(1498);
		when "0010111011011" => data_out <= rom_array(1499);
		when "0010111011100" => data_out <= rom_array(1500);
		when "0010111011101" => data_out <= rom_array(1501);
		when "0010111011110" => data_out <= rom_array(1502);
		when "0010111011111" => data_out <= rom_array(1503);
		when "0010111100000" => data_out <= rom_array(1504);
		when "0010111100001" => data_out <= rom_array(1505);
		when "0010111100010" => data_out <= rom_array(1506);
		when "0010111100011" => data_out <= rom_array(1507);
		when "0010111100100" => data_out <= rom_array(1508);
		when "0010111100101" => data_out <= rom_array(1509);
		when "0010111100110" => data_out <= rom_array(1510);
		when "0010111100111" => data_out <= rom_array(1511);
		when "0010111101000" => data_out <= rom_array(1512);
		when "0010111101001" => data_out <= rom_array(1513);
		when "0010111101010" => data_out <= rom_array(1514);
		when "0010111101011" => data_out <= rom_array(1515);
		when "0010111101100" => data_out <= rom_array(1516);
		when "0010111101101" => data_out <= rom_array(1517);
		when "0010111101110" => data_out <= rom_array(1518);
		when "0010111101111" => data_out <= rom_array(1519);
		when "0010111110000" => data_out <= rom_array(1520);
		when "0010111110001" => data_out <= rom_array(1521);
		when "0010111110010" => data_out <= rom_array(1522);
		when "0010111110011" => data_out <= rom_array(1523);
		when "0010111110100" => data_out <= rom_array(1524);
		when "0010111110101" => data_out <= rom_array(1525);
		when "0010111110110" => data_out <= rom_array(1526);
		when "0010111110111" => data_out <= rom_array(1527);
		when "0010111111000" => data_out <= rom_array(1528);
		when "0010111111001" => data_out <= rom_array(1529);
		when "0010111111010" => data_out <= rom_array(1530);
		when "0010111111011" => data_out <= rom_array(1531);
		when "0010111111100" => data_out <= rom_array(1532);
		when "0010111111101" => data_out <= rom_array(1533);
		when "0010111111110" => data_out <= rom_array(1534);
		when "0010111111111" => data_out <= rom_array(1535);
		when "0011000000000" => data_out <= rom_array(1536);
		when "0011000000001" => data_out <= rom_array(1537);
		when "0011000000010" => data_out <= rom_array(1538);
		when "0011000000011" => data_out <= rom_array(1539);
		when "0011000000100" => data_out <= rom_array(1540);
		when "0011000000101" => data_out <= rom_array(1541);
		when "0011000000110" => data_out <= rom_array(1542);
		when "0011000000111" => data_out <= rom_array(1543);
		when "0011000001000" => data_out <= rom_array(1544);
		when "0011000001001" => data_out <= rom_array(1545);
		when "0011000001010" => data_out <= rom_array(1546);
		when "0011000001011" => data_out <= rom_array(1547);
		when "0011000001100" => data_out <= rom_array(1548);
		when "0011000001101" => data_out <= rom_array(1549);
		when "0011000001110" => data_out <= rom_array(1550);
		when "0011000001111" => data_out <= rom_array(1551);
		when "0011000010000" => data_out <= rom_array(1552);
		when "0011000010001" => data_out <= rom_array(1553);
		when "0011000010010" => data_out <= rom_array(1554);
		when "0011000010011" => data_out <= rom_array(1555);
		when "0011000010100" => data_out <= rom_array(1556);
		when "0011000010101" => data_out <= rom_array(1557);
		when "0011000010110" => data_out <= rom_array(1558);
		when "0011000010111" => data_out <= rom_array(1559);
		when "0011000011000" => data_out <= rom_array(1560);
		when "0011000011001" => data_out <= rom_array(1561);
		when "0011000011010" => data_out <= rom_array(1562);
		when "0011000011011" => data_out <= rom_array(1563);
		when "0011000011100" => data_out <= rom_array(1564);
		when "0011000011101" => data_out <= rom_array(1565);
		when "0011000011110" => data_out <= rom_array(1566);
		when "0011000011111" => data_out <= rom_array(1567);
		when "0011000100000" => data_out <= rom_array(1568);
		when "0011000100001" => data_out <= rom_array(1569);
		when "0011000100010" => data_out <= rom_array(1570);
		when "0011000100011" => data_out <= rom_array(1571);
		when "0011000100100" => data_out <= rom_array(1572);
		when "0011000100101" => data_out <= rom_array(1573);
		when "0011000100110" => data_out <= rom_array(1574);
		when "0011000100111" => data_out <= rom_array(1575);
		when "0011000101000" => data_out <= rom_array(1576);
		when "0011000101001" => data_out <= rom_array(1577);
		when "0011000101010" => data_out <= rom_array(1578);
		when "0011000101011" => data_out <= rom_array(1579);
		when "0011000101100" => data_out <= rom_array(1580);
		when "0011000101101" => data_out <= rom_array(1581);
		when "0011000101110" => data_out <= rom_array(1582);
		when "0011000101111" => data_out <= rom_array(1583);
		when "0011000110000" => data_out <= rom_array(1584);
		when "0011000110001" => data_out <= rom_array(1585);
		when "0011000110010" => data_out <= rom_array(1586);
		when "0011000110011" => data_out <= rom_array(1587);
		when "0011000110100" => data_out <= rom_array(1588);
		when "0011000110101" => data_out <= rom_array(1589);
		when "0011000110110" => data_out <= rom_array(1590);
		when "0011000110111" => data_out <= rom_array(1591);
		when "0011000111000" => data_out <= rom_array(1592);
		when "0011000111001" => data_out <= rom_array(1593);
		when "0011000111010" => data_out <= rom_array(1594);
		when "0011000111011" => data_out <= rom_array(1595);
		when "0011000111100" => data_out <= rom_array(1596);
		when "0011000111101" => data_out <= rom_array(1597);
		when "0011000111110" => data_out <= rom_array(1598);
		when "0011000111111" => data_out <= rom_array(1599);
		when "0011001000000" => data_out <= rom_array(1600);
		when "0011001000001" => data_out <= rom_array(1601);
		when "0011001000010" => data_out <= rom_array(1602);
		when "0011001000011" => data_out <= rom_array(1603);
		when "0011001000100" => data_out <= rom_array(1604);
		when "0011001000101" => data_out <= rom_array(1605);
		when "0011001000110" => data_out <= rom_array(1606);
		when "0011001000111" => data_out <= rom_array(1607);
		when "0011001001000" => data_out <= rom_array(1608);
		when "0011001001001" => data_out <= rom_array(1609);
		when "0011001001010" => data_out <= rom_array(1610);
		when "0011001001011" => data_out <= rom_array(1611);
		when "0011001001100" => data_out <= rom_array(1612);
		when "0011001001101" => data_out <= rom_array(1613);
		when "0011001001110" => data_out <= rom_array(1614);
		when "0011001001111" => data_out <= rom_array(1615);
		when "0011001010000" => data_out <= rom_array(1616);
		when "0011001010001" => data_out <= rom_array(1617);
		when "0011001010010" => data_out <= rom_array(1618);
		when "0011001010011" => data_out <= rom_array(1619);
		when "0011001010100" => data_out <= rom_array(1620);
		when "0011001010101" => data_out <= rom_array(1621);
		when "0011001010110" => data_out <= rom_array(1622);
		when "0011001010111" => data_out <= rom_array(1623);
		when "0011001011000" => data_out <= rom_array(1624);
		when "0011001011001" => data_out <= rom_array(1625);
		when "0011001011010" => data_out <= rom_array(1626);
		when "0011001011011" => data_out <= rom_array(1627);
		when "0011001011100" => data_out <= rom_array(1628);
		when "0011001011101" => data_out <= rom_array(1629);
		when "0011001011110" => data_out <= rom_array(1630);
		when "0011001011111" => data_out <= rom_array(1631);
		when "0011001100000" => data_out <= rom_array(1632);
		when "0011001100001" => data_out <= rom_array(1633);
		when "0011001100010" => data_out <= rom_array(1634);
		when "0011001100011" => data_out <= rom_array(1635);
		when "0011001100100" => data_out <= rom_array(1636);
		when "0011001100101" => data_out <= rom_array(1637);
		when "0011001100110" => data_out <= rom_array(1638);
		when "0011001100111" => data_out <= rom_array(1639);
		when "0011001101000" => data_out <= rom_array(1640);
		when "0011001101001" => data_out <= rom_array(1641);
		when "0011001101010" => data_out <= rom_array(1642);
		when "0011001101011" => data_out <= rom_array(1643);
		when "0011001101100" => data_out <= rom_array(1644);
		when "0011001101101" => data_out <= rom_array(1645);
		when "0011001101110" => data_out <= rom_array(1646);
		when "0011001101111" => data_out <= rom_array(1647);
		when "0011001110000" => data_out <= rom_array(1648);
		when "0011001110001" => data_out <= rom_array(1649);
		when "0011001110010" => data_out <= rom_array(1650);
		when "0011001110011" => data_out <= rom_array(1651);
		when "0011001110100" => data_out <= rom_array(1652);
		when "0011001110101" => data_out <= rom_array(1653);
		when "0011001110110" => data_out <= rom_array(1654);
		when "0011001110111" => data_out <= rom_array(1655);
		when "0011001111000" => data_out <= rom_array(1656);
		when "0011001111001" => data_out <= rom_array(1657);
		when "0011001111010" => data_out <= rom_array(1658);
		when "0011001111011" => data_out <= rom_array(1659);
		when "0011001111100" => data_out <= rom_array(1660);
		when "0011001111101" => data_out <= rom_array(1661);
		when "0011001111110" => data_out <= rom_array(1662);
		when "0011001111111" => data_out <= rom_array(1663);
		when "0011010000000" => data_out <= rom_array(1664);
		when "0011010000001" => data_out <= rom_array(1665);
		when "0011010000010" => data_out <= rom_array(1666);
		when "0011010000011" => data_out <= rom_array(1667);
		when "0011010000100" => data_out <= rom_array(1668);
		when "0011010000101" => data_out <= rom_array(1669);
		when "0011010000110" => data_out <= rom_array(1670);
		when "0011010000111" => data_out <= rom_array(1671);
		when "0011010001000" => data_out <= rom_array(1672);
		when "0011010001001" => data_out <= rom_array(1673);
		when "0011010001010" => data_out <= rom_array(1674);
		when "0011010001011" => data_out <= rom_array(1675);
		when "0011010001100" => data_out <= rom_array(1676);
		when "0011010001101" => data_out <= rom_array(1677);
		when "0011010001110" => data_out <= rom_array(1678);
		when "0011010001111" => data_out <= rom_array(1679);
		when "0011010010000" => data_out <= rom_array(1680);
		when "0011010010001" => data_out <= rom_array(1681);
		when "0011010010010" => data_out <= rom_array(1682);
		when "0011010010011" => data_out <= rom_array(1683);
		when "0011010010100" => data_out <= rom_array(1684);
		when "0011010010101" => data_out <= rom_array(1685);
		when "0011010010110" => data_out <= rom_array(1686);
		when "0011010010111" => data_out <= rom_array(1687);
		when "0011010011000" => data_out <= rom_array(1688);
		when "0011010011001" => data_out <= rom_array(1689);
		when "0011010011010" => data_out <= rom_array(1690);
		when "0011010011011" => data_out <= rom_array(1691);
		when "0011010011100" => data_out <= rom_array(1692);
		when "0011010011101" => data_out <= rom_array(1693);
		when "0011010011110" => data_out <= rom_array(1694);
		when "0011010011111" => data_out <= rom_array(1695);
		when "0011010100000" => data_out <= rom_array(1696);
		when "0011010100001" => data_out <= rom_array(1697);
		when "0011010100010" => data_out <= rom_array(1698);
		when "0011010100011" => data_out <= rom_array(1699);
		when "0011010100100" => data_out <= rom_array(1700);
		when "0011010100101" => data_out <= rom_array(1701);
		when "0011010100110" => data_out <= rom_array(1702);
		when "0011010100111" => data_out <= rom_array(1703);
		when "0011010101000" => data_out <= rom_array(1704);
		when "0011010101001" => data_out <= rom_array(1705);
		when "0011010101010" => data_out <= rom_array(1706);
		when "0011010101011" => data_out <= rom_array(1707);
		when "0011010101100" => data_out <= rom_array(1708);
		when "0011010101101" => data_out <= rom_array(1709);
		when "0011010101110" => data_out <= rom_array(1710);
		when "0011010101111" => data_out <= rom_array(1711);
		when "0011010110000" => data_out <= rom_array(1712);
		when "0011010110001" => data_out <= rom_array(1713);
		when "0011010110010" => data_out <= rom_array(1714);
		when "0011010110011" => data_out <= rom_array(1715);
		when "0011010110100" => data_out <= rom_array(1716);
		when "0011010110101" => data_out <= rom_array(1717);
		when "0011010110110" => data_out <= rom_array(1718);
		when "0011010110111" => data_out <= rom_array(1719);
		when "0011010111000" => data_out <= rom_array(1720);
		when "0011010111001" => data_out <= rom_array(1721);
		when "0011010111010" => data_out <= rom_array(1722);
		when "0011010111011" => data_out <= rom_array(1723);
		when "0011010111100" => data_out <= rom_array(1724);
		when "0011010111101" => data_out <= rom_array(1725);
		when "0011010111110" => data_out <= rom_array(1726);
		when "0011010111111" => data_out <= rom_array(1727);
		when "0011011000000" => data_out <= rom_array(1728);
		when "0011011000001" => data_out <= rom_array(1729);
		when "0011011000010" => data_out <= rom_array(1730);
		when "0011011000011" => data_out <= rom_array(1731);
		when "0011011000100" => data_out <= rom_array(1732);
		when "0011011000101" => data_out <= rom_array(1733);
		when "0011011000110" => data_out <= rom_array(1734);
		when "0011011000111" => data_out <= rom_array(1735);
		when "0011011001000" => data_out <= rom_array(1736);
		when "0011011001001" => data_out <= rom_array(1737);
		when "0011011001010" => data_out <= rom_array(1738);
		when "0011011001011" => data_out <= rom_array(1739);
		when "0011011001100" => data_out <= rom_array(1740);
		when "0011011001101" => data_out <= rom_array(1741);
		when "0011011001110" => data_out <= rom_array(1742);
		when "0011011001111" => data_out <= rom_array(1743);
		when "0011011010000" => data_out <= rom_array(1744);
		when "0011011010001" => data_out <= rom_array(1745);
		when "0011011010010" => data_out <= rom_array(1746);
		when "0011011010011" => data_out <= rom_array(1747);
		when "0011011010100" => data_out <= rom_array(1748);
		when "0011011010101" => data_out <= rom_array(1749);
		when "0011011010110" => data_out <= rom_array(1750);
		when "0011011010111" => data_out <= rom_array(1751);
		when "0011011011000" => data_out <= rom_array(1752);
		when "0011011011001" => data_out <= rom_array(1753);
		when "0011011011010" => data_out <= rom_array(1754);
		when "0011011011011" => data_out <= rom_array(1755);
		when "0011011011100" => data_out <= rom_array(1756);
		when "0011011011101" => data_out <= rom_array(1757);
		when "0011011011110" => data_out <= rom_array(1758);
		when "0011011011111" => data_out <= rom_array(1759);
		when "0011011100000" => data_out <= rom_array(1760);
		when "0011011100001" => data_out <= rom_array(1761);
		when "0011011100010" => data_out <= rom_array(1762);
		when "0011011100011" => data_out <= rom_array(1763);
		when "0011011100100" => data_out <= rom_array(1764);
		when "0011011100101" => data_out <= rom_array(1765);
		when "0011011100110" => data_out <= rom_array(1766);
		when "0011011100111" => data_out <= rom_array(1767);
		when "0011011101000" => data_out <= rom_array(1768);
		when "0011011101001" => data_out <= rom_array(1769);
		when "0011011101010" => data_out <= rom_array(1770);
		when "0011011101011" => data_out <= rom_array(1771);
		when "0011011101100" => data_out <= rom_array(1772);
		when "0011011101101" => data_out <= rom_array(1773);
		when "0011011101110" => data_out <= rom_array(1774);
		when "0011011101111" => data_out <= rom_array(1775);
		when "0011011110000" => data_out <= rom_array(1776);
		when "0011011110001" => data_out <= rom_array(1777);
		when "0011011110010" => data_out <= rom_array(1778);
		when "0011011110011" => data_out <= rom_array(1779);
		when "0011011110100" => data_out <= rom_array(1780);
		when "0011011110101" => data_out <= rom_array(1781);
		when "0011011110110" => data_out <= rom_array(1782);
		when "0011011110111" => data_out <= rom_array(1783);
		when "0011011111000" => data_out <= rom_array(1784);
		when "0011011111001" => data_out <= rom_array(1785);
		when "0011011111010" => data_out <= rom_array(1786);
		when "0011011111011" => data_out <= rom_array(1787);
		when "0011011111100" => data_out <= rom_array(1788);
		when "0011011111101" => data_out <= rom_array(1789);
		when "0011011111110" => data_out <= rom_array(1790);
		when "0011011111111" => data_out <= rom_array(1791);
		when "0011100000000" => data_out <= rom_array(1792);
		when "0011100000001" => data_out <= rom_array(1793);
		when "0011100000010" => data_out <= rom_array(1794);
		when "0011100000011" => data_out <= rom_array(1795);
		when "0011100000100" => data_out <= rom_array(1796);
		when "0011100000101" => data_out <= rom_array(1797);
		when "0011100000110" => data_out <= rom_array(1798);
		when "0011100000111" => data_out <= rom_array(1799);
		when "0011100001000" => data_out <= rom_array(1800);
		when "0011100001001" => data_out <= rom_array(1801);
		when "0011100001010" => data_out <= rom_array(1802);
		when "0011100001011" => data_out <= rom_array(1803);
		when "0011100001100" => data_out <= rom_array(1804);
		when "0011100001101" => data_out <= rom_array(1805);
		when "0011100001110" => data_out <= rom_array(1806);
		when "0011100001111" => data_out <= rom_array(1807);
		when "0011100010000" => data_out <= rom_array(1808);
		when "0011100010001" => data_out <= rom_array(1809);
		when "0011100010010" => data_out <= rom_array(1810);
		when "0011100010011" => data_out <= rom_array(1811);
		when "0011100010100" => data_out <= rom_array(1812);
		when "0011100010101" => data_out <= rom_array(1813);
		when "0011100010110" => data_out <= rom_array(1814);
		when "0011100010111" => data_out <= rom_array(1815);
		when "0011100011000" => data_out <= rom_array(1816);
		when "0011100011001" => data_out <= rom_array(1817);
		when "0011100011010" => data_out <= rom_array(1818);
		when "0011100011011" => data_out <= rom_array(1819);
		when "0011100011100" => data_out <= rom_array(1820);
		when "0011100011101" => data_out <= rom_array(1821);
		when "0011100011110" => data_out <= rom_array(1822);
		when "0011100011111" => data_out <= rom_array(1823);
		when "0011100100000" => data_out <= rom_array(1824);
		when "0011100100001" => data_out <= rom_array(1825);
		when "0011100100010" => data_out <= rom_array(1826);
		when "0011100100011" => data_out <= rom_array(1827);
		when "0011100100100" => data_out <= rom_array(1828);
		when "0011100100101" => data_out <= rom_array(1829);
		when "0011100100110" => data_out <= rom_array(1830);
		when "0011100100111" => data_out <= rom_array(1831);
		when "0011100101000" => data_out <= rom_array(1832);
		when "0011100101001" => data_out <= rom_array(1833);
		when "0011100101010" => data_out <= rom_array(1834);
		when "0011100101011" => data_out <= rom_array(1835);
		when "0011100101100" => data_out <= rom_array(1836);
		when "0011100101101" => data_out <= rom_array(1837);
		when "0011100101110" => data_out <= rom_array(1838);
		when "0011100101111" => data_out <= rom_array(1839);
		when "0011100110000" => data_out <= rom_array(1840);
		when "0011100110001" => data_out <= rom_array(1841);
		when "0011100110010" => data_out <= rom_array(1842);
		when "0011100110011" => data_out <= rom_array(1843);
		when "0011100110100" => data_out <= rom_array(1844);
		when "0011100110101" => data_out <= rom_array(1845);
		when "0011100110110" => data_out <= rom_array(1846);
		when "0011100110111" => data_out <= rom_array(1847);
		when "0011100111000" => data_out <= rom_array(1848);
		when "0011100111001" => data_out <= rom_array(1849);
		when "0011100111010" => data_out <= rom_array(1850);
		when "0011100111011" => data_out <= rom_array(1851);
		when "0011100111100" => data_out <= rom_array(1852);
		when "0011100111101" => data_out <= rom_array(1853);
		when "0011100111110" => data_out <= rom_array(1854);
		when "0011100111111" => data_out <= rom_array(1855);
		when "0011101000000" => data_out <= rom_array(1856);
		when "0011101000001" => data_out <= rom_array(1857);
		when "0011101000010" => data_out <= rom_array(1858);
		when "0011101000011" => data_out <= rom_array(1859);
		when "0011101000100" => data_out <= rom_array(1860);
		when "0011101000101" => data_out <= rom_array(1861);
		when "0011101000110" => data_out <= rom_array(1862);
		when "0011101000111" => data_out <= rom_array(1863);
		when "0011101001000" => data_out <= rom_array(1864);
		when "0011101001001" => data_out <= rom_array(1865);
		when "0011101001010" => data_out <= rom_array(1866);
		when "0011101001011" => data_out <= rom_array(1867);
		when "0011101001100" => data_out <= rom_array(1868);
		when "0011101001101" => data_out <= rom_array(1869);
		when "0011101001110" => data_out <= rom_array(1870);
		when "0011101001111" => data_out <= rom_array(1871);
		when "0011101010000" => data_out <= rom_array(1872);
		when "0011101010001" => data_out <= rom_array(1873);
		when "0011101010010" => data_out <= rom_array(1874);
		when "0011101010011" => data_out <= rom_array(1875);
		when "0011101010100" => data_out <= rom_array(1876);
		when "0011101010101" => data_out <= rom_array(1877);
		when "0011101010110" => data_out <= rom_array(1878);
		when "0011101010111" => data_out <= rom_array(1879);
		when "0011101011000" => data_out <= rom_array(1880);
		when "0011101011001" => data_out <= rom_array(1881);
		when "0011101011010" => data_out <= rom_array(1882);
		when "0011101011011" => data_out <= rom_array(1883);
		when "0011101011100" => data_out <= rom_array(1884);
		when "0011101011101" => data_out <= rom_array(1885);
		when "0011101011110" => data_out <= rom_array(1886);
		when "0011101011111" => data_out <= rom_array(1887);
		when "0011101100000" => data_out <= rom_array(1888);
		when "0011101100001" => data_out <= rom_array(1889);
		when "0011101100010" => data_out <= rom_array(1890);
		when "0011101100011" => data_out <= rom_array(1891);
		when "0011101100100" => data_out <= rom_array(1892);
		when "0011101100101" => data_out <= rom_array(1893);
		when "0011101100110" => data_out <= rom_array(1894);
		when "0011101100111" => data_out <= rom_array(1895);
		when "0011101101000" => data_out <= rom_array(1896);
		when "0011101101001" => data_out <= rom_array(1897);
		when "0011101101010" => data_out <= rom_array(1898);
		when "0011101101011" => data_out <= rom_array(1899);
		when "0011101101100" => data_out <= rom_array(1900);
		when "0011101101101" => data_out <= rom_array(1901);
		when "0011101101110" => data_out <= rom_array(1902);
		when "0011101101111" => data_out <= rom_array(1903);
		when "0011101110000" => data_out <= rom_array(1904);
		when "0011101110001" => data_out <= rom_array(1905);
		when "0011101110010" => data_out <= rom_array(1906);
		when "0011101110011" => data_out <= rom_array(1907);
		when "0011101110100" => data_out <= rom_array(1908);
		when "0011101110101" => data_out <= rom_array(1909);
		when "0011101110110" => data_out <= rom_array(1910);
		when "0011101110111" => data_out <= rom_array(1911);
		when "0011101111000" => data_out <= rom_array(1912);
		when "0011101111001" => data_out <= rom_array(1913);
		when "0011101111010" => data_out <= rom_array(1914);
		when "0011101111011" => data_out <= rom_array(1915);
		when "0011101111100" => data_out <= rom_array(1916);
		when "0011101111101" => data_out <= rom_array(1917);
		when "0011101111110" => data_out <= rom_array(1918);
		when "0011101111111" => data_out <= rom_array(1919);
		when "0011110000000" => data_out <= rom_array(1920);
		when "0011110000001" => data_out <= rom_array(1921);
		when "0011110000010" => data_out <= rom_array(1922);
		when "0011110000011" => data_out <= rom_array(1923);
		when "0011110000100" => data_out <= rom_array(1924);
		when "0011110000101" => data_out <= rom_array(1925);
		when "0011110000110" => data_out <= rom_array(1926);
		when "0011110000111" => data_out <= rom_array(1927);
		when "0011110001000" => data_out <= rom_array(1928);
		when "0011110001001" => data_out <= rom_array(1929);
		when "0011110001010" => data_out <= rom_array(1930);
		when "0011110001011" => data_out <= rom_array(1931);
		when "0011110001100" => data_out <= rom_array(1932);
		when "0011110001101" => data_out <= rom_array(1933);
		when "0011110001110" => data_out <= rom_array(1934);
		when "0011110001111" => data_out <= rom_array(1935);
		when "0011110010000" => data_out <= rom_array(1936);
		when "0011110010001" => data_out <= rom_array(1937);
		when "0011110010010" => data_out <= rom_array(1938);
		when "0011110010011" => data_out <= rom_array(1939);
		when "0011110010100" => data_out <= rom_array(1940);
		when "0011110010101" => data_out <= rom_array(1941);
		when "0011110010110" => data_out <= rom_array(1942);
		when "0011110010111" => data_out <= rom_array(1943);
		when "0011110011000" => data_out <= rom_array(1944);
		when "0011110011001" => data_out <= rom_array(1945);
		when "0011110011010" => data_out <= rom_array(1946);
		when "0011110011011" => data_out <= rom_array(1947);
		when "0011110011100" => data_out <= rom_array(1948);
		when "0011110011101" => data_out <= rom_array(1949);
		when "0011110011110" => data_out <= rom_array(1950);
		when "0011110011111" => data_out <= rom_array(1951);
		when "0011110100000" => data_out <= rom_array(1952);
		when "0011110100001" => data_out <= rom_array(1953);
		when "0011110100010" => data_out <= rom_array(1954);
		when "0011110100011" => data_out <= rom_array(1955);
		when "0011110100100" => data_out <= rom_array(1956);
		when "0011110100101" => data_out <= rom_array(1957);
		when "0011110100110" => data_out <= rom_array(1958);
		when "0011110100111" => data_out <= rom_array(1959);
		when "0011110101000" => data_out <= rom_array(1960);
		when "0011110101001" => data_out <= rom_array(1961);
		when "0011110101010" => data_out <= rom_array(1962);
		when "0011110101011" => data_out <= rom_array(1963);
		when "0011110101100" => data_out <= rom_array(1964);
		when "0011110101101" => data_out <= rom_array(1965);
		when "0011110101110" => data_out <= rom_array(1966);
		when "0011110101111" => data_out <= rom_array(1967);
		when "0011110110000" => data_out <= rom_array(1968);
		when "0011110110001" => data_out <= rom_array(1969);
		when "0011110110010" => data_out <= rom_array(1970);
		when "0011110110011" => data_out <= rom_array(1971);
		when "0011110110100" => data_out <= rom_array(1972);
		when "0011110110101" => data_out <= rom_array(1973);
		when "0011110110110" => data_out <= rom_array(1974);
		when "0011110110111" => data_out <= rom_array(1975);
		when "0011110111000" => data_out <= rom_array(1976);
		when "0011110111001" => data_out <= rom_array(1977);
		when "0011110111010" => data_out <= rom_array(1978);
		when "0011110111011" => data_out <= rom_array(1979);
		when "0011110111100" => data_out <= rom_array(1980);
		when "0011110111101" => data_out <= rom_array(1981);
		when "0011110111110" => data_out <= rom_array(1982);
		when "0011110111111" => data_out <= rom_array(1983);
		when "0011111000000" => data_out <= rom_array(1984);
		when "0011111000001" => data_out <= rom_array(1985);
		when "0011111000010" => data_out <= rom_array(1986);
		when "0011111000011" => data_out <= rom_array(1987);
		when "0011111000100" => data_out <= rom_array(1988);
		when "0011111000101" => data_out <= rom_array(1989);
		when "0011111000110" => data_out <= rom_array(1990);
		when "0011111000111" => data_out <= rom_array(1991);
		when "0011111001000" => data_out <= rom_array(1992);
		when "0011111001001" => data_out <= rom_array(1993);
		when "0011111001010" => data_out <= rom_array(1994);
		when "0011111001011" => data_out <= rom_array(1995);
		when "0011111001100" => data_out <= rom_array(1996);
		when "0011111001101" => data_out <= rom_array(1997);
		when "0011111001110" => data_out <= rom_array(1998);
		when "0011111001111" => data_out <= rom_array(1999);
		when "0011111010000" => data_out <= rom_array(2000);
		when "0011111010001" => data_out <= rom_array(2001);
		when "0011111010010" => data_out <= rom_array(2002);
		when "0011111010011" => data_out <= rom_array(2003);
		when "0011111010100" => data_out <= rom_array(2004);
		when "0011111010101" => data_out <= rom_array(2005);
		when "0011111010110" => data_out <= rom_array(2006);
		when "0011111010111" => data_out <= rom_array(2007);
		when "0011111011000" => data_out <= rom_array(2008);
		when "0011111011001" => data_out <= rom_array(2009);
		when "0011111011010" => data_out <= rom_array(2010);
		when "0011111011011" => data_out <= rom_array(2011);
		when "0011111011100" => data_out <= rom_array(2012);
		when "0011111011101" => data_out <= rom_array(2013);
		when "0011111011110" => data_out <= rom_array(2014);
		when "0011111011111" => data_out <= rom_array(2015);
		when "0011111100000" => data_out <= rom_array(2016);
		when "0011111100001" => data_out <= rom_array(2017);
		when "0011111100010" => data_out <= rom_array(2018);
		when "0011111100011" => data_out <= rom_array(2019);
		when "0011111100100" => data_out <= rom_array(2020);
		when "0011111100101" => data_out <= rom_array(2021);
		when "0011111100110" => data_out <= rom_array(2022);
		when "0011111100111" => data_out <= rom_array(2023);
		when "0011111101000" => data_out <= rom_array(2024);
		when "0011111101001" => data_out <= rom_array(2025);
		when "0011111101010" => data_out <= rom_array(2026);
		when "0011111101011" => data_out <= rom_array(2027);
		when "0011111101100" => data_out <= rom_array(2028);
		when "0011111101101" => data_out <= rom_array(2029);
		when "0011111101110" => data_out <= rom_array(2030);
		when "0011111101111" => data_out <= rom_array(2031);
		when "0011111110000" => data_out <= rom_array(2032);
		when "0011111110001" => data_out <= rom_array(2033);
		when "0011111110010" => data_out <= rom_array(2034);
		when "0011111110011" => data_out <= rom_array(2035);
		when "0011111110100" => data_out <= rom_array(2036);
		when "0011111110101" => data_out <= rom_array(2037);
		when "0011111110110" => data_out <= rom_array(2038);
		when "0011111110111" => data_out <= rom_array(2039);
		when "0011111111000" => data_out <= rom_array(2040);
		when "0011111111001" => data_out <= rom_array(2041);
		when "0011111111010" => data_out <= rom_array(2042);
		when "0011111111011" => data_out <= rom_array(2043);
		when "0011111111100" => data_out <= rom_array(2044);
		when "0011111111101" => data_out <= rom_array(2045);
		when "0011111111110" => data_out <= rom_array(2046);
		when "0011111111111" => data_out <= rom_array(2047);
		when "0100000000000" => data_out <= rom_array(2048);
		when "0100000000001" => data_out <= rom_array(2049);
		when "0100000000010" => data_out <= rom_array(2050);
		when "0100000000011" => data_out <= rom_array(2051);
		when "0100000000100" => data_out <= rom_array(2052);
		when "0100000000101" => data_out <= rom_array(2053);
		when "0100000000110" => data_out <= rom_array(2054);
		when "0100000000111" => data_out <= rom_array(2055);
		when "0100000001000" => data_out <= rom_array(2056);
		when "0100000001001" => data_out <= rom_array(2057);
		when "0100000001010" => data_out <= rom_array(2058);
		when "0100000001011" => data_out <= rom_array(2059);
		when "0100000001100" => data_out <= rom_array(2060);
		when "0100000001101" => data_out <= rom_array(2061);
		when "0100000001110" => data_out <= rom_array(2062);
		when "0100000001111" => data_out <= rom_array(2063);
		when "0100000010000" => data_out <= rom_array(2064);
		when "0100000010001" => data_out <= rom_array(2065);
		when "0100000010010" => data_out <= rom_array(2066);
		when "0100000010011" => data_out <= rom_array(2067);
		when "0100000010100" => data_out <= rom_array(2068);
		when "0100000010101" => data_out <= rom_array(2069);
		when "0100000010110" => data_out <= rom_array(2070);
		when "0100000010111" => data_out <= rom_array(2071);
		when "0100000011000" => data_out <= rom_array(2072);
		when "0100000011001" => data_out <= rom_array(2073);
		when "0100000011010" => data_out <= rom_array(2074);
		when "0100000011011" => data_out <= rom_array(2075);
		when "0100000011100" => data_out <= rom_array(2076);
		when "0100000011101" => data_out <= rom_array(2077);
		when "0100000011110" => data_out <= rom_array(2078);
		when "0100000011111" => data_out <= rom_array(2079);
		when "0100000100000" => data_out <= rom_array(2080);
		when "0100000100001" => data_out <= rom_array(2081);
		when "0100000100010" => data_out <= rom_array(2082);
		when "0100000100011" => data_out <= rom_array(2083);
		when "0100000100100" => data_out <= rom_array(2084);
		when "0100000100101" => data_out <= rom_array(2085);
		when "0100000100110" => data_out <= rom_array(2086);
		when "0100000100111" => data_out <= rom_array(2087);
		when "0100000101000" => data_out <= rom_array(2088);
		when "0100000101001" => data_out <= rom_array(2089);
		when "0100000101010" => data_out <= rom_array(2090);
		when "0100000101011" => data_out <= rom_array(2091);
		when "0100000101100" => data_out <= rom_array(2092);
		when "0100000101101" => data_out <= rom_array(2093);
		when "0100000101110" => data_out <= rom_array(2094);
		when "0100000101111" => data_out <= rom_array(2095);
		when "0100000110000" => data_out <= rom_array(2096);
		when "0100000110001" => data_out <= rom_array(2097);
		when "0100000110010" => data_out <= rom_array(2098);
		when "0100000110011" => data_out <= rom_array(2099);
		when "0100000110100" => data_out <= rom_array(2100);
		when "0100000110101" => data_out <= rom_array(2101);
		when "0100000110110" => data_out <= rom_array(2102);
		when "0100000110111" => data_out <= rom_array(2103);
		when "0100000111000" => data_out <= rom_array(2104);
		when "0100000111001" => data_out <= rom_array(2105);
		when "0100000111010" => data_out <= rom_array(2106);
		when "0100000111011" => data_out <= rom_array(2107);
		when "0100000111100" => data_out <= rom_array(2108);
		when "0100000111101" => data_out <= rom_array(2109);
		when "0100000111110" => data_out <= rom_array(2110);
		when "0100000111111" => data_out <= rom_array(2111);
		when "0100001000000" => data_out <= rom_array(2112);
		when "0100001000001" => data_out <= rom_array(2113);
		when "0100001000010" => data_out <= rom_array(2114);
		when "0100001000011" => data_out <= rom_array(2115);
		when "0100001000100" => data_out <= rom_array(2116);
		when "0100001000101" => data_out <= rom_array(2117);
		when "0100001000110" => data_out <= rom_array(2118);
		when "0100001000111" => data_out <= rom_array(2119);
		when "0100001001000" => data_out <= rom_array(2120);
		when "0100001001001" => data_out <= rom_array(2121);
		when "0100001001010" => data_out <= rom_array(2122);
		when "0100001001011" => data_out <= rom_array(2123);
		when "0100001001100" => data_out <= rom_array(2124);
		when "0100001001101" => data_out <= rom_array(2125);
		when "0100001001110" => data_out <= rom_array(2126);
		when "0100001001111" => data_out <= rom_array(2127);
		when "0100001010000" => data_out <= rom_array(2128);
		when "0100001010001" => data_out <= rom_array(2129);
		when "0100001010010" => data_out <= rom_array(2130);
		when "0100001010011" => data_out <= rom_array(2131);
		when "0100001010100" => data_out <= rom_array(2132);
		when "0100001010101" => data_out <= rom_array(2133);
		when "0100001010110" => data_out <= rom_array(2134);
		when "0100001010111" => data_out <= rom_array(2135);
		when "0100001011000" => data_out <= rom_array(2136);
		when "0100001011001" => data_out <= rom_array(2137);
		when "0100001011010" => data_out <= rom_array(2138);
		when "0100001011011" => data_out <= rom_array(2139);
		when "0100001011100" => data_out <= rom_array(2140);
		when "0100001011101" => data_out <= rom_array(2141);
		when "0100001011110" => data_out <= rom_array(2142);
		when "0100001011111" => data_out <= rom_array(2143);
		when "0100001100000" => data_out <= rom_array(2144);
		when "0100001100001" => data_out <= rom_array(2145);
		when "0100001100010" => data_out <= rom_array(2146);
		when "0100001100011" => data_out <= rom_array(2147);
		when "0100001100100" => data_out <= rom_array(2148);
		when "0100001100101" => data_out <= rom_array(2149);
		when "0100001100110" => data_out <= rom_array(2150);
		when "0100001100111" => data_out <= rom_array(2151);
		when "0100001101000" => data_out <= rom_array(2152);
		when "0100001101001" => data_out <= rom_array(2153);
		when "0100001101010" => data_out <= rom_array(2154);
		when "0100001101011" => data_out <= rom_array(2155);
		when "0100001101100" => data_out <= rom_array(2156);
		when "0100001101101" => data_out <= rom_array(2157);
		when "0100001101110" => data_out <= rom_array(2158);
		when "0100001101111" => data_out <= rom_array(2159);
		when "0100001110000" => data_out <= rom_array(2160);
		when "0100001110001" => data_out <= rom_array(2161);
		when "0100001110010" => data_out <= rom_array(2162);
		when "0100001110011" => data_out <= rom_array(2163);
		when "0100001110100" => data_out <= rom_array(2164);
		when "0100001110101" => data_out <= rom_array(2165);
		when "0100001110110" => data_out <= rom_array(2166);
		when "0100001110111" => data_out <= rom_array(2167);
		when "0100001111000" => data_out <= rom_array(2168);
		when "0100001111001" => data_out <= rom_array(2169);
		when "0100001111010" => data_out <= rom_array(2170);
		when "0100001111011" => data_out <= rom_array(2171);
		when "0100001111100" => data_out <= rom_array(2172);
		when "0100001111101" => data_out <= rom_array(2173);
		when "0100001111110" => data_out <= rom_array(2174);
		when "0100001111111" => data_out <= rom_array(2175);
		when "0100010000000" => data_out <= rom_array(2176);
		when "0100010000001" => data_out <= rom_array(2177);
		when "0100010000010" => data_out <= rom_array(2178);
		when "0100010000011" => data_out <= rom_array(2179);
		when "0100010000100" => data_out <= rom_array(2180);
		when "0100010000101" => data_out <= rom_array(2181);
		when "0100010000110" => data_out <= rom_array(2182);
		when "0100010000111" => data_out <= rom_array(2183);
		when "0100010001000" => data_out <= rom_array(2184);
		when "0100010001001" => data_out <= rom_array(2185);
		when "0100010001010" => data_out <= rom_array(2186);
		when "0100010001011" => data_out <= rom_array(2187);
		when "0100010001100" => data_out <= rom_array(2188);
		when "0100010001101" => data_out <= rom_array(2189);
		when "0100010001110" => data_out <= rom_array(2190);
		when "0100010001111" => data_out <= rom_array(2191);
		when "0100010010000" => data_out <= rom_array(2192);
		when "0100010010001" => data_out <= rom_array(2193);
		when "0100010010010" => data_out <= rom_array(2194);
		when "0100010010011" => data_out <= rom_array(2195);
		when "0100010010100" => data_out <= rom_array(2196);
		when "0100010010101" => data_out <= rom_array(2197);
		when "0100010010110" => data_out <= rom_array(2198);
		when "0100010010111" => data_out <= rom_array(2199);
		when "0100010011000" => data_out <= rom_array(2200);
		when "0100010011001" => data_out <= rom_array(2201);
		when "0100010011010" => data_out <= rom_array(2202);
		when "0100010011011" => data_out <= rom_array(2203);
		when "0100010011100" => data_out <= rom_array(2204);
		when "0100010011101" => data_out <= rom_array(2205);
		when "0100010011110" => data_out <= rom_array(2206);
		when "0100010011111" => data_out <= rom_array(2207);
		when "0100010100000" => data_out <= rom_array(2208);
		when "0100010100001" => data_out <= rom_array(2209);
		when "0100010100010" => data_out <= rom_array(2210);
		when "0100010100011" => data_out <= rom_array(2211);
		when "0100010100100" => data_out <= rom_array(2212);
		when "0100010100101" => data_out <= rom_array(2213);
		when "0100010100110" => data_out <= rom_array(2214);
		when "0100010100111" => data_out <= rom_array(2215);
		when "0100010101000" => data_out <= rom_array(2216);
		when "0100010101001" => data_out <= rom_array(2217);
		when "0100010101010" => data_out <= rom_array(2218);
		when "0100010101011" => data_out <= rom_array(2219);
		when "0100010101100" => data_out <= rom_array(2220);
		when "0100010101101" => data_out <= rom_array(2221);
		when "0100010101110" => data_out <= rom_array(2222);
		when "0100010101111" => data_out <= rom_array(2223);
		when "0100010110000" => data_out <= rom_array(2224);
		when "0100010110001" => data_out <= rom_array(2225);
		when "0100010110010" => data_out <= rom_array(2226);
		when "0100010110011" => data_out <= rom_array(2227);
		when "0100010110100" => data_out <= rom_array(2228);
		when "0100010110101" => data_out <= rom_array(2229);
		when "0100010110110" => data_out <= rom_array(2230);
		when "0100010110111" => data_out <= rom_array(2231);
		when "0100010111000" => data_out <= rom_array(2232);
		when "0100010111001" => data_out <= rom_array(2233);
		when "0100010111010" => data_out <= rom_array(2234);
		when "0100010111011" => data_out <= rom_array(2235);
		when "0100010111100" => data_out <= rom_array(2236);
		when "0100010111101" => data_out <= rom_array(2237);
		when "0100010111110" => data_out <= rom_array(2238);
		when "0100010111111" => data_out <= rom_array(2239);
		when "0100011000000" => data_out <= rom_array(2240);
		when "0100011000001" => data_out <= rom_array(2241);
		when "0100011000010" => data_out <= rom_array(2242);
		when "0100011000011" => data_out <= rom_array(2243);
		when "0100011000100" => data_out <= rom_array(2244);
		when "0100011000101" => data_out <= rom_array(2245);
		when "0100011000110" => data_out <= rom_array(2246);
		when "0100011000111" => data_out <= rom_array(2247);
		when "0100011001000" => data_out <= rom_array(2248);
		when "0100011001001" => data_out <= rom_array(2249);
		when "0100011001010" => data_out <= rom_array(2250);
		when "0100011001011" => data_out <= rom_array(2251);
		when "0100011001100" => data_out <= rom_array(2252);
		when "0100011001101" => data_out <= rom_array(2253);
		when "0100011001110" => data_out <= rom_array(2254);
		when "0100011001111" => data_out <= rom_array(2255);
		when "0100011010000" => data_out <= rom_array(2256);
		when "0100011010001" => data_out <= rom_array(2257);
		when "0100011010010" => data_out <= rom_array(2258);
		when "0100011010011" => data_out <= rom_array(2259);
		when "0100011010100" => data_out <= rom_array(2260);
		when "0100011010101" => data_out <= rom_array(2261);
		when "0100011010110" => data_out <= rom_array(2262);
		when "0100011010111" => data_out <= rom_array(2263);
		when "0100011011000" => data_out <= rom_array(2264);
		when "0100011011001" => data_out <= rom_array(2265);
		when "0100011011010" => data_out <= rom_array(2266);
		when "0100011011011" => data_out <= rom_array(2267);
		when "0100011011100" => data_out <= rom_array(2268);
		when "0100011011101" => data_out <= rom_array(2269);
		when "0100011011110" => data_out <= rom_array(2270);
		when "0100011011111" => data_out <= rom_array(2271);
		when "0100011100000" => data_out <= rom_array(2272);
		when "0100011100001" => data_out <= rom_array(2273);
		when "0100011100010" => data_out <= rom_array(2274);
		when "0100011100011" => data_out <= rom_array(2275);
		when "0100011100100" => data_out <= rom_array(2276);
		when "0100011100101" => data_out <= rom_array(2277);
		when "0100011100110" => data_out <= rom_array(2278);
		when "0100011100111" => data_out <= rom_array(2279);
		when "0100011101000" => data_out <= rom_array(2280);
		when "0100011101001" => data_out <= rom_array(2281);
		when "0100011101010" => data_out <= rom_array(2282);
		when "0100011101011" => data_out <= rom_array(2283);
		when "0100011101100" => data_out <= rom_array(2284);
		when "0100011101101" => data_out <= rom_array(2285);
		when "0100011101110" => data_out <= rom_array(2286);
		when "0100011101111" => data_out <= rom_array(2287);
		when "0100011110000" => data_out <= rom_array(2288);
		when "0100011110001" => data_out <= rom_array(2289);
		when "0100011110010" => data_out <= rom_array(2290);
		when "0100011110011" => data_out <= rom_array(2291);
		when "0100011110100" => data_out <= rom_array(2292);
		when "0100011110101" => data_out <= rom_array(2293);
		when "0100011110110" => data_out <= rom_array(2294);
		when "0100011110111" => data_out <= rom_array(2295);
		when "0100011111000" => data_out <= rom_array(2296);
		when "0100011111001" => data_out <= rom_array(2297);
		when "0100011111010" => data_out <= rom_array(2298);
		when "0100011111011" => data_out <= rom_array(2299);
		when "0100011111100" => data_out <= rom_array(2300);
		when "0100011111101" => data_out <= rom_array(2301);
		when "0100011111110" => data_out <= rom_array(2302);
		when "0100011111111" => data_out <= rom_array(2303);
		when "0100100000000" => data_out <= rom_array(2304);
		when "0100100000001" => data_out <= rom_array(2305);
		when "0100100000010" => data_out <= rom_array(2306);
		when "0100100000011" => data_out <= rom_array(2307);
		when "0100100000100" => data_out <= rom_array(2308);
		when "0100100000101" => data_out <= rom_array(2309);
		when "0100100000110" => data_out <= rom_array(2310);
		when "0100100000111" => data_out <= rom_array(2311);
		when "0100100001000" => data_out <= rom_array(2312);
		when "0100100001001" => data_out <= rom_array(2313);
		when "0100100001010" => data_out <= rom_array(2314);
		when "0100100001011" => data_out <= rom_array(2315);
		when "0100100001100" => data_out <= rom_array(2316);
		when "0100100001101" => data_out <= rom_array(2317);
		when "0100100001110" => data_out <= rom_array(2318);
		when "0100100001111" => data_out <= rom_array(2319);
		when "0100100010000" => data_out <= rom_array(2320);
		when "0100100010001" => data_out <= rom_array(2321);
		when "0100100010010" => data_out <= rom_array(2322);
		when "0100100010011" => data_out <= rom_array(2323);
		when "0100100010100" => data_out <= rom_array(2324);
		when "0100100010101" => data_out <= rom_array(2325);
		when "0100100010110" => data_out <= rom_array(2326);
		when "0100100010111" => data_out <= rom_array(2327);
		when "0100100011000" => data_out <= rom_array(2328);
		when "0100100011001" => data_out <= rom_array(2329);
		when "0100100011010" => data_out <= rom_array(2330);
		when "0100100011011" => data_out <= rom_array(2331);
		when "0100100011100" => data_out <= rom_array(2332);
		when "0100100011101" => data_out <= rom_array(2333);
		when "0100100011110" => data_out <= rom_array(2334);
		when "0100100011111" => data_out <= rom_array(2335);
		when "0100100100000" => data_out <= rom_array(2336);
		when "0100100100001" => data_out <= rom_array(2337);
		when "0100100100010" => data_out <= rom_array(2338);
		when "0100100100011" => data_out <= rom_array(2339);
		when "0100100100100" => data_out <= rom_array(2340);
		when "0100100100101" => data_out <= rom_array(2341);
		when "0100100100110" => data_out <= rom_array(2342);
		when "0100100100111" => data_out <= rom_array(2343);
		when "0100100101000" => data_out <= rom_array(2344);
		when "0100100101001" => data_out <= rom_array(2345);
		when "0100100101010" => data_out <= rom_array(2346);
		when "0100100101011" => data_out <= rom_array(2347);
		when "0100100101100" => data_out <= rom_array(2348);
		when "0100100101101" => data_out <= rom_array(2349);
		when "0100100101110" => data_out <= rom_array(2350);
		when "0100100101111" => data_out <= rom_array(2351);
		when "0100100110000" => data_out <= rom_array(2352);
		when "0100100110001" => data_out <= rom_array(2353);
		when "0100100110010" => data_out <= rom_array(2354);
		when "0100100110011" => data_out <= rom_array(2355);
		when "0100100110100" => data_out <= rom_array(2356);
		when "0100100110101" => data_out <= rom_array(2357);
		when "0100100110110" => data_out <= rom_array(2358);
		when "0100100110111" => data_out <= rom_array(2359);
		when "0100100111000" => data_out <= rom_array(2360);
		when "0100100111001" => data_out <= rom_array(2361);
		when "0100100111010" => data_out <= rom_array(2362);
		when "0100100111011" => data_out <= rom_array(2363);
		when "0100100111100" => data_out <= rom_array(2364);
		when "0100100111101" => data_out <= rom_array(2365);
		when "0100100111110" => data_out <= rom_array(2366);
		when "0100100111111" => data_out <= rom_array(2367);
		when "0100101000000" => data_out <= rom_array(2368);
		when "0100101000001" => data_out <= rom_array(2369);
		when "0100101000010" => data_out <= rom_array(2370);
		when "0100101000011" => data_out <= rom_array(2371);
		when "0100101000100" => data_out <= rom_array(2372);
		when "0100101000101" => data_out <= rom_array(2373);
		when "0100101000110" => data_out <= rom_array(2374);
		when "0100101000111" => data_out <= rom_array(2375);
		when "0100101001000" => data_out <= rom_array(2376);
		when "0100101001001" => data_out <= rom_array(2377);
		when "0100101001010" => data_out <= rom_array(2378);
		when "0100101001011" => data_out <= rom_array(2379);
		when "0100101001100" => data_out <= rom_array(2380);
		when "0100101001101" => data_out <= rom_array(2381);
		when "0100101001110" => data_out <= rom_array(2382);
		when "0100101001111" => data_out <= rom_array(2383);
		when "0100101010000" => data_out <= rom_array(2384);
		when "0100101010001" => data_out <= rom_array(2385);
		when "0100101010010" => data_out <= rom_array(2386);
		when "0100101010011" => data_out <= rom_array(2387);
		when "0100101010100" => data_out <= rom_array(2388);
		when "0100101010101" => data_out <= rom_array(2389);
		when "0100101010110" => data_out <= rom_array(2390);
		when "0100101010111" => data_out <= rom_array(2391);
		when "0100101011000" => data_out <= rom_array(2392);
		when "0100101011001" => data_out <= rom_array(2393);
		when "0100101011010" => data_out <= rom_array(2394);
		when "0100101011011" => data_out <= rom_array(2395);
		when "0100101011100" => data_out <= rom_array(2396);
		when "0100101011101" => data_out <= rom_array(2397);
		when "0100101011110" => data_out <= rom_array(2398);
		when "0100101011111" => data_out <= rom_array(2399);
		when "0100101100000" => data_out <= rom_array(2400);
		when "0100101100001" => data_out <= rom_array(2401);
		when "0100101100010" => data_out <= rom_array(2402);
		when "0100101100011" => data_out <= rom_array(2403);
		when "0100101100100" => data_out <= rom_array(2404);
		when "0100101100101" => data_out <= rom_array(2405);
		when "0100101100110" => data_out <= rom_array(2406);
		when "0100101100111" => data_out <= rom_array(2407);
		when "0100101101000" => data_out <= rom_array(2408);
		when "0100101101001" => data_out <= rom_array(2409);
		when "0100101101010" => data_out <= rom_array(2410);
		when "0100101101011" => data_out <= rom_array(2411);
		when "0100101101100" => data_out <= rom_array(2412);
		when "0100101101101" => data_out <= rom_array(2413);
		when "0100101101110" => data_out <= rom_array(2414);
		when "0100101101111" => data_out <= rom_array(2415);
		when "0100101110000" => data_out <= rom_array(2416);
		when "0100101110001" => data_out <= rom_array(2417);
		when "0100101110010" => data_out <= rom_array(2418);
		when "0100101110011" => data_out <= rom_array(2419);
		when "0100101110100" => data_out <= rom_array(2420);
		when "0100101110101" => data_out <= rom_array(2421);
		when "0100101110110" => data_out <= rom_array(2422);
		when "0100101110111" => data_out <= rom_array(2423);
		when "0100101111000" => data_out <= rom_array(2424);
		when "0100101111001" => data_out <= rom_array(2425);
		when "0100101111010" => data_out <= rom_array(2426);
		when "0100101111011" => data_out <= rom_array(2427);
		when "0100101111100" => data_out <= rom_array(2428);
		when "0100101111101" => data_out <= rom_array(2429);
		when "0100101111110" => data_out <= rom_array(2430);
		when "0100101111111" => data_out <= rom_array(2431);
		when "0100110000000" => data_out <= rom_array(2432);
		when "0100110000001" => data_out <= rom_array(2433);
		when "0100110000010" => data_out <= rom_array(2434);
		when "0100110000011" => data_out <= rom_array(2435);
		when "0100110000100" => data_out <= rom_array(2436);
		when "0100110000101" => data_out <= rom_array(2437);
		when "0100110000110" => data_out <= rom_array(2438);
		when "0100110000111" => data_out <= rom_array(2439);
		when "0100110001000" => data_out <= rom_array(2440);
		when "0100110001001" => data_out <= rom_array(2441);
		when "0100110001010" => data_out <= rom_array(2442);
		when "0100110001011" => data_out <= rom_array(2443);
		when "0100110001100" => data_out <= rom_array(2444);
		when "0100110001101" => data_out <= rom_array(2445);
		when "0100110001110" => data_out <= rom_array(2446);
		when "0100110001111" => data_out <= rom_array(2447);
		when "0100110010000" => data_out <= rom_array(2448);
		when "0100110010001" => data_out <= rom_array(2449);
		when "0100110010010" => data_out <= rom_array(2450);
		when "0100110010011" => data_out <= rom_array(2451);
		when "0100110010100" => data_out <= rom_array(2452);
		when "0100110010101" => data_out <= rom_array(2453);
		when "0100110010110" => data_out <= rom_array(2454);
		when "0100110010111" => data_out <= rom_array(2455);
		when "0100110011000" => data_out <= rom_array(2456);
		when "0100110011001" => data_out <= rom_array(2457);
		when "0100110011010" => data_out <= rom_array(2458);
		when "0100110011011" => data_out <= rom_array(2459);
		when "0100110011100" => data_out <= rom_array(2460);
		when "0100110011101" => data_out <= rom_array(2461);
		when "0100110011110" => data_out <= rom_array(2462);
		when "0100110011111" => data_out <= rom_array(2463);
		when "0100110100000" => data_out <= rom_array(2464);
		when "0100110100001" => data_out <= rom_array(2465);
		when "0100110100010" => data_out <= rom_array(2466);
		when "0100110100011" => data_out <= rom_array(2467);
		when "0100110100100" => data_out <= rom_array(2468);
		when "0100110100101" => data_out <= rom_array(2469);
		when "0100110100110" => data_out <= rom_array(2470);
		when "0100110100111" => data_out <= rom_array(2471);
		when "0100110101000" => data_out <= rom_array(2472);
		when "0100110101001" => data_out <= rom_array(2473);
		when "0100110101010" => data_out <= rom_array(2474);
		when "0100110101011" => data_out <= rom_array(2475);
		when "0100110101100" => data_out <= rom_array(2476);
		when "0100110101101" => data_out <= rom_array(2477);
		when "0100110101110" => data_out <= rom_array(2478);
		when "0100110101111" => data_out <= rom_array(2479);
		when "0100110110000" => data_out <= rom_array(2480);
		when "0100110110001" => data_out <= rom_array(2481);
		when "0100110110010" => data_out <= rom_array(2482);
		when "0100110110011" => data_out <= rom_array(2483);
		when "0100110110100" => data_out <= rom_array(2484);
		when "0100110110101" => data_out <= rom_array(2485);
		when "0100110110110" => data_out <= rom_array(2486);
		when "0100110110111" => data_out <= rom_array(2487);
		when "0100110111000" => data_out <= rom_array(2488);
		when "0100110111001" => data_out <= rom_array(2489);
		when "0100110111010" => data_out <= rom_array(2490);
		when "0100110111011" => data_out <= rom_array(2491);
		when "0100110111100" => data_out <= rom_array(2492);
		when "0100110111101" => data_out <= rom_array(2493);
		when "0100110111110" => data_out <= rom_array(2494);
		when "0100110111111" => data_out <= rom_array(2495);
		when "0100111000000" => data_out <= rom_array(2496);
		when "0100111000001" => data_out <= rom_array(2497);
		when "0100111000010" => data_out <= rom_array(2498);
		when "0100111000011" => data_out <= rom_array(2499);
		when "0100111000100" => data_out <= rom_array(2500);
		when "0100111000101" => data_out <= rom_array(2501);
		when "0100111000110" => data_out <= rom_array(2502);
		when "0100111000111" => data_out <= rom_array(2503);
		when "0100111001000" => data_out <= rom_array(2504);
		when "0100111001001" => data_out <= rom_array(2505);
		when "0100111001010" => data_out <= rom_array(2506);
		when "0100111001011" => data_out <= rom_array(2507);
		when "0100111001100" => data_out <= rom_array(2508);
		when "0100111001101" => data_out <= rom_array(2509);
		when "0100111001110" => data_out <= rom_array(2510);
		when "0100111001111" => data_out <= rom_array(2511);
		when "0100111010000" => data_out <= rom_array(2512);
		when "0100111010001" => data_out <= rom_array(2513);
		when "0100111010010" => data_out <= rom_array(2514);
		when "0100111010011" => data_out <= rom_array(2515);
		when "0100111010100" => data_out <= rom_array(2516);
		when "0100111010101" => data_out <= rom_array(2517);
		when "0100111010110" => data_out <= rom_array(2518);
		when "0100111010111" => data_out <= rom_array(2519);
		when "0100111011000" => data_out <= rom_array(2520);
		when "0100111011001" => data_out <= rom_array(2521);
		when "0100111011010" => data_out <= rom_array(2522);
		when "0100111011011" => data_out <= rom_array(2523);
		when "0100111011100" => data_out <= rom_array(2524);
		when "0100111011101" => data_out <= rom_array(2525);
		when "0100111011110" => data_out <= rom_array(2526);
		when "0100111011111" => data_out <= rom_array(2527);
		when "0100111100000" => data_out <= rom_array(2528);
		when "0100111100001" => data_out <= rom_array(2529);
		when "0100111100010" => data_out <= rom_array(2530);
		when "0100111100011" => data_out <= rom_array(2531);
		when "0100111100100" => data_out <= rom_array(2532);
		when "0100111100101" => data_out <= rom_array(2533);
		when "0100111100110" => data_out <= rom_array(2534);
		when "0100111100111" => data_out <= rom_array(2535);
		when "0100111101000" => data_out <= rom_array(2536);
		when "0100111101001" => data_out <= rom_array(2537);
		when "0100111101010" => data_out <= rom_array(2538);
		when "0100111101011" => data_out <= rom_array(2539);
		when "0100111101100" => data_out <= rom_array(2540);
		when "0100111101101" => data_out <= rom_array(2541);
		when "0100111101110" => data_out <= rom_array(2542);
		when "0100111101111" => data_out <= rom_array(2543);
		when "0100111110000" => data_out <= rom_array(2544);
		when "0100111110001" => data_out <= rom_array(2545);
		when "0100111110010" => data_out <= rom_array(2546);
		when "0100111110011" => data_out <= rom_array(2547);
		when "0100111110100" => data_out <= rom_array(2548);
		when "0100111110101" => data_out <= rom_array(2549);
		when "0100111110110" => data_out <= rom_array(2550);
		when "0100111110111" => data_out <= rom_array(2551);
		when "0100111111000" => data_out <= rom_array(2552);
		when "0100111111001" => data_out <= rom_array(2553);
		when "0100111111010" => data_out <= rom_array(2554);
		when "0100111111011" => data_out <= rom_array(2555);
		when "0100111111100" => data_out <= rom_array(2556);
		when "0100111111101" => data_out <= rom_array(2557);
		when "0100111111110" => data_out <= rom_array(2558);
		when "0100111111111" => data_out <= rom_array(2559);
		when "0101000000000" => data_out <= rom_array(2560);
		when "0101000000001" => data_out <= rom_array(2561);
		when "0101000000010" => data_out <= rom_array(2562);
		when "0101000000011" => data_out <= rom_array(2563);
		when "0101000000100" => data_out <= rom_array(2564);
		when "0101000000101" => data_out <= rom_array(2565);
		when "0101000000110" => data_out <= rom_array(2566);
		when "0101000000111" => data_out <= rom_array(2567);
		when "0101000001000" => data_out <= rom_array(2568);
		when "0101000001001" => data_out <= rom_array(2569);
		when "0101000001010" => data_out <= rom_array(2570);
		when "0101000001011" => data_out <= rom_array(2571);
		when "0101000001100" => data_out <= rom_array(2572);
		when "0101000001101" => data_out <= rom_array(2573);
		when "0101000001110" => data_out <= rom_array(2574);
		when "0101000001111" => data_out <= rom_array(2575);
		when "0101000010000" => data_out <= rom_array(2576);
		when "0101000010001" => data_out <= rom_array(2577);
		when "0101000010010" => data_out <= rom_array(2578);
		when "0101000010011" => data_out <= rom_array(2579);
		when "0101000010100" => data_out <= rom_array(2580);
		when "0101000010101" => data_out <= rom_array(2581);
		when "0101000010110" => data_out <= rom_array(2582);
		when "0101000010111" => data_out <= rom_array(2583);
		when "0101000011000" => data_out <= rom_array(2584);
		when "0101000011001" => data_out <= rom_array(2585);
		when "0101000011010" => data_out <= rom_array(2586);
		when "0101000011011" => data_out <= rom_array(2587);
		when "0101000011100" => data_out <= rom_array(2588);
		when "0101000011101" => data_out <= rom_array(2589);
		when "0101000011110" => data_out <= rom_array(2590);
		when "0101000011111" => data_out <= rom_array(2591);
		when "0101000100000" => data_out <= rom_array(2592);
		when "0101000100001" => data_out <= rom_array(2593);
		when "0101000100010" => data_out <= rom_array(2594);
		when "0101000100011" => data_out <= rom_array(2595);
		when "0101000100100" => data_out <= rom_array(2596);
		when "0101000100101" => data_out <= rom_array(2597);
		when "0101000100110" => data_out <= rom_array(2598);
		when "0101000100111" => data_out <= rom_array(2599);
		when "0101000101000" => data_out <= rom_array(2600);
		when "0101000101001" => data_out <= rom_array(2601);
		when "0101000101010" => data_out <= rom_array(2602);
		when "0101000101011" => data_out <= rom_array(2603);
		when "0101000101100" => data_out <= rom_array(2604);
		when "0101000101101" => data_out <= rom_array(2605);
		when "0101000101110" => data_out <= rom_array(2606);
		when "0101000101111" => data_out <= rom_array(2607);
		when "0101000110000" => data_out <= rom_array(2608);
		when "0101000110001" => data_out <= rom_array(2609);
		when "0101000110010" => data_out <= rom_array(2610);
		when "0101000110011" => data_out <= rom_array(2611);
		when "0101000110100" => data_out <= rom_array(2612);
		when "0101000110101" => data_out <= rom_array(2613);
		when "0101000110110" => data_out <= rom_array(2614);
		when "0101000110111" => data_out <= rom_array(2615);
		when "0101000111000" => data_out <= rom_array(2616);
		when "0101000111001" => data_out <= rom_array(2617);
		when "0101000111010" => data_out <= rom_array(2618);
		when "0101000111011" => data_out <= rom_array(2619);
		when "0101000111100" => data_out <= rom_array(2620);
		when "0101000111101" => data_out <= rom_array(2621);
		when "0101000111110" => data_out <= rom_array(2622);
		when "0101000111111" => data_out <= rom_array(2623);
		when "0101001000000" => data_out <= rom_array(2624);
		when "0101001000001" => data_out <= rom_array(2625);
		when "0101001000010" => data_out <= rom_array(2626);
		when "0101001000011" => data_out <= rom_array(2627);
		when "0101001000100" => data_out <= rom_array(2628);
		when "0101001000101" => data_out <= rom_array(2629);
		when "0101001000110" => data_out <= rom_array(2630);
		when "0101001000111" => data_out <= rom_array(2631);
		when "0101001001000" => data_out <= rom_array(2632);
		when "0101001001001" => data_out <= rom_array(2633);
		when "0101001001010" => data_out <= rom_array(2634);
		when "0101001001011" => data_out <= rom_array(2635);
		when "0101001001100" => data_out <= rom_array(2636);
		when "0101001001101" => data_out <= rom_array(2637);
		when "0101001001110" => data_out <= rom_array(2638);
		when "0101001001111" => data_out <= rom_array(2639);
		when "0101001010000" => data_out <= rom_array(2640);
		when "0101001010001" => data_out <= rom_array(2641);
		when "0101001010010" => data_out <= rom_array(2642);
		when "0101001010011" => data_out <= rom_array(2643);
		when "0101001010100" => data_out <= rom_array(2644);
		when "0101001010101" => data_out <= rom_array(2645);
		when "0101001010110" => data_out <= rom_array(2646);
		when "0101001010111" => data_out <= rom_array(2647);
		when "0101001011000" => data_out <= rom_array(2648);
		when "0101001011001" => data_out <= rom_array(2649);
		when "0101001011010" => data_out <= rom_array(2650);
		when "0101001011011" => data_out <= rom_array(2651);
		when "0101001011100" => data_out <= rom_array(2652);
		when "0101001011101" => data_out <= rom_array(2653);
		when "0101001011110" => data_out <= rom_array(2654);
		when "0101001011111" => data_out <= rom_array(2655);
		when "0101001100000" => data_out <= rom_array(2656);
		when "0101001100001" => data_out <= rom_array(2657);
		when "0101001100010" => data_out <= rom_array(2658);
		when "0101001100011" => data_out <= rom_array(2659);
		when "0101001100100" => data_out <= rom_array(2660);
		when "0101001100101" => data_out <= rom_array(2661);
		when "0101001100110" => data_out <= rom_array(2662);
		when "0101001100111" => data_out <= rom_array(2663);
		when "0101001101000" => data_out <= rom_array(2664);
		when "0101001101001" => data_out <= rom_array(2665);
		when "0101001101010" => data_out <= rom_array(2666);
		when "0101001101011" => data_out <= rom_array(2667);
		when "0101001101100" => data_out <= rom_array(2668);
		when "0101001101101" => data_out <= rom_array(2669);
		when "0101001101110" => data_out <= rom_array(2670);
		when "0101001101111" => data_out <= rom_array(2671);
		when "0101001110000" => data_out <= rom_array(2672);
		when "0101001110001" => data_out <= rom_array(2673);
		when "0101001110010" => data_out <= rom_array(2674);
		when "0101001110011" => data_out <= rom_array(2675);
		when "0101001110100" => data_out <= rom_array(2676);
		when "0101001110101" => data_out <= rom_array(2677);
		when "0101001110110" => data_out <= rom_array(2678);
		when "0101001110111" => data_out <= rom_array(2679);
		when "0101001111000" => data_out <= rom_array(2680);
		when "0101001111001" => data_out <= rom_array(2681);
		when "0101001111010" => data_out <= rom_array(2682);
		when "0101001111011" => data_out <= rom_array(2683);
		when "0101001111100" => data_out <= rom_array(2684);
		when "0101001111101" => data_out <= rom_array(2685);
		when "0101001111110" => data_out <= rom_array(2686);
		when "0101001111111" => data_out <= rom_array(2687);
		when "0101010000000" => data_out <= rom_array(2688);
		when "0101010000001" => data_out <= rom_array(2689);
		when "0101010000010" => data_out <= rom_array(2690);
		when "0101010000011" => data_out <= rom_array(2691);
		when "0101010000100" => data_out <= rom_array(2692);
		when "0101010000101" => data_out <= rom_array(2693);
		when "0101010000110" => data_out <= rom_array(2694);
		when "0101010000111" => data_out <= rom_array(2695);
		when "0101010001000" => data_out <= rom_array(2696);
		when "0101010001001" => data_out <= rom_array(2697);
		when "0101010001010" => data_out <= rom_array(2698);
		when "0101010001011" => data_out <= rom_array(2699);
		when "0101010001100" => data_out <= rom_array(2700);
		when "0101010001101" => data_out <= rom_array(2701);
		when "0101010001110" => data_out <= rom_array(2702);
		when "0101010001111" => data_out <= rom_array(2703);
		when "0101010010000" => data_out <= rom_array(2704);
		when "0101010010001" => data_out <= rom_array(2705);
		when "0101010010010" => data_out <= rom_array(2706);
		when "0101010010011" => data_out <= rom_array(2707);
		when "0101010010100" => data_out <= rom_array(2708);
		when "0101010010101" => data_out <= rom_array(2709);
		when "0101010010110" => data_out <= rom_array(2710);
		when "0101010010111" => data_out <= rom_array(2711);
		when "0101010011000" => data_out <= rom_array(2712);
		when "0101010011001" => data_out <= rom_array(2713);
		when "0101010011010" => data_out <= rom_array(2714);
		when "0101010011011" => data_out <= rom_array(2715);
		when "0101010011100" => data_out <= rom_array(2716);
		when "0101010011101" => data_out <= rom_array(2717);
		when "0101010011110" => data_out <= rom_array(2718);
		when "0101010011111" => data_out <= rom_array(2719);
		when "0101010100000" => data_out <= rom_array(2720);
		when "0101010100001" => data_out <= rom_array(2721);
		when "0101010100010" => data_out <= rom_array(2722);
		when "0101010100011" => data_out <= rom_array(2723);
		when "0101010100100" => data_out <= rom_array(2724);
		when "0101010100101" => data_out <= rom_array(2725);
		when "0101010100110" => data_out <= rom_array(2726);
		when "0101010100111" => data_out <= rom_array(2727);
		when "0101010101000" => data_out <= rom_array(2728);
		when "0101010101001" => data_out <= rom_array(2729);
		when "0101010101010" => data_out <= rom_array(2730);
		when "0101010101011" => data_out <= rom_array(2731);
		when "0101010101100" => data_out <= rom_array(2732);
		when "0101010101101" => data_out <= rom_array(2733);
		when "0101010101110" => data_out <= rom_array(2734);
		when "0101010101111" => data_out <= rom_array(2735);
		when "0101010110000" => data_out <= rom_array(2736);
		when "0101010110001" => data_out <= rom_array(2737);
		when "0101010110010" => data_out <= rom_array(2738);
		when "0101010110011" => data_out <= rom_array(2739);
		when "0101010110100" => data_out <= rom_array(2740);
		when "0101010110101" => data_out <= rom_array(2741);
		when "0101010110110" => data_out <= rom_array(2742);
		when "0101010110111" => data_out <= rom_array(2743);
		when "0101010111000" => data_out <= rom_array(2744);
		when "0101010111001" => data_out <= rom_array(2745);
		when "0101010111010" => data_out <= rom_array(2746);
		when "0101010111011" => data_out <= rom_array(2747);
		when "0101010111100" => data_out <= rom_array(2748);
		when "0101010111101" => data_out <= rom_array(2749);
		when "0101010111110" => data_out <= rom_array(2750);
		when "0101010111111" => data_out <= rom_array(2751);
		when "0101011000000" => data_out <= rom_array(2752);
		when "0101011000001" => data_out <= rom_array(2753);
		when "0101011000010" => data_out <= rom_array(2754);
		when "0101011000011" => data_out <= rom_array(2755);
		when "0101011000100" => data_out <= rom_array(2756);
		when "0101011000101" => data_out <= rom_array(2757);
		when "0101011000110" => data_out <= rom_array(2758);
		when "0101011000111" => data_out <= rom_array(2759);
		when "0101011001000" => data_out <= rom_array(2760);
		when "0101011001001" => data_out <= rom_array(2761);
		when "0101011001010" => data_out <= rom_array(2762);
		when "0101011001011" => data_out <= rom_array(2763);
		when "0101011001100" => data_out <= rom_array(2764);
		when "0101011001101" => data_out <= rom_array(2765);
		when "0101011001110" => data_out <= rom_array(2766);
		when "0101011001111" => data_out <= rom_array(2767);
		when "0101011010000" => data_out <= rom_array(2768);
		when "0101011010001" => data_out <= rom_array(2769);
		when "0101011010010" => data_out <= rom_array(2770);
		when "0101011010011" => data_out <= rom_array(2771);
		when "0101011010100" => data_out <= rom_array(2772);
		when "0101011010101" => data_out <= rom_array(2773);
		when "0101011010110" => data_out <= rom_array(2774);
		when "0101011010111" => data_out <= rom_array(2775);
		when "0101011011000" => data_out <= rom_array(2776);
		when "0101011011001" => data_out <= rom_array(2777);
		when "0101011011010" => data_out <= rom_array(2778);
		when "0101011011011" => data_out <= rom_array(2779);
		when "0101011011100" => data_out <= rom_array(2780);
		when "0101011011101" => data_out <= rom_array(2781);
		when "0101011011110" => data_out <= rom_array(2782);
		when "0101011011111" => data_out <= rom_array(2783);
		when "0101011100000" => data_out <= rom_array(2784);
		when "0101011100001" => data_out <= rom_array(2785);
		when "0101011100010" => data_out <= rom_array(2786);
		when "0101011100011" => data_out <= rom_array(2787);
		when "0101011100100" => data_out <= rom_array(2788);
		when "0101011100101" => data_out <= rom_array(2789);
		when "0101011100110" => data_out <= rom_array(2790);
		when "0101011100111" => data_out <= rom_array(2791);
		when "0101011101000" => data_out <= rom_array(2792);
		when "0101011101001" => data_out <= rom_array(2793);
		when "0101011101010" => data_out <= rom_array(2794);
		when "0101011101011" => data_out <= rom_array(2795);
		when "0101011101100" => data_out <= rom_array(2796);
		when "0101011101101" => data_out <= rom_array(2797);
		when "0101011101110" => data_out <= rom_array(2798);
		when "0101011101111" => data_out <= rom_array(2799);
		when "0101011110000" => data_out <= rom_array(2800);
		when "0101011110001" => data_out <= rom_array(2801);
		when "0101011110010" => data_out <= rom_array(2802);
		when "0101011110011" => data_out <= rom_array(2803);
		when "0101011110100" => data_out <= rom_array(2804);
		when "0101011110101" => data_out <= rom_array(2805);
		when "0101011110110" => data_out <= rom_array(2806);
		when "0101011110111" => data_out <= rom_array(2807);
		when "0101011111000" => data_out <= rom_array(2808);
		when "0101011111001" => data_out <= rom_array(2809);
		when "0101011111010" => data_out <= rom_array(2810);
		when "0101011111011" => data_out <= rom_array(2811);
		when "0101011111100" => data_out <= rom_array(2812);
		when "0101011111101" => data_out <= rom_array(2813);
		when "0101011111110" => data_out <= rom_array(2814);
		when "0101011111111" => data_out <= rom_array(2815);
		when "0101100000000" => data_out <= rom_array(2816);
		when "0101100000001" => data_out <= rom_array(2817);
		when "0101100000010" => data_out <= rom_array(2818);
		when "0101100000011" => data_out <= rom_array(2819);
		when "0101100000100" => data_out <= rom_array(2820);
		when "0101100000101" => data_out <= rom_array(2821);
		when "0101100000110" => data_out <= rom_array(2822);
		when "0101100000111" => data_out <= rom_array(2823);
		when "0101100001000" => data_out <= rom_array(2824);
		when "0101100001001" => data_out <= rom_array(2825);
		when "0101100001010" => data_out <= rom_array(2826);
		when "0101100001011" => data_out <= rom_array(2827);
		when "0101100001100" => data_out <= rom_array(2828);
		when "0101100001101" => data_out <= rom_array(2829);
		when "0101100001110" => data_out <= rom_array(2830);
		when "0101100001111" => data_out <= rom_array(2831);
		when "0101100010000" => data_out <= rom_array(2832);
		when "0101100010001" => data_out <= rom_array(2833);
		when "0101100010010" => data_out <= rom_array(2834);
		when "0101100010011" => data_out <= rom_array(2835);
		when "0101100010100" => data_out <= rom_array(2836);
		when "0101100010101" => data_out <= rom_array(2837);
		when "0101100010110" => data_out <= rom_array(2838);
		when "0101100010111" => data_out <= rom_array(2839);
		when "0101100011000" => data_out <= rom_array(2840);
		when "0101100011001" => data_out <= rom_array(2841);
		when "0101100011010" => data_out <= rom_array(2842);
		when "0101100011011" => data_out <= rom_array(2843);
		when "0101100011100" => data_out <= rom_array(2844);
		when "0101100011101" => data_out <= rom_array(2845);
		when "0101100011110" => data_out <= rom_array(2846);
		when "0101100011111" => data_out <= rom_array(2847);
		when "0101100100000" => data_out <= rom_array(2848);
		when "0101100100001" => data_out <= rom_array(2849);
		when "0101100100010" => data_out <= rom_array(2850);
		when "0101100100011" => data_out <= rom_array(2851);
		when "0101100100100" => data_out <= rom_array(2852);
		when "0101100100101" => data_out <= rom_array(2853);
		when "0101100100110" => data_out <= rom_array(2854);
		when "0101100100111" => data_out <= rom_array(2855);
		when "0101100101000" => data_out <= rom_array(2856);
		when "0101100101001" => data_out <= rom_array(2857);
		when "0101100101010" => data_out <= rom_array(2858);
		when "0101100101011" => data_out <= rom_array(2859);
		when "0101100101100" => data_out <= rom_array(2860);
		when "0101100101101" => data_out <= rom_array(2861);
		when "0101100101110" => data_out <= rom_array(2862);
		when "0101100101111" => data_out <= rom_array(2863);
		when "0101100110000" => data_out <= rom_array(2864);
		when "0101100110001" => data_out <= rom_array(2865);
		when "0101100110010" => data_out <= rom_array(2866);
		when "0101100110011" => data_out <= rom_array(2867);
		when "0101100110100" => data_out <= rom_array(2868);
		when "0101100110101" => data_out <= rom_array(2869);
		when "0101100110110" => data_out <= rom_array(2870);
		when "0101100110111" => data_out <= rom_array(2871);
		when "0101100111000" => data_out <= rom_array(2872);
		when "0101100111001" => data_out <= rom_array(2873);
		when "0101100111010" => data_out <= rom_array(2874);
		when "0101100111011" => data_out <= rom_array(2875);
		when "0101100111100" => data_out <= rom_array(2876);
		when "0101100111101" => data_out <= rom_array(2877);
		when "0101100111110" => data_out <= rom_array(2878);
		when "0101100111111" => data_out <= rom_array(2879);
		when "0101101000000" => data_out <= rom_array(2880);
		when "0101101000001" => data_out <= rom_array(2881);
		when "0101101000010" => data_out <= rom_array(2882);
		when "0101101000011" => data_out <= rom_array(2883);
		when "0101101000100" => data_out <= rom_array(2884);
		when "0101101000101" => data_out <= rom_array(2885);
		when "0101101000110" => data_out <= rom_array(2886);
		when "0101101000111" => data_out <= rom_array(2887);
		when "0101101001000" => data_out <= rom_array(2888);
		when "0101101001001" => data_out <= rom_array(2889);
		when "0101101001010" => data_out <= rom_array(2890);
		when "0101101001011" => data_out <= rom_array(2891);
		when "0101101001100" => data_out <= rom_array(2892);
		when "0101101001101" => data_out <= rom_array(2893);
		when "0101101001110" => data_out <= rom_array(2894);
		when "0101101001111" => data_out <= rom_array(2895);
		when "0101101010000" => data_out <= rom_array(2896);
		when "0101101010001" => data_out <= rom_array(2897);
		when "0101101010010" => data_out <= rom_array(2898);
		when "0101101010011" => data_out <= rom_array(2899);
		when "0101101010100" => data_out <= rom_array(2900);
		when "0101101010101" => data_out <= rom_array(2901);
		when "0101101010110" => data_out <= rom_array(2902);
		when "0101101010111" => data_out <= rom_array(2903);
		when "0101101011000" => data_out <= rom_array(2904);
		when "0101101011001" => data_out <= rom_array(2905);
		when "0101101011010" => data_out <= rom_array(2906);
		when "0101101011011" => data_out <= rom_array(2907);
		when "0101101011100" => data_out <= rom_array(2908);
		when "0101101011101" => data_out <= rom_array(2909);
		when "0101101011110" => data_out <= rom_array(2910);
		when "0101101011111" => data_out <= rom_array(2911);
		when "0101101100000" => data_out <= rom_array(2912);
		when "0101101100001" => data_out <= rom_array(2913);
		when "0101101100010" => data_out <= rom_array(2914);
		when "0101101100011" => data_out <= rom_array(2915);
		when "0101101100100" => data_out <= rom_array(2916);
		when "0101101100101" => data_out <= rom_array(2917);
		when "0101101100110" => data_out <= rom_array(2918);
		when "0101101100111" => data_out <= rom_array(2919);
		when "0101101101000" => data_out <= rom_array(2920);
		when "0101101101001" => data_out <= rom_array(2921);
		when "0101101101010" => data_out <= rom_array(2922);
		when "0101101101011" => data_out <= rom_array(2923);
		when "0101101101100" => data_out <= rom_array(2924);
		when "0101101101101" => data_out <= rom_array(2925);
		when "0101101101110" => data_out <= rom_array(2926);
		when "0101101101111" => data_out <= rom_array(2927);
		when "0101101110000" => data_out <= rom_array(2928);
		when "0101101110001" => data_out <= rom_array(2929);
		when "0101101110010" => data_out <= rom_array(2930);
		when "0101101110011" => data_out <= rom_array(2931);
		when "0101101110100" => data_out <= rom_array(2932);
		when "0101101110101" => data_out <= rom_array(2933);
		when "0101101110110" => data_out <= rom_array(2934);
		when "0101101110111" => data_out <= rom_array(2935);
		when "0101101111000" => data_out <= rom_array(2936);
		when "0101101111001" => data_out <= rom_array(2937);
		when "0101101111010" => data_out <= rom_array(2938);
		when "0101101111011" => data_out <= rom_array(2939);
		when "0101101111100" => data_out <= rom_array(2940);
		when "0101101111101" => data_out <= rom_array(2941);
		when "0101101111110" => data_out <= rom_array(2942);
		when "0101101111111" => data_out <= rom_array(2943);
		when "0101110000000" => data_out <= rom_array(2944);
		when "0101110000001" => data_out <= rom_array(2945);
		when "0101110000010" => data_out <= rom_array(2946);
		when "0101110000011" => data_out <= rom_array(2947);
		when "0101110000100" => data_out <= rom_array(2948);
		when "0101110000101" => data_out <= rom_array(2949);
		when "0101110000110" => data_out <= rom_array(2950);
		when "0101110000111" => data_out <= rom_array(2951);
		when "0101110001000" => data_out <= rom_array(2952);
		when "0101110001001" => data_out <= rom_array(2953);
		when "0101110001010" => data_out <= rom_array(2954);
		when "0101110001011" => data_out <= rom_array(2955);
		when "0101110001100" => data_out <= rom_array(2956);
		when "0101110001101" => data_out <= rom_array(2957);
		when "0101110001110" => data_out <= rom_array(2958);
		when "0101110001111" => data_out <= rom_array(2959);
		when "0101110010000" => data_out <= rom_array(2960);
		when "0101110010001" => data_out <= rom_array(2961);
		when "0101110010010" => data_out <= rom_array(2962);
		when "0101110010011" => data_out <= rom_array(2963);
		when "0101110010100" => data_out <= rom_array(2964);
		when "0101110010101" => data_out <= rom_array(2965);
		when "0101110010110" => data_out <= rom_array(2966);
		when "0101110010111" => data_out <= rom_array(2967);
		when "0101110011000" => data_out <= rom_array(2968);
		when "0101110011001" => data_out <= rom_array(2969);
		when "0101110011010" => data_out <= rom_array(2970);
		when "0101110011011" => data_out <= rom_array(2971);
		when "0101110011100" => data_out <= rom_array(2972);
		when "0101110011101" => data_out <= rom_array(2973);
		when "0101110011110" => data_out <= rom_array(2974);
		when "0101110011111" => data_out <= rom_array(2975);
		when "0101110100000" => data_out <= rom_array(2976);
		when "0101110100001" => data_out <= rom_array(2977);
		when "0101110100010" => data_out <= rom_array(2978);
		when "0101110100011" => data_out <= rom_array(2979);
		when "0101110100100" => data_out <= rom_array(2980);
		when "0101110100101" => data_out <= rom_array(2981);
		when "0101110100110" => data_out <= rom_array(2982);
		when "0101110100111" => data_out <= rom_array(2983);
		when "0101110101000" => data_out <= rom_array(2984);
		when "0101110101001" => data_out <= rom_array(2985);
		when "0101110101010" => data_out <= rom_array(2986);
		when "0101110101011" => data_out <= rom_array(2987);
		when "0101110101100" => data_out <= rom_array(2988);
		when "0101110101101" => data_out <= rom_array(2989);
		when "0101110101110" => data_out <= rom_array(2990);
		when "0101110101111" => data_out <= rom_array(2991);
		when "0101110110000" => data_out <= rom_array(2992);
		when "0101110110001" => data_out <= rom_array(2993);
		when "0101110110010" => data_out <= rom_array(2994);
		when "0101110110011" => data_out <= rom_array(2995);
		when "0101110110100" => data_out <= rom_array(2996);
		when "0101110110101" => data_out <= rom_array(2997);
		when "0101110110110" => data_out <= rom_array(2998);
		when "0101110110111" => data_out <= rom_array(2999);
		when "0101110111000" => data_out <= rom_array(3000);
		when "0101110111001" => data_out <= rom_array(3001);
		when "0101110111010" => data_out <= rom_array(3002);
		when "0101110111011" => data_out <= rom_array(3003);
		when "0101110111100" => data_out <= rom_array(3004);
		when "0101110111101" => data_out <= rom_array(3005);
		when "0101110111110" => data_out <= rom_array(3006);
		when "0101110111111" => data_out <= rom_array(3007);
		when "0101111000000" => data_out <= rom_array(3008);
		when "0101111000001" => data_out <= rom_array(3009);
		when "0101111000010" => data_out <= rom_array(3010);
		when "0101111000011" => data_out <= rom_array(3011);
		when "0101111000100" => data_out <= rom_array(3012);
		when "0101111000101" => data_out <= rom_array(3013);
		when "0101111000110" => data_out <= rom_array(3014);
		when "0101111000111" => data_out <= rom_array(3015);
		when "0101111001000" => data_out <= rom_array(3016);
		when "0101111001001" => data_out <= rom_array(3017);
		when "0101111001010" => data_out <= rom_array(3018);
		when "0101111001011" => data_out <= rom_array(3019);
		when "0101111001100" => data_out <= rom_array(3020);
		when "0101111001101" => data_out <= rom_array(3021);
		when "0101111001110" => data_out <= rom_array(3022);
		when "0101111001111" => data_out <= rom_array(3023);
		when "0101111010000" => data_out <= rom_array(3024);
		when "0101111010001" => data_out <= rom_array(3025);
		when "0101111010010" => data_out <= rom_array(3026);
		when "0101111010011" => data_out <= rom_array(3027);
		when "0101111010100" => data_out <= rom_array(3028);
		when "0101111010101" => data_out <= rom_array(3029);
		when "0101111010110" => data_out <= rom_array(3030);
		when "0101111010111" => data_out <= rom_array(3031);
		when "0101111011000" => data_out <= rom_array(3032);
		when "0101111011001" => data_out <= rom_array(3033);
		when "0101111011010" => data_out <= rom_array(3034);
		when "0101111011011" => data_out <= rom_array(3035);
		when "0101111011100" => data_out <= rom_array(3036);
		when "0101111011101" => data_out <= rom_array(3037);
		when "0101111011110" => data_out <= rom_array(3038);
		when "0101111011111" => data_out <= rom_array(3039);
		when "0101111100000" => data_out <= rom_array(3040);
		when "0101111100001" => data_out <= rom_array(3041);
		when "0101111100010" => data_out <= rom_array(3042);
		when "0101111100011" => data_out <= rom_array(3043);
		when "0101111100100" => data_out <= rom_array(3044);
		when "0101111100101" => data_out <= rom_array(3045);
		when "0101111100110" => data_out <= rom_array(3046);
		when "0101111100111" => data_out <= rom_array(3047);
		when "0101111101000" => data_out <= rom_array(3048);
		when "0101111101001" => data_out <= rom_array(3049);
		when "0101111101010" => data_out <= rom_array(3050);
		when "0101111101011" => data_out <= rom_array(3051);
		when "0101111101100" => data_out <= rom_array(3052);
		when "0101111101101" => data_out <= rom_array(3053);
		when "0101111101110" => data_out <= rom_array(3054);
		when "0101111101111" => data_out <= rom_array(3055);
		when "0101111110000" => data_out <= rom_array(3056);
		when "0101111110001" => data_out <= rom_array(3057);
		when "0101111110010" => data_out <= rom_array(3058);
		when "0101111110011" => data_out <= rom_array(3059);
		when "0101111110100" => data_out <= rom_array(3060);
		when "0101111110101" => data_out <= rom_array(3061);
		when "0101111110110" => data_out <= rom_array(3062);
		when "0101111110111" => data_out <= rom_array(3063);
		when "0101111111000" => data_out <= rom_array(3064);
		when "0101111111001" => data_out <= rom_array(3065);
		when "0101111111010" => data_out <= rom_array(3066);
		when "0101111111011" => data_out <= rom_array(3067);
		when "0101111111100" => data_out <= rom_array(3068);
		when "0101111111101" => data_out <= rom_array(3069);
		when "0101111111110" => data_out <= rom_array(3070);
		when "0101111111111" => data_out <= rom_array(3071);
		when "0110000000000" => data_out <= rom_array(3072);
		when "0110000000001" => data_out <= rom_array(3073);
		when "0110000000010" => data_out <= rom_array(3074);
		when "0110000000011" => data_out <= rom_array(3075);
		when "0110000000100" => data_out <= rom_array(3076);
		when "0110000000101" => data_out <= rom_array(3077);
		when "0110000000110" => data_out <= rom_array(3078);
		when "0110000000111" => data_out <= rom_array(3079);
		when "0110000001000" => data_out <= rom_array(3080);
		when "0110000001001" => data_out <= rom_array(3081);
		when "0110000001010" => data_out <= rom_array(3082);
		when "0110000001011" => data_out <= rom_array(3083);
		when "0110000001100" => data_out <= rom_array(3084);
		when "0110000001101" => data_out <= rom_array(3085);
		when "0110000001110" => data_out <= rom_array(3086);
		when "0110000001111" => data_out <= rom_array(3087);
		when "0110000010000" => data_out <= rom_array(3088);
		when "0110000010001" => data_out <= rom_array(3089);
		when "0110000010010" => data_out <= rom_array(3090);
		when "0110000010011" => data_out <= rom_array(3091);
		when "0110000010100" => data_out <= rom_array(3092);
		when "0110000010101" => data_out <= rom_array(3093);
		when "0110000010110" => data_out <= rom_array(3094);
		when "0110000010111" => data_out <= rom_array(3095);
		when "0110000011000" => data_out <= rom_array(3096);
		when "0110000011001" => data_out <= rom_array(3097);
		when "0110000011010" => data_out <= rom_array(3098);
		when "0110000011011" => data_out <= rom_array(3099);
		when "0110000011100" => data_out <= rom_array(3100);
		when "0110000011101" => data_out <= rom_array(3101);
		when "0110000011110" => data_out <= rom_array(3102);
		when "0110000011111" => data_out <= rom_array(3103);
		when "0110000100000" => data_out <= rom_array(3104);
		when "0110000100001" => data_out <= rom_array(3105);
		when "0110000100010" => data_out <= rom_array(3106);
		when "0110000100011" => data_out <= rom_array(3107);
		when "0110000100100" => data_out <= rom_array(3108);
		when "0110000100101" => data_out <= rom_array(3109);
		when "0110000100110" => data_out <= rom_array(3110);
		when "0110000100111" => data_out <= rom_array(3111);
		when "0110000101000" => data_out <= rom_array(3112);
		when "0110000101001" => data_out <= rom_array(3113);
		when "0110000101010" => data_out <= rom_array(3114);
		when "0110000101011" => data_out <= rom_array(3115);
		when "0110000101100" => data_out <= rom_array(3116);
		when "0110000101101" => data_out <= rom_array(3117);
		when "0110000101110" => data_out <= rom_array(3118);
		when "0110000101111" => data_out <= rom_array(3119);
		when "0110000110000" => data_out <= rom_array(3120);
		when "0110000110001" => data_out <= rom_array(3121);
		when "0110000110010" => data_out <= rom_array(3122);
		when "0110000110011" => data_out <= rom_array(3123);
		when "0110000110100" => data_out <= rom_array(3124);
		when "0110000110101" => data_out <= rom_array(3125);
		when "0110000110110" => data_out <= rom_array(3126);
		when "0110000110111" => data_out <= rom_array(3127);
		when "0110000111000" => data_out <= rom_array(3128);
		when "0110000111001" => data_out <= rom_array(3129);
		when "0110000111010" => data_out <= rom_array(3130);
		when "0110000111011" => data_out <= rom_array(3131);
		when "0110000111100" => data_out <= rom_array(3132);
		when "0110000111101" => data_out <= rom_array(3133);
		when "0110000111110" => data_out <= rom_array(3134);
		when "0110000111111" => data_out <= rom_array(3135);
		when "0110001000000" => data_out <= rom_array(3136);
		when "0110001000001" => data_out <= rom_array(3137);
		when "0110001000010" => data_out <= rom_array(3138);
		when "0110001000011" => data_out <= rom_array(3139);
		when "0110001000100" => data_out <= rom_array(3140);
		when "0110001000101" => data_out <= rom_array(3141);
		when "0110001000110" => data_out <= rom_array(3142);
		when "0110001000111" => data_out <= rom_array(3143);
		when "0110001001000" => data_out <= rom_array(3144);
		when "0110001001001" => data_out <= rom_array(3145);
		when "0110001001010" => data_out <= rom_array(3146);
		when "0110001001011" => data_out <= rom_array(3147);
		when "0110001001100" => data_out <= rom_array(3148);
		when "0110001001101" => data_out <= rom_array(3149);
		when "0110001001110" => data_out <= rom_array(3150);
		when "0110001001111" => data_out <= rom_array(3151);
		when "0110001010000" => data_out <= rom_array(3152);
		when "0110001010001" => data_out <= rom_array(3153);
		when "0110001010010" => data_out <= rom_array(3154);
		when "0110001010011" => data_out <= rom_array(3155);
		when "0110001010100" => data_out <= rom_array(3156);
		when "0110001010101" => data_out <= rom_array(3157);
		when "0110001010110" => data_out <= rom_array(3158);
		when "0110001010111" => data_out <= rom_array(3159);
		when "0110001011000" => data_out <= rom_array(3160);
		when "0110001011001" => data_out <= rom_array(3161);
		when "0110001011010" => data_out <= rom_array(3162);
		when "0110001011011" => data_out <= rom_array(3163);
		when "0110001011100" => data_out <= rom_array(3164);
		when "0110001011101" => data_out <= rom_array(3165);
		when "0110001011110" => data_out <= rom_array(3166);
		when "0110001011111" => data_out <= rom_array(3167);
		when "0110001100000" => data_out <= rom_array(3168);
		when "0110001100001" => data_out <= rom_array(3169);
		when "0110001100010" => data_out <= rom_array(3170);
		when "0110001100011" => data_out <= rom_array(3171);
		when "0110001100100" => data_out <= rom_array(3172);
		when "0110001100101" => data_out <= rom_array(3173);
		when "0110001100110" => data_out <= rom_array(3174);
		when "0110001100111" => data_out <= rom_array(3175);
		when "0110001101000" => data_out <= rom_array(3176);
		when "0110001101001" => data_out <= rom_array(3177);
		when "0110001101010" => data_out <= rom_array(3178);
		when "0110001101011" => data_out <= rom_array(3179);
		when "0110001101100" => data_out <= rom_array(3180);
		when "0110001101101" => data_out <= rom_array(3181);
		when "0110001101110" => data_out <= rom_array(3182);
		when "0110001101111" => data_out <= rom_array(3183);
		when "0110001110000" => data_out <= rom_array(3184);
		when "0110001110001" => data_out <= rom_array(3185);
		when "0110001110010" => data_out <= rom_array(3186);
		when "0110001110011" => data_out <= rom_array(3187);
		when "0110001110100" => data_out <= rom_array(3188);
		when "0110001110101" => data_out <= rom_array(3189);
		when "0110001110110" => data_out <= rom_array(3190);
		when "0110001110111" => data_out <= rom_array(3191);
		when "0110001111000" => data_out <= rom_array(3192);
		when "0110001111001" => data_out <= rom_array(3193);
		when "0110001111010" => data_out <= rom_array(3194);
		when "0110001111011" => data_out <= rom_array(3195);
		when "0110001111100" => data_out <= rom_array(3196);
		when "0110001111101" => data_out <= rom_array(3197);
		when "0110001111110" => data_out <= rom_array(3198);
		when "0110001111111" => data_out <= rom_array(3199);
		when "0110010000000" => data_out <= rom_array(3200);
		when "0110010000001" => data_out <= rom_array(3201);
		when "0110010000010" => data_out <= rom_array(3202);
		when "0110010000011" => data_out <= rom_array(3203);
		when "0110010000100" => data_out <= rom_array(3204);
		when "0110010000101" => data_out <= rom_array(3205);
		when "0110010000110" => data_out <= rom_array(3206);
		when "0110010000111" => data_out <= rom_array(3207);
		when "0110010001000" => data_out <= rom_array(3208);
		when "0110010001001" => data_out <= rom_array(3209);
		when "0110010001010" => data_out <= rom_array(3210);
		when "0110010001011" => data_out <= rom_array(3211);
		when "0110010001100" => data_out <= rom_array(3212);
		when "0110010001101" => data_out <= rom_array(3213);
		when "0110010001110" => data_out <= rom_array(3214);
		when "0110010001111" => data_out <= rom_array(3215);
		when "0110010010000" => data_out <= rom_array(3216);
		when "0110010010001" => data_out <= rom_array(3217);
		when "0110010010010" => data_out <= rom_array(3218);
		when "0110010010011" => data_out <= rom_array(3219);
		when "0110010010100" => data_out <= rom_array(3220);
		when "0110010010101" => data_out <= rom_array(3221);
		when "0110010010110" => data_out <= rom_array(3222);
		when "0110010010111" => data_out <= rom_array(3223);
		when "0110010011000" => data_out <= rom_array(3224);
		when "0110010011001" => data_out <= rom_array(3225);
		when "0110010011010" => data_out <= rom_array(3226);
		when "0110010011011" => data_out <= rom_array(3227);
		when "0110010011100" => data_out <= rom_array(3228);
		when "0110010011101" => data_out <= rom_array(3229);
		when "0110010011110" => data_out <= rom_array(3230);
		when "0110010011111" => data_out <= rom_array(3231);
		when "0110010100000" => data_out <= rom_array(3232);
		when "0110010100001" => data_out <= rom_array(3233);
		when "0110010100010" => data_out <= rom_array(3234);
		when "0110010100011" => data_out <= rom_array(3235);
		when "0110010100100" => data_out <= rom_array(3236);
		when "0110010100101" => data_out <= rom_array(3237);
		when "0110010100110" => data_out <= rom_array(3238);
		when "0110010100111" => data_out <= rom_array(3239);
		when "0110010101000" => data_out <= rom_array(3240);
		when "0110010101001" => data_out <= rom_array(3241);
		when "0110010101010" => data_out <= rom_array(3242);
		when "0110010101011" => data_out <= rom_array(3243);
		when "0110010101100" => data_out <= rom_array(3244);
		when "0110010101101" => data_out <= rom_array(3245);
		when "0110010101110" => data_out <= rom_array(3246);
		when "0110010101111" => data_out <= rom_array(3247);
		when "0110010110000" => data_out <= rom_array(3248);
		when "0110010110001" => data_out <= rom_array(3249);
		when "0110010110010" => data_out <= rom_array(3250);
		when "0110010110011" => data_out <= rom_array(3251);
		when "0110010110100" => data_out <= rom_array(3252);
		when "0110010110101" => data_out <= rom_array(3253);
		when "0110010110110" => data_out <= rom_array(3254);
		when "0110010110111" => data_out <= rom_array(3255);
		when "0110010111000" => data_out <= rom_array(3256);
		when "0110010111001" => data_out <= rom_array(3257);
		when "0110010111010" => data_out <= rom_array(3258);
		when "0110010111011" => data_out <= rom_array(3259);
		when "0110010111100" => data_out <= rom_array(3260);
		when "0110010111101" => data_out <= rom_array(3261);
		when "0110010111110" => data_out <= rom_array(3262);
		when "0110010111111" => data_out <= rom_array(3263);
		when "0110011000000" => data_out <= rom_array(3264);
		when "0110011000001" => data_out <= rom_array(3265);
		when "0110011000010" => data_out <= rom_array(3266);
		when "0110011000011" => data_out <= rom_array(3267);
		when "0110011000100" => data_out <= rom_array(3268);
		when "0110011000101" => data_out <= rom_array(3269);
		when "0110011000110" => data_out <= rom_array(3270);
		when "0110011000111" => data_out <= rom_array(3271);
		when "0110011001000" => data_out <= rom_array(3272);
		when "0110011001001" => data_out <= rom_array(3273);
		when "0110011001010" => data_out <= rom_array(3274);
		when "0110011001011" => data_out <= rom_array(3275);
		when "0110011001100" => data_out <= rom_array(3276);
		when "0110011001101" => data_out <= rom_array(3277);
		when "0110011001110" => data_out <= rom_array(3278);
		when "0110011001111" => data_out <= rom_array(3279);
		when "0110011010000" => data_out <= rom_array(3280);
		when "0110011010001" => data_out <= rom_array(3281);
		when "0110011010010" => data_out <= rom_array(3282);
		when "0110011010011" => data_out <= rom_array(3283);
		when "0110011010100" => data_out <= rom_array(3284);
		when "0110011010101" => data_out <= rom_array(3285);
		when "0110011010110" => data_out <= rom_array(3286);
		when "0110011010111" => data_out <= rom_array(3287);
		when "0110011011000" => data_out <= rom_array(3288);
		when "0110011011001" => data_out <= rom_array(3289);
		when "0110011011010" => data_out <= rom_array(3290);
		when "0110011011011" => data_out <= rom_array(3291);
		when "0110011011100" => data_out <= rom_array(3292);
		when "0110011011101" => data_out <= rom_array(3293);
		when "0110011011110" => data_out <= rom_array(3294);
		when "0110011011111" => data_out <= rom_array(3295);
		when "0110011100000" => data_out <= rom_array(3296);
		when "0110011100001" => data_out <= rom_array(3297);
		when "0110011100010" => data_out <= rom_array(3298);
		when "0110011100011" => data_out <= rom_array(3299);
		when "0110011100100" => data_out <= rom_array(3300);
		when "0110011100101" => data_out <= rom_array(3301);
		when "0110011100110" => data_out <= rom_array(3302);
		when "0110011100111" => data_out <= rom_array(3303);
		when "0110011101000" => data_out <= rom_array(3304);
		when "0110011101001" => data_out <= rom_array(3305);
		when "0110011101010" => data_out <= rom_array(3306);
		when "0110011101011" => data_out <= rom_array(3307);
		when "0110011101100" => data_out <= rom_array(3308);
		when "0110011101101" => data_out <= rom_array(3309);
		when "0110011101110" => data_out <= rom_array(3310);
		when "0110011101111" => data_out <= rom_array(3311);
		when "0110011110000" => data_out <= rom_array(3312);
		when "0110011110001" => data_out <= rom_array(3313);
		when "0110011110010" => data_out <= rom_array(3314);
		when "0110011110011" => data_out <= rom_array(3315);
		when "0110011110100" => data_out <= rom_array(3316);
		when "0110011110101" => data_out <= rom_array(3317);
		when "0110011110110" => data_out <= rom_array(3318);
		when "0110011110111" => data_out <= rom_array(3319);
		when "0110011111000" => data_out <= rom_array(3320);
		when "0110011111001" => data_out <= rom_array(3321);
		when "0110011111010" => data_out <= rom_array(3322);
		when "0110011111011" => data_out <= rom_array(3323);
		when "0110011111100" => data_out <= rom_array(3324);
		when "0110011111101" => data_out <= rom_array(3325);
		when "0110011111110" => data_out <= rom_array(3326);
		when "0110011111111" => data_out <= rom_array(3327);
		when "0110100000000" => data_out <= rom_array(3328);
		when "0110100000001" => data_out <= rom_array(3329);
		when "0110100000010" => data_out <= rom_array(3330);
		when "0110100000011" => data_out <= rom_array(3331);
		when "0110100000100" => data_out <= rom_array(3332);
		when "0110100000101" => data_out <= rom_array(3333);
		when "0110100000110" => data_out <= rom_array(3334);
		when "0110100000111" => data_out <= rom_array(3335);
		when "0110100001000" => data_out <= rom_array(3336);
		when "0110100001001" => data_out <= rom_array(3337);
		when "0110100001010" => data_out <= rom_array(3338);
		when "0110100001011" => data_out <= rom_array(3339);
		when "0110100001100" => data_out <= rom_array(3340);
		when "0110100001101" => data_out <= rom_array(3341);
		when "0110100001110" => data_out <= rom_array(3342);
		when "0110100001111" => data_out <= rom_array(3343);
		when "0110100010000" => data_out <= rom_array(3344);
		when "0110100010001" => data_out <= rom_array(3345);
		when "0110100010010" => data_out <= rom_array(3346);
		when "0110100010011" => data_out <= rom_array(3347);
		when "0110100010100" => data_out <= rom_array(3348);
		when "0110100010101" => data_out <= rom_array(3349);
		when "0110100010110" => data_out <= rom_array(3350);
		when "0110100010111" => data_out <= rom_array(3351);
		when "0110100011000" => data_out <= rom_array(3352);
		when "0110100011001" => data_out <= rom_array(3353);
		when "0110100011010" => data_out <= rom_array(3354);
		when "0110100011011" => data_out <= rom_array(3355);
		when "0110100011100" => data_out <= rom_array(3356);
		when "0110100011101" => data_out <= rom_array(3357);
		when "0110100011110" => data_out <= rom_array(3358);
		when "0110100011111" => data_out <= rom_array(3359);
		when "0110100100000" => data_out <= rom_array(3360);
		when "0110100100001" => data_out <= rom_array(3361);
		when "0110100100010" => data_out <= rom_array(3362);
		when "0110100100011" => data_out <= rom_array(3363);
		when "0110100100100" => data_out <= rom_array(3364);
		when "0110100100101" => data_out <= rom_array(3365);
		when "0110100100110" => data_out <= rom_array(3366);
		when "0110100100111" => data_out <= rom_array(3367);
		when "0110100101000" => data_out <= rom_array(3368);
		when "0110100101001" => data_out <= rom_array(3369);
		when "0110100101010" => data_out <= rom_array(3370);
		when "0110100101011" => data_out <= rom_array(3371);
		when "0110100101100" => data_out <= rom_array(3372);
		when "0110100101101" => data_out <= rom_array(3373);
		when "0110100101110" => data_out <= rom_array(3374);
		when "0110100101111" => data_out <= rom_array(3375);
		when "0110100110000" => data_out <= rom_array(3376);
		when "0110100110001" => data_out <= rom_array(3377);
		when "0110100110010" => data_out <= rom_array(3378);
		when "0110100110011" => data_out <= rom_array(3379);
		when "0110100110100" => data_out <= rom_array(3380);
		when "0110100110101" => data_out <= rom_array(3381);
		when "0110100110110" => data_out <= rom_array(3382);
		when "0110100110111" => data_out <= rom_array(3383);
		when "0110100111000" => data_out <= rom_array(3384);
		when "0110100111001" => data_out <= rom_array(3385);
		when "0110100111010" => data_out <= rom_array(3386);
		when "0110100111011" => data_out <= rom_array(3387);
		when "0110100111100" => data_out <= rom_array(3388);
		when "0110100111101" => data_out <= rom_array(3389);
		when "0110100111110" => data_out <= rom_array(3390);
		when "0110100111111" => data_out <= rom_array(3391);
		when "0110101000000" => data_out <= rom_array(3392);
		when "0110101000001" => data_out <= rom_array(3393);
		when "0110101000010" => data_out <= rom_array(3394);
		when "0110101000011" => data_out <= rom_array(3395);
		when "0110101000100" => data_out <= rom_array(3396);
		when "0110101000101" => data_out <= rom_array(3397);
		when "0110101000110" => data_out <= rom_array(3398);
		when "0110101000111" => data_out <= rom_array(3399);
		when "0110101001000" => data_out <= rom_array(3400);
		when "0110101001001" => data_out <= rom_array(3401);
		when "0110101001010" => data_out <= rom_array(3402);
		when "0110101001011" => data_out <= rom_array(3403);
		when "0110101001100" => data_out <= rom_array(3404);
		when "0110101001101" => data_out <= rom_array(3405);
		when "0110101001110" => data_out <= rom_array(3406);
		when "0110101001111" => data_out <= rom_array(3407);
		when "0110101010000" => data_out <= rom_array(3408);
		when "0110101010001" => data_out <= rom_array(3409);
		when "0110101010010" => data_out <= rom_array(3410);
		when "0110101010011" => data_out <= rom_array(3411);
		when "0110101010100" => data_out <= rom_array(3412);
		when "0110101010101" => data_out <= rom_array(3413);
		when "0110101010110" => data_out <= rom_array(3414);
		when "0110101010111" => data_out <= rom_array(3415);
		when "0110101011000" => data_out <= rom_array(3416);
		when "0110101011001" => data_out <= rom_array(3417);
		when "0110101011010" => data_out <= rom_array(3418);
		when "0110101011011" => data_out <= rom_array(3419);
		when "0110101011100" => data_out <= rom_array(3420);
		when "0110101011101" => data_out <= rom_array(3421);
		when "0110101011110" => data_out <= rom_array(3422);
		when "0110101011111" => data_out <= rom_array(3423);
		when "0110101100000" => data_out <= rom_array(3424);
		when "0110101100001" => data_out <= rom_array(3425);
		when "0110101100010" => data_out <= rom_array(3426);
		when "0110101100011" => data_out <= rom_array(3427);
		when "0110101100100" => data_out <= rom_array(3428);
		when "0110101100101" => data_out <= rom_array(3429);
		when "0110101100110" => data_out <= rom_array(3430);
		when "0110101100111" => data_out <= rom_array(3431);
		when "0110101101000" => data_out <= rom_array(3432);
		when "0110101101001" => data_out <= rom_array(3433);
		when "0110101101010" => data_out <= rom_array(3434);
		when "0110101101011" => data_out <= rom_array(3435);
		when "0110101101100" => data_out <= rom_array(3436);
		when "0110101101101" => data_out <= rom_array(3437);
		when "0110101101110" => data_out <= rom_array(3438);
		when "0110101101111" => data_out <= rom_array(3439);
		when "0110101110000" => data_out <= rom_array(3440);
		when "0110101110001" => data_out <= rom_array(3441);
		when "0110101110010" => data_out <= rom_array(3442);
		when "0110101110011" => data_out <= rom_array(3443);
		when "0110101110100" => data_out <= rom_array(3444);
		when "0110101110101" => data_out <= rom_array(3445);
		when "0110101110110" => data_out <= rom_array(3446);
		when "0110101110111" => data_out <= rom_array(3447);
		when "0110101111000" => data_out <= rom_array(3448);
		when "0110101111001" => data_out <= rom_array(3449);
		when "0110101111010" => data_out <= rom_array(3450);
		when "0110101111011" => data_out <= rom_array(3451);
		when "0110101111100" => data_out <= rom_array(3452);
		when "0110101111101" => data_out <= rom_array(3453);
		when "0110101111110" => data_out <= rom_array(3454);
		when "0110101111111" => data_out <= rom_array(3455);
		when "0110110000000" => data_out <= rom_array(3456);
		when "0110110000001" => data_out <= rom_array(3457);
		when "0110110000010" => data_out <= rom_array(3458);
		when "0110110000011" => data_out <= rom_array(3459);
		when "0110110000100" => data_out <= rom_array(3460);
		when "0110110000101" => data_out <= rom_array(3461);
		when "0110110000110" => data_out <= rom_array(3462);
		when "0110110000111" => data_out <= rom_array(3463);
		when "0110110001000" => data_out <= rom_array(3464);
		when "0110110001001" => data_out <= rom_array(3465);
		when "0110110001010" => data_out <= rom_array(3466);
		when "0110110001011" => data_out <= rom_array(3467);
		when "0110110001100" => data_out <= rom_array(3468);
		when "0110110001101" => data_out <= rom_array(3469);
		when "0110110001110" => data_out <= rom_array(3470);
		when "0110110001111" => data_out <= rom_array(3471);
		when "0110110010000" => data_out <= rom_array(3472);
		when "0110110010001" => data_out <= rom_array(3473);
		when "0110110010010" => data_out <= rom_array(3474);
		when "0110110010011" => data_out <= rom_array(3475);
		when "0110110010100" => data_out <= rom_array(3476);
		when "0110110010101" => data_out <= rom_array(3477);
		when "0110110010110" => data_out <= rom_array(3478);
		when "0110110010111" => data_out <= rom_array(3479);
		when "0110110011000" => data_out <= rom_array(3480);
		when "0110110011001" => data_out <= rom_array(3481);
		when "0110110011010" => data_out <= rom_array(3482);
		when "0110110011011" => data_out <= rom_array(3483);
		when "0110110011100" => data_out <= rom_array(3484);
		when "0110110011101" => data_out <= rom_array(3485);
		when "0110110011110" => data_out <= rom_array(3486);
		when "0110110011111" => data_out <= rom_array(3487);
		when "0110110100000" => data_out <= rom_array(3488);
		when "0110110100001" => data_out <= rom_array(3489);
		when "0110110100010" => data_out <= rom_array(3490);
		when "0110110100011" => data_out <= rom_array(3491);
		when "0110110100100" => data_out <= rom_array(3492);
		when "0110110100101" => data_out <= rom_array(3493);
		when "0110110100110" => data_out <= rom_array(3494);
		when "0110110100111" => data_out <= rom_array(3495);
		when "0110110101000" => data_out <= rom_array(3496);
		when "0110110101001" => data_out <= rom_array(3497);
		when "0110110101010" => data_out <= rom_array(3498);
		when "0110110101011" => data_out <= rom_array(3499);
		when "0110110101100" => data_out <= rom_array(3500);
		when "0110110101101" => data_out <= rom_array(3501);
		when "0110110101110" => data_out <= rom_array(3502);
		when "0110110101111" => data_out <= rom_array(3503);
		when "0110110110000" => data_out <= rom_array(3504);
		when "0110110110001" => data_out <= rom_array(3505);
		when "0110110110010" => data_out <= rom_array(3506);
		when "0110110110011" => data_out <= rom_array(3507);
		when "0110110110100" => data_out <= rom_array(3508);
		when "0110110110101" => data_out <= rom_array(3509);
		when "0110110110110" => data_out <= rom_array(3510);
		when "0110110110111" => data_out <= rom_array(3511);
		when "0110110111000" => data_out <= rom_array(3512);
		when "0110110111001" => data_out <= rom_array(3513);
		when "0110110111010" => data_out <= rom_array(3514);
		when "0110110111011" => data_out <= rom_array(3515);
		when "0110110111100" => data_out <= rom_array(3516);
		when "0110110111101" => data_out <= rom_array(3517);
		when "0110110111110" => data_out <= rom_array(3518);
		when "0110110111111" => data_out <= rom_array(3519);
		when "0110111000000" => data_out <= rom_array(3520);
		when "0110111000001" => data_out <= rom_array(3521);
		when "0110111000010" => data_out <= rom_array(3522);
		when "0110111000011" => data_out <= rom_array(3523);
		when "0110111000100" => data_out <= rom_array(3524);
		when "0110111000101" => data_out <= rom_array(3525);
		when "0110111000110" => data_out <= rom_array(3526);
		when "0110111000111" => data_out <= rom_array(3527);
		when "0110111001000" => data_out <= rom_array(3528);
		when "0110111001001" => data_out <= rom_array(3529);
		when "0110111001010" => data_out <= rom_array(3530);
		when "0110111001011" => data_out <= rom_array(3531);
		when "0110111001100" => data_out <= rom_array(3532);
		when "0110111001101" => data_out <= rom_array(3533);
		when "0110111001110" => data_out <= rom_array(3534);
		when "0110111001111" => data_out <= rom_array(3535);
		when "0110111010000" => data_out <= rom_array(3536);
		when "0110111010001" => data_out <= rom_array(3537);
		when "0110111010010" => data_out <= rom_array(3538);
		when "0110111010011" => data_out <= rom_array(3539);
		when "0110111010100" => data_out <= rom_array(3540);
		when "0110111010101" => data_out <= rom_array(3541);
		when "0110111010110" => data_out <= rom_array(3542);
		when "0110111010111" => data_out <= rom_array(3543);
		when "0110111011000" => data_out <= rom_array(3544);
		when "0110111011001" => data_out <= rom_array(3545);
		when "0110111011010" => data_out <= rom_array(3546);
		when "0110111011011" => data_out <= rom_array(3547);
		when "0110111011100" => data_out <= rom_array(3548);
		when "0110111011101" => data_out <= rom_array(3549);
		when "0110111011110" => data_out <= rom_array(3550);
		when "0110111011111" => data_out <= rom_array(3551);
		when "0110111100000" => data_out <= rom_array(3552);
		when "0110111100001" => data_out <= rom_array(3553);
		when "0110111100010" => data_out <= rom_array(3554);
		when "0110111100011" => data_out <= rom_array(3555);
		when "0110111100100" => data_out <= rom_array(3556);
		when "0110111100101" => data_out <= rom_array(3557);
		when "0110111100110" => data_out <= rom_array(3558);
		when "0110111100111" => data_out <= rom_array(3559);
		when "0110111101000" => data_out <= rom_array(3560);
		when "0110111101001" => data_out <= rom_array(3561);
		when "0110111101010" => data_out <= rom_array(3562);
		when "0110111101011" => data_out <= rom_array(3563);
		when "0110111101100" => data_out <= rom_array(3564);
		when "0110111101101" => data_out <= rom_array(3565);
		when "0110111101110" => data_out <= rom_array(3566);
		when "0110111101111" => data_out <= rom_array(3567);
		when "0110111110000" => data_out <= rom_array(3568);
		when "0110111110001" => data_out <= rom_array(3569);
		when "0110111110010" => data_out <= rom_array(3570);
		when "0110111110011" => data_out <= rom_array(3571);
		when "0110111110100" => data_out <= rom_array(3572);
		when "0110111110101" => data_out <= rom_array(3573);
		when "0110111110110" => data_out <= rom_array(3574);
		when "0110111110111" => data_out <= rom_array(3575);
		when "0110111111000" => data_out <= rom_array(3576);
		when "0110111111001" => data_out <= rom_array(3577);
		when "0110111111010" => data_out <= rom_array(3578);
		when "0110111111011" => data_out <= rom_array(3579);
		when "0110111111100" => data_out <= rom_array(3580);
		when "0110111111101" => data_out <= rom_array(3581);
		when "0110111111110" => data_out <= rom_array(3582);
		when "0110111111111" => data_out <= rom_array(3583);
		when "0111000000000" => data_out <= rom_array(3584);
		when "0111000000001" => data_out <= rom_array(3585);
		when "0111000000010" => data_out <= rom_array(3586);
		when "0111000000011" => data_out <= rom_array(3587);
		when "0111000000100" => data_out <= rom_array(3588);
		when "0111000000101" => data_out <= rom_array(3589);
		when "0111000000110" => data_out <= rom_array(3590);
		when "0111000000111" => data_out <= rom_array(3591);
		when "0111000001000" => data_out <= rom_array(3592);
		when "0111000001001" => data_out <= rom_array(3593);
		when "0111000001010" => data_out <= rom_array(3594);
		when "0111000001011" => data_out <= rom_array(3595);
		when "0111000001100" => data_out <= rom_array(3596);
		when "0111000001101" => data_out <= rom_array(3597);
		when "0111000001110" => data_out <= rom_array(3598);
		when "0111000001111" => data_out <= rom_array(3599);
		when "0111000010000" => data_out <= rom_array(3600);
		when "0111000010001" => data_out <= rom_array(3601);
		when "0111000010010" => data_out <= rom_array(3602);
		when "0111000010011" => data_out <= rom_array(3603);
		when "0111000010100" => data_out <= rom_array(3604);
		when "0111000010101" => data_out <= rom_array(3605);
		when "0111000010110" => data_out <= rom_array(3606);
		when "0111000010111" => data_out <= rom_array(3607);
		when "0111000011000" => data_out <= rom_array(3608);
		when "0111000011001" => data_out <= rom_array(3609);
		when "0111000011010" => data_out <= rom_array(3610);
		when "0111000011011" => data_out <= rom_array(3611);
		when "0111000011100" => data_out <= rom_array(3612);
		when "0111000011101" => data_out <= rom_array(3613);
		when "0111000011110" => data_out <= rom_array(3614);
		when "0111000011111" => data_out <= rom_array(3615);
		when "0111000100000" => data_out <= rom_array(3616);
		when "0111000100001" => data_out <= rom_array(3617);
		when "0111000100010" => data_out <= rom_array(3618);
		when "0111000100011" => data_out <= rom_array(3619);
		when "0111000100100" => data_out <= rom_array(3620);
		when "0111000100101" => data_out <= rom_array(3621);
		when "0111000100110" => data_out <= rom_array(3622);
		when "0111000100111" => data_out <= rom_array(3623);
		when "0111000101000" => data_out <= rom_array(3624);
		when "0111000101001" => data_out <= rom_array(3625);
		when "0111000101010" => data_out <= rom_array(3626);
		when "0111000101011" => data_out <= rom_array(3627);
		when "0111000101100" => data_out <= rom_array(3628);
		when "0111000101101" => data_out <= rom_array(3629);
		when "0111000101110" => data_out <= rom_array(3630);
		when "0111000101111" => data_out <= rom_array(3631);
		when "0111000110000" => data_out <= rom_array(3632);
		when "0111000110001" => data_out <= rom_array(3633);
		when "0111000110010" => data_out <= rom_array(3634);
		when "0111000110011" => data_out <= rom_array(3635);
		when "0111000110100" => data_out <= rom_array(3636);
		when "0111000110101" => data_out <= rom_array(3637);
		when "0111000110110" => data_out <= rom_array(3638);
		when "0111000110111" => data_out <= rom_array(3639);
		when "0111000111000" => data_out <= rom_array(3640);
		when "0111000111001" => data_out <= rom_array(3641);
		when "0111000111010" => data_out <= rom_array(3642);
		when "0111000111011" => data_out <= rom_array(3643);
		when "0111000111100" => data_out <= rom_array(3644);
		when "0111000111101" => data_out <= rom_array(3645);
		when "0111000111110" => data_out <= rom_array(3646);
		when "0111000111111" => data_out <= rom_array(3647);
		when "0111001000000" => data_out <= rom_array(3648);
		when "0111001000001" => data_out <= rom_array(3649);
		when "0111001000010" => data_out <= rom_array(3650);
		when "0111001000011" => data_out <= rom_array(3651);
		when "0111001000100" => data_out <= rom_array(3652);
		when "0111001000101" => data_out <= rom_array(3653);
		when "0111001000110" => data_out <= rom_array(3654);
		when "0111001000111" => data_out <= rom_array(3655);
		when "0111001001000" => data_out <= rom_array(3656);
		when "0111001001001" => data_out <= rom_array(3657);
		when "0111001001010" => data_out <= rom_array(3658);
		when "0111001001011" => data_out <= rom_array(3659);
		when "0111001001100" => data_out <= rom_array(3660);
		when "0111001001101" => data_out <= rom_array(3661);
		when "0111001001110" => data_out <= rom_array(3662);
		when "0111001001111" => data_out <= rom_array(3663);
		when "0111001010000" => data_out <= rom_array(3664);
		when "0111001010001" => data_out <= rom_array(3665);
		when "0111001010010" => data_out <= rom_array(3666);
		when "0111001010011" => data_out <= rom_array(3667);
		when "0111001010100" => data_out <= rom_array(3668);
		when "0111001010101" => data_out <= rom_array(3669);
		when "0111001010110" => data_out <= rom_array(3670);
		when "0111001010111" => data_out <= rom_array(3671);
		when "0111001011000" => data_out <= rom_array(3672);
		when "0111001011001" => data_out <= rom_array(3673);
		when "0111001011010" => data_out <= rom_array(3674);
		when "0111001011011" => data_out <= rom_array(3675);
		when "0111001011100" => data_out <= rom_array(3676);
		when "0111001011101" => data_out <= rom_array(3677);
		when "0111001011110" => data_out <= rom_array(3678);
		when "0111001011111" => data_out <= rom_array(3679);
		when "0111001100000" => data_out <= rom_array(3680);
		when "0111001100001" => data_out <= rom_array(3681);
		when "0111001100010" => data_out <= rom_array(3682);
		when "0111001100011" => data_out <= rom_array(3683);
		when "0111001100100" => data_out <= rom_array(3684);
		when "0111001100101" => data_out <= rom_array(3685);
		when "0111001100110" => data_out <= rom_array(3686);
		when "0111001100111" => data_out <= rom_array(3687);
		when "0111001101000" => data_out <= rom_array(3688);
		when "0111001101001" => data_out <= rom_array(3689);
		when "0111001101010" => data_out <= rom_array(3690);
		when "0111001101011" => data_out <= rom_array(3691);
		when "0111001101100" => data_out <= rom_array(3692);
		when "0111001101101" => data_out <= rom_array(3693);
		when "0111001101110" => data_out <= rom_array(3694);
		when "0111001101111" => data_out <= rom_array(3695);
		when "0111001110000" => data_out <= rom_array(3696);
		when "0111001110001" => data_out <= rom_array(3697);
		when "0111001110010" => data_out <= rom_array(3698);
		when "0111001110011" => data_out <= rom_array(3699);
		when "0111001110100" => data_out <= rom_array(3700);
		when "0111001110101" => data_out <= rom_array(3701);
		when "0111001110110" => data_out <= rom_array(3702);
		when "0111001110111" => data_out <= rom_array(3703);
		when "0111001111000" => data_out <= rom_array(3704);
		when "0111001111001" => data_out <= rom_array(3705);
		when "0111001111010" => data_out <= rom_array(3706);
		when "0111001111011" => data_out <= rom_array(3707);
		when "0111001111100" => data_out <= rom_array(3708);
		when "0111001111101" => data_out <= rom_array(3709);
		when "0111001111110" => data_out <= rom_array(3710);
		when "0111001111111" => data_out <= rom_array(3711);
		when "0111010000000" => data_out <= rom_array(3712);
		when "0111010000001" => data_out <= rom_array(3713);
		when "0111010000010" => data_out <= rom_array(3714);
		when "0111010000011" => data_out <= rom_array(3715);
		when "0111010000100" => data_out <= rom_array(3716);
		when "0111010000101" => data_out <= rom_array(3717);
		when "0111010000110" => data_out <= rom_array(3718);
		when "0111010000111" => data_out <= rom_array(3719);
		when "0111010001000" => data_out <= rom_array(3720);
		when "0111010001001" => data_out <= rom_array(3721);
		when "0111010001010" => data_out <= rom_array(3722);
		when "0111010001011" => data_out <= rom_array(3723);
		when "0111010001100" => data_out <= rom_array(3724);
		when "0111010001101" => data_out <= rom_array(3725);
		when "0111010001110" => data_out <= rom_array(3726);
		when "0111010001111" => data_out <= rom_array(3727);
		when "0111010010000" => data_out <= rom_array(3728);
		when "0111010010001" => data_out <= rom_array(3729);
		when "0111010010010" => data_out <= rom_array(3730);
		when "0111010010011" => data_out <= rom_array(3731);
		when "0111010010100" => data_out <= rom_array(3732);
		when "0111010010101" => data_out <= rom_array(3733);
		when "0111010010110" => data_out <= rom_array(3734);
		when "0111010010111" => data_out <= rom_array(3735);
		when "0111010011000" => data_out <= rom_array(3736);
		when "0111010011001" => data_out <= rom_array(3737);
		when "0111010011010" => data_out <= rom_array(3738);
		when "0111010011011" => data_out <= rom_array(3739);
		when "0111010011100" => data_out <= rom_array(3740);
		when "0111010011101" => data_out <= rom_array(3741);
		when "0111010011110" => data_out <= rom_array(3742);
		when "0111010011111" => data_out <= rom_array(3743);
		when "0111010100000" => data_out <= rom_array(3744);
		when "0111010100001" => data_out <= rom_array(3745);
		when "0111010100010" => data_out <= rom_array(3746);
		when "0111010100011" => data_out <= rom_array(3747);
		when "0111010100100" => data_out <= rom_array(3748);
		when "0111010100101" => data_out <= rom_array(3749);
		when "0111010100110" => data_out <= rom_array(3750);
		when "0111010100111" => data_out <= rom_array(3751);
		when "0111010101000" => data_out <= rom_array(3752);
		when "0111010101001" => data_out <= rom_array(3753);
		when "0111010101010" => data_out <= rom_array(3754);
		when "0111010101011" => data_out <= rom_array(3755);
		when "0111010101100" => data_out <= rom_array(3756);
		when "0111010101101" => data_out <= rom_array(3757);
		when "0111010101110" => data_out <= rom_array(3758);
		when "0111010101111" => data_out <= rom_array(3759);
		when "0111010110000" => data_out <= rom_array(3760);
		when "0111010110001" => data_out <= rom_array(3761);
		when "0111010110010" => data_out <= rom_array(3762);
		when "0111010110011" => data_out <= rom_array(3763);
		when "0111010110100" => data_out <= rom_array(3764);
		when "0111010110101" => data_out <= rom_array(3765);
		when "0111010110110" => data_out <= rom_array(3766);
		when "0111010110111" => data_out <= rom_array(3767);
		when "0111010111000" => data_out <= rom_array(3768);
		when "0111010111001" => data_out <= rom_array(3769);
		when "0111010111010" => data_out <= rom_array(3770);
		when "0111010111011" => data_out <= rom_array(3771);
		when "0111010111100" => data_out <= rom_array(3772);
		when "0111010111101" => data_out <= rom_array(3773);
		when "0111010111110" => data_out <= rom_array(3774);
		when "0111010111111" => data_out <= rom_array(3775);
		when "0111011000000" => data_out <= rom_array(3776);
		when "0111011000001" => data_out <= rom_array(3777);
		when "0111011000010" => data_out <= rom_array(3778);
		when "0111011000011" => data_out <= rom_array(3779);
		when "0111011000100" => data_out <= rom_array(3780);
		when "0111011000101" => data_out <= rom_array(3781);
		when "0111011000110" => data_out <= rom_array(3782);
		when "0111011000111" => data_out <= rom_array(3783);
		when "0111011001000" => data_out <= rom_array(3784);
		when "0111011001001" => data_out <= rom_array(3785);
		when "0111011001010" => data_out <= rom_array(3786);
		when "0111011001011" => data_out <= rom_array(3787);
		when "0111011001100" => data_out <= rom_array(3788);
		when "0111011001101" => data_out <= rom_array(3789);
		when "0111011001110" => data_out <= rom_array(3790);
		when "0111011001111" => data_out <= rom_array(3791);
		when "0111011010000" => data_out <= rom_array(3792);
		when "0111011010001" => data_out <= rom_array(3793);
		when "0111011010010" => data_out <= rom_array(3794);
		when "0111011010011" => data_out <= rom_array(3795);
		when "0111011010100" => data_out <= rom_array(3796);
		when "0111011010101" => data_out <= rom_array(3797);
		when "0111011010110" => data_out <= rom_array(3798);
		when "0111011010111" => data_out <= rom_array(3799);
		when "0111011011000" => data_out <= rom_array(3800);
		when "0111011011001" => data_out <= rom_array(3801);
		when "0111011011010" => data_out <= rom_array(3802);
		when "0111011011011" => data_out <= rom_array(3803);
		when "0111011011100" => data_out <= rom_array(3804);
		when "0111011011101" => data_out <= rom_array(3805);
		when "0111011011110" => data_out <= rom_array(3806);
		when "0111011011111" => data_out <= rom_array(3807);
		when "0111011100000" => data_out <= rom_array(3808);
		when "0111011100001" => data_out <= rom_array(3809);
		when "0111011100010" => data_out <= rom_array(3810);
		when "0111011100011" => data_out <= rom_array(3811);
		when "0111011100100" => data_out <= rom_array(3812);
		when "0111011100101" => data_out <= rom_array(3813);
		when "0111011100110" => data_out <= rom_array(3814);
		when "0111011100111" => data_out <= rom_array(3815);
		when "0111011101000" => data_out <= rom_array(3816);
		when "0111011101001" => data_out <= rom_array(3817);
		when "0111011101010" => data_out <= rom_array(3818);
		when "0111011101011" => data_out <= rom_array(3819);
		when "0111011101100" => data_out <= rom_array(3820);
		when "0111011101101" => data_out <= rom_array(3821);
		when "0111011101110" => data_out <= rom_array(3822);
		when "0111011101111" => data_out <= rom_array(3823);
		when "0111011110000" => data_out <= rom_array(3824);
		when "0111011110001" => data_out <= rom_array(3825);
		when "0111011110010" => data_out <= rom_array(3826);
		when "0111011110011" => data_out <= rom_array(3827);
		when "0111011110100" => data_out <= rom_array(3828);
		when "0111011110101" => data_out <= rom_array(3829);
		when "0111011110110" => data_out <= rom_array(3830);
		when "0111011110111" => data_out <= rom_array(3831);
		when "0111011111000" => data_out <= rom_array(3832);
		when "0111011111001" => data_out <= rom_array(3833);
		when "0111011111010" => data_out <= rom_array(3834);
		when "0111011111011" => data_out <= rom_array(3835);
		when "0111011111100" => data_out <= rom_array(3836);
		when "0111011111101" => data_out <= rom_array(3837);
		when "0111011111110" => data_out <= rom_array(3838);
		when "0111011111111" => data_out <= rom_array(3839);
		when "0111100000000" => data_out <= rom_array(3840);
		when "0111100000001" => data_out <= rom_array(3841);
		when "0111100000010" => data_out <= rom_array(3842);
		when "0111100000011" => data_out <= rom_array(3843);
		when "0111100000100" => data_out <= rom_array(3844);
		when "0111100000101" => data_out <= rom_array(3845);
		when "0111100000110" => data_out <= rom_array(3846);
		when "0111100000111" => data_out <= rom_array(3847);
		when "0111100001000" => data_out <= rom_array(3848);
		when "0111100001001" => data_out <= rom_array(3849);
		when "0111100001010" => data_out <= rom_array(3850);
		when "0111100001011" => data_out <= rom_array(3851);
		when "0111100001100" => data_out <= rom_array(3852);
		when "0111100001101" => data_out <= rom_array(3853);
		when "0111100001110" => data_out <= rom_array(3854);
		when "0111100001111" => data_out <= rom_array(3855);
		when "0111100010000" => data_out <= rom_array(3856);
		when "0111100010001" => data_out <= rom_array(3857);
		when "0111100010010" => data_out <= rom_array(3858);
		when "0111100010011" => data_out <= rom_array(3859);
		when "0111100010100" => data_out <= rom_array(3860);
		when "0111100010101" => data_out <= rom_array(3861);
		when "0111100010110" => data_out <= rom_array(3862);
		when "0111100010111" => data_out <= rom_array(3863);
		when "0111100011000" => data_out <= rom_array(3864);
		when "0111100011001" => data_out <= rom_array(3865);
		when "0111100011010" => data_out <= rom_array(3866);
		when "0111100011011" => data_out <= rom_array(3867);
		when "0111100011100" => data_out <= rom_array(3868);
		when "0111100011101" => data_out <= rom_array(3869);
		when "0111100011110" => data_out <= rom_array(3870);
		when "0111100011111" => data_out <= rom_array(3871);
		when "0111100100000" => data_out <= rom_array(3872);
		when "0111100100001" => data_out <= rom_array(3873);
		when "0111100100010" => data_out <= rom_array(3874);
		when "0111100100011" => data_out <= rom_array(3875);
		when "0111100100100" => data_out <= rom_array(3876);
		when "0111100100101" => data_out <= rom_array(3877);
		when "0111100100110" => data_out <= rom_array(3878);
		when "0111100100111" => data_out <= rom_array(3879);
		when "0111100101000" => data_out <= rom_array(3880);
		when "0111100101001" => data_out <= rom_array(3881);
		when "0111100101010" => data_out <= rom_array(3882);
		when "0111100101011" => data_out <= rom_array(3883);
		when "0111100101100" => data_out <= rom_array(3884);
		when "0111100101101" => data_out <= rom_array(3885);
		when "0111100101110" => data_out <= rom_array(3886);
		when "0111100101111" => data_out <= rom_array(3887);
		when "0111100110000" => data_out <= rom_array(3888);
		when "0111100110001" => data_out <= rom_array(3889);
		when "0111100110010" => data_out <= rom_array(3890);
		when "0111100110011" => data_out <= rom_array(3891);
		when "0111100110100" => data_out <= rom_array(3892);
		when "0111100110101" => data_out <= rom_array(3893);
		when "0111100110110" => data_out <= rom_array(3894);
		when "0111100110111" => data_out <= rom_array(3895);
		when "0111100111000" => data_out <= rom_array(3896);
		when "0111100111001" => data_out <= rom_array(3897);
		when "0111100111010" => data_out <= rom_array(3898);
		when "0111100111011" => data_out <= rom_array(3899);
		when "0111100111100" => data_out <= rom_array(3900);
		when "0111100111101" => data_out <= rom_array(3901);
		when "0111100111110" => data_out <= rom_array(3902);
		when "0111100111111" => data_out <= rom_array(3903);
		when "0111101000000" => data_out <= rom_array(3904);
		when "0111101000001" => data_out <= rom_array(3905);
		when "0111101000010" => data_out <= rom_array(3906);
		when "0111101000011" => data_out <= rom_array(3907);
		when "0111101000100" => data_out <= rom_array(3908);
		when "0111101000101" => data_out <= rom_array(3909);
		when "0111101000110" => data_out <= rom_array(3910);
		when "0111101000111" => data_out <= rom_array(3911);
		when "0111101001000" => data_out <= rom_array(3912);
		when "0111101001001" => data_out <= rom_array(3913);
		when "0111101001010" => data_out <= rom_array(3914);
		when "0111101001011" => data_out <= rom_array(3915);
		when "0111101001100" => data_out <= rom_array(3916);
		when "0111101001101" => data_out <= rom_array(3917);
		when "0111101001110" => data_out <= rom_array(3918);
		when "0111101001111" => data_out <= rom_array(3919);
		when "0111101010000" => data_out <= rom_array(3920);
		when "0111101010001" => data_out <= rom_array(3921);
		when "0111101010010" => data_out <= rom_array(3922);
		when "0111101010011" => data_out <= rom_array(3923);
		when "0111101010100" => data_out <= rom_array(3924);
		when "0111101010101" => data_out <= rom_array(3925);
		when "0111101010110" => data_out <= rom_array(3926);
		when "0111101010111" => data_out <= rom_array(3927);
		when "0111101011000" => data_out <= rom_array(3928);
		when "0111101011001" => data_out <= rom_array(3929);
		when "0111101011010" => data_out <= rom_array(3930);
		when "0111101011011" => data_out <= rom_array(3931);
		when "0111101011100" => data_out <= rom_array(3932);
		when "0111101011101" => data_out <= rom_array(3933);
		when "0111101011110" => data_out <= rom_array(3934);
		when "0111101011111" => data_out <= rom_array(3935);
		when "0111101100000" => data_out <= rom_array(3936);
		when "0111101100001" => data_out <= rom_array(3937);
		when "0111101100010" => data_out <= rom_array(3938);
		when "0111101100011" => data_out <= rom_array(3939);
		when "0111101100100" => data_out <= rom_array(3940);
		when "0111101100101" => data_out <= rom_array(3941);
		when "0111101100110" => data_out <= rom_array(3942);
		when "0111101100111" => data_out <= rom_array(3943);
		when "0111101101000" => data_out <= rom_array(3944);
		when "0111101101001" => data_out <= rom_array(3945);
		when "0111101101010" => data_out <= rom_array(3946);
		when "0111101101011" => data_out <= rom_array(3947);
		when "0111101101100" => data_out <= rom_array(3948);
		when "0111101101101" => data_out <= rom_array(3949);
		when "0111101101110" => data_out <= rom_array(3950);
		when "0111101101111" => data_out <= rom_array(3951);
		when "0111101110000" => data_out <= rom_array(3952);
		when "0111101110001" => data_out <= rom_array(3953);
		when "0111101110010" => data_out <= rom_array(3954);
		when "0111101110011" => data_out <= rom_array(3955);
		when "0111101110100" => data_out <= rom_array(3956);
		when "0111101110101" => data_out <= rom_array(3957);
		when "0111101110110" => data_out <= rom_array(3958);
		when "0111101110111" => data_out <= rom_array(3959);
		when "0111101111000" => data_out <= rom_array(3960);
		when "0111101111001" => data_out <= rom_array(3961);
		when "0111101111010" => data_out <= rom_array(3962);
		when "0111101111011" => data_out <= rom_array(3963);
		when "0111101111100" => data_out <= rom_array(3964);
		when "0111101111101" => data_out <= rom_array(3965);
		when "0111101111110" => data_out <= rom_array(3966);
		when "0111101111111" => data_out <= rom_array(3967);
		when "0111110000000" => data_out <= rom_array(3968);
		when "0111110000001" => data_out <= rom_array(3969);
		when "0111110000010" => data_out <= rom_array(3970);
		when "0111110000011" => data_out <= rom_array(3971);
		when "0111110000100" => data_out <= rom_array(3972);
		when "0111110000101" => data_out <= rom_array(3973);
		when "0111110000110" => data_out <= rom_array(3974);
		when "0111110000111" => data_out <= rom_array(3975);
		when "0111110001000" => data_out <= rom_array(3976);
		when "0111110001001" => data_out <= rom_array(3977);
		when "0111110001010" => data_out <= rom_array(3978);
		when "0111110001011" => data_out <= rom_array(3979);
		when "0111110001100" => data_out <= rom_array(3980);
		when "0111110001101" => data_out <= rom_array(3981);
		when "0111110001110" => data_out <= rom_array(3982);
		when "0111110001111" => data_out <= rom_array(3983);
		when "0111110010000" => data_out <= rom_array(3984);
		when "0111110010001" => data_out <= rom_array(3985);
		when "0111110010010" => data_out <= rom_array(3986);
		when "0111110010011" => data_out <= rom_array(3987);
		when "0111110010100" => data_out <= rom_array(3988);
		when "0111110010101" => data_out <= rom_array(3989);
		when "0111110010110" => data_out <= rom_array(3990);
		when "0111110010111" => data_out <= rom_array(3991);
		when "0111110011000" => data_out <= rom_array(3992);
		when "0111110011001" => data_out <= rom_array(3993);
		when "0111110011010" => data_out <= rom_array(3994);
		when "0111110011011" => data_out <= rom_array(3995);
		when "0111110011100" => data_out <= rom_array(3996);
		when "0111110011101" => data_out <= rom_array(3997);
		when "0111110011110" => data_out <= rom_array(3998);
		when "0111110011111" => data_out <= rom_array(3999);
		when "0111110100000" => data_out <= rom_array(4000);
		when "0111110100001" => data_out <= rom_array(4001);
		when "0111110100010" => data_out <= rom_array(4002);
		when "0111110100011" => data_out <= rom_array(4003);
		when "0111110100100" => data_out <= rom_array(4004);
		when "0111110100101" => data_out <= rom_array(4005);
		when "0111110100110" => data_out <= rom_array(4006);
		when "0111110100111" => data_out <= rom_array(4007);
		when "0111110101000" => data_out <= rom_array(4008);
		when "0111110101001" => data_out <= rom_array(4009);
		when "0111110101010" => data_out <= rom_array(4010);
		when "0111110101011" => data_out <= rom_array(4011);
		when "0111110101100" => data_out <= rom_array(4012);
		when "0111110101101" => data_out <= rom_array(4013);
		when "0111110101110" => data_out <= rom_array(4014);
		when "0111110101111" => data_out <= rom_array(4015);
		when "0111110110000" => data_out <= rom_array(4016);
		when "0111110110001" => data_out <= rom_array(4017);
		when "0111110110010" => data_out <= rom_array(4018);
		when "0111110110011" => data_out <= rom_array(4019);
		when "0111110110100" => data_out <= rom_array(4020);
		when "0111110110101" => data_out <= rom_array(4021);
		when "0111110110110" => data_out <= rom_array(4022);
		when "0111110110111" => data_out <= rom_array(4023);
		when "0111110111000" => data_out <= rom_array(4024);
		when "0111110111001" => data_out <= rom_array(4025);
		when "0111110111010" => data_out <= rom_array(4026);
		when "0111110111011" => data_out <= rom_array(4027);
		when "0111110111100" => data_out <= rom_array(4028);
		when "0111110111101" => data_out <= rom_array(4029);
		when "0111110111110" => data_out <= rom_array(4030);
		when "0111110111111" => data_out <= rom_array(4031);
		when "0111111000000" => data_out <= rom_array(4032);
		when "0111111000001" => data_out <= rom_array(4033);
		when "0111111000010" => data_out <= rom_array(4034);
		when "0111111000011" => data_out <= rom_array(4035);
		when "0111111000100" => data_out <= rom_array(4036);
		when "0111111000101" => data_out <= rom_array(4037);
		when "0111111000110" => data_out <= rom_array(4038);
		when "0111111000111" => data_out <= rom_array(4039);
		when "0111111001000" => data_out <= rom_array(4040);
		when "0111111001001" => data_out <= rom_array(4041);
		when "0111111001010" => data_out <= rom_array(4042);
		when "0111111001011" => data_out <= rom_array(4043);
		when "0111111001100" => data_out <= rom_array(4044);
		when "0111111001101" => data_out <= rom_array(4045);
		when "0111111001110" => data_out <= rom_array(4046);
		when "0111111001111" => data_out <= rom_array(4047);
		when "0111111010000" => data_out <= rom_array(4048);
		when "0111111010001" => data_out <= rom_array(4049);
		when "0111111010010" => data_out <= rom_array(4050);
		when "0111111010011" => data_out <= rom_array(4051);
		when "0111111010100" => data_out <= rom_array(4052);
		when "0111111010101" => data_out <= rom_array(4053);
		when "0111111010110" => data_out <= rom_array(4054);
		when "0111111010111" => data_out <= rom_array(4055);
		when "0111111011000" => data_out <= rom_array(4056);
		when "0111111011001" => data_out <= rom_array(4057);
		when "0111111011010" => data_out <= rom_array(4058);
		when "0111111011011" => data_out <= rom_array(4059);
		when "0111111011100" => data_out <= rom_array(4060);
		when "0111111011101" => data_out <= rom_array(4061);
		when "0111111011110" => data_out <= rom_array(4062);
		when "0111111011111" => data_out <= rom_array(4063);
		when "0111111100000" => data_out <= rom_array(4064);
		when "0111111100001" => data_out <= rom_array(4065);
		when "0111111100010" => data_out <= rom_array(4066);
		when "0111111100011" => data_out <= rom_array(4067);
		when "0111111100100" => data_out <= rom_array(4068);
		when "0111111100101" => data_out <= rom_array(4069);
		when "0111111100110" => data_out <= rom_array(4070);
		when "0111111100111" => data_out <= rom_array(4071);
		when "0111111101000" => data_out <= rom_array(4072);
		when "0111111101001" => data_out <= rom_array(4073);
		when "0111111101010" => data_out <= rom_array(4074);
		when "0111111101011" => data_out <= rom_array(4075);
		when "0111111101100" => data_out <= rom_array(4076);
		when "0111111101101" => data_out <= rom_array(4077);
		when "0111111101110" => data_out <= rom_array(4078);
		when "0111111101111" => data_out <= rom_array(4079);
		when "0111111110000" => data_out <= rom_array(4080);
		when "0111111110001" => data_out <= rom_array(4081);
		when "0111111110010" => data_out <= rom_array(4082);
		when "0111111110011" => data_out <= rom_array(4083);
		when "0111111110100" => data_out <= rom_array(4084);
		when "0111111110101" => data_out <= rom_array(4085);
		when "0111111110110" => data_out <= rom_array(4086);
		when "0111111110111" => data_out <= rom_array(4087);
		when "0111111111000" => data_out <= rom_array(4088);
		when "0111111111001" => data_out <= rom_array(4089);
		when "0111111111010" => data_out <= rom_array(4090);
		when "0111111111011" => data_out <= rom_array(4091);
		when "0111111111100" => data_out <= rom_array(4092);
		when "0111111111101" => data_out <= rom_array(4093);
		when "0111111111110" => data_out <= rom_array(4094);
		when "0111111111111" => data_out <= rom_array(4095);
		when "1000000000000" => data_out <= rom_array(4096);
		when "1000000000001" => data_out <= rom_array(4097);
		when "1000000000010" => data_out <= rom_array(4098);
		when "1000000000011" => data_out <= rom_array(4099);
		when "1000000000100" => data_out <= rom_array(4100);
		when "1000000000101" => data_out <= rom_array(4101);
		when "1000000000110" => data_out <= rom_array(4102);
		when "1000000000111" => data_out <= rom_array(4103);
		when "1000000001000" => data_out <= rom_array(4104);
		when "1000000001001" => data_out <= rom_array(4105);
		when "1000000001010" => data_out <= rom_array(4106);
		when "1000000001011" => data_out <= rom_array(4107);
		when "1000000001100" => data_out <= rom_array(4108);
		when "1000000001101" => data_out <= rom_array(4109);
		when "1000000001110" => data_out <= rom_array(4110);
		when "1000000001111" => data_out <= rom_array(4111);
		when "1000000010000" => data_out <= rom_array(4112);
		when "1000000010001" => data_out <= rom_array(4113);
		when "1000000010010" => data_out <= rom_array(4114);
		when "1000000010011" => data_out <= rom_array(4115);
		when "1000000010100" => data_out <= rom_array(4116);
		when "1000000010101" => data_out <= rom_array(4117);
		when "1000000010110" => data_out <= rom_array(4118);
		when "1000000010111" => data_out <= rom_array(4119);
		when "1000000011000" => data_out <= rom_array(4120);
		when "1000000011001" => data_out <= rom_array(4121);
		when "1000000011010" => data_out <= rom_array(4122);
		when "1000000011011" => data_out <= rom_array(4123);
		when "1000000011100" => data_out <= rom_array(4124);
		when "1000000011101" => data_out <= rom_array(4125);
		when "1000000011110" => data_out <= rom_array(4126);
		when "1000000011111" => data_out <= rom_array(4127);
		when "1000000100000" => data_out <= rom_array(4128);
		when "1000000100001" => data_out <= rom_array(4129);
		when "1000000100010" => data_out <= rom_array(4130);
		when "1000000100011" => data_out <= rom_array(4131);
		when "1000000100100" => data_out <= rom_array(4132);
		when "1000000100101" => data_out <= rom_array(4133);
		when "1000000100110" => data_out <= rom_array(4134);
		when "1000000100111" => data_out <= rom_array(4135);
		when "1000000101000" => data_out <= rom_array(4136);
		when "1000000101001" => data_out <= rom_array(4137);
		when "1000000101010" => data_out <= rom_array(4138);
		when "1000000101011" => data_out <= rom_array(4139);
		when "1000000101100" => data_out <= rom_array(4140);
		when "1000000101101" => data_out <= rom_array(4141);
		when "1000000101110" => data_out <= rom_array(4142);
		when "1000000101111" => data_out <= rom_array(4143);
		when "1000000110000" => data_out <= rom_array(4144);
		when "1000000110001" => data_out <= rom_array(4145);
		when "1000000110010" => data_out <= rom_array(4146);
		when "1000000110011" => data_out <= rom_array(4147);
		when "1000000110100" => data_out <= rom_array(4148);
		when "1000000110101" => data_out <= rom_array(4149);
		when "1000000110110" => data_out <= rom_array(4150);
		when "1000000110111" => data_out <= rom_array(4151);
		when "1000000111000" => data_out <= rom_array(4152);
		when "1000000111001" => data_out <= rom_array(4153);
		when "1000000111010" => data_out <= rom_array(4154);
		when "1000000111011" => data_out <= rom_array(4155);
		when "1000000111100" => data_out <= rom_array(4156);
		when "1000000111101" => data_out <= rom_array(4157);
		when "1000000111110" => data_out <= rom_array(4158);
		when "1000000111111" => data_out <= rom_array(4159);
		when "1000001000000" => data_out <= rom_array(4160);
		when "1000001000001" => data_out <= rom_array(4161);
		when "1000001000010" => data_out <= rom_array(4162);
		when "1000001000011" => data_out <= rom_array(4163);
		when "1000001000100" => data_out <= rom_array(4164);
		when "1000001000101" => data_out <= rom_array(4165);
		when "1000001000110" => data_out <= rom_array(4166);
		when "1000001000111" => data_out <= rom_array(4167);
		when "1000001001000" => data_out <= rom_array(4168);
		when "1000001001001" => data_out <= rom_array(4169);
		when "1000001001010" => data_out <= rom_array(4170);
		when "1000001001011" => data_out <= rom_array(4171);
		when "1000001001100" => data_out <= rom_array(4172);
		when "1000001001101" => data_out <= rom_array(4173);
		when "1000001001110" => data_out <= rom_array(4174);
		when "1000001001111" => data_out <= rom_array(4175);
		when "1000001010000" => data_out <= rom_array(4176);
		when "1000001010001" => data_out <= rom_array(4177);
		when "1000001010010" => data_out <= rom_array(4178);
		when "1000001010011" => data_out <= rom_array(4179);
		when "1000001010100" => data_out <= rom_array(4180);
		when "1000001010101" => data_out <= rom_array(4181);
		when "1000001010110" => data_out <= rom_array(4182);
		when "1000001010111" => data_out <= rom_array(4183);
		when "1000001011000" => data_out <= rom_array(4184);
		when "1000001011001" => data_out <= rom_array(4185);
		when "1000001011010" => data_out <= rom_array(4186);
		when "1000001011011" => data_out <= rom_array(4187);
		when "1000001011100" => data_out <= rom_array(4188);
		when "1000001011101" => data_out <= rom_array(4189);
		when "1000001011110" => data_out <= rom_array(4190);
		when "1000001011111" => data_out <= rom_array(4191);
		when "1000001100000" => data_out <= rom_array(4192);
		when "1000001100001" => data_out <= rom_array(4193);
		when "1000001100010" => data_out <= rom_array(4194);
		when "1000001100011" => data_out <= rom_array(4195);
		when "1000001100100" => data_out <= rom_array(4196);
		when "1000001100101" => data_out <= rom_array(4197);
		when "1000001100110" => data_out <= rom_array(4198);
		when "1000001100111" => data_out <= rom_array(4199);
		when "1000001101000" => data_out <= rom_array(4200);
		when "1000001101001" => data_out <= rom_array(4201);
		when "1000001101010" => data_out <= rom_array(4202);
		when "1000001101011" => data_out <= rom_array(4203);
		when "1000001101100" => data_out <= rom_array(4204);
		when "1000001101101" => data_out <= rom_array(4205);
		when "1000001101110" => data_out <= rom_array(4206);
		when "1000001101111" => data_out <= rom_array(4207);
		when "1000001110000" => data_out <= rom_array(4208);
		when "1000001110001" => data_out <= rom_array(4209);
		when "1000001110010" => data_out <= rom_array(4210);
		when "1000001110011" => data_out <= rom_array(4211);
		when "1000001110100" => data_out <= rom_array(4212);
		when "1000001110101" => data_out <= rom_array(4213);
		when "1000001110110" => data_out <= rom_array(4214);
		when "1000001110111" => data_out <= rom_array(4215);
		when "1000001111000" => data_out <= rom_array(4216);
		when "1000001111001" => data_out <= rom_array(4217);
		when "1000001111010" => data_out <= rom_array(4218);
		when "1000001111011" => data_out <= rom_array(4219);
		when "1000001111100" => data_out <= rom_array(4220);
		when "1000001111101" => data_out <= rom_array(4221);
		when "1000001111110" => data_out <= rom_array(4222);
		when "1000001111111" => data_out <= rom_array(4223);
		when "1000010000000" => data_out <= rom_array(4224);
		when "1000010000001" => data_out <= rom_array(4225);
		when "1000010000010" => data_out <= rom_array(4226);
		when "1000010000011" => data_out <= rom_array(4227);
		when "1000010000100" => data_out <= rom_array(4228);
		when "1000010000101" => data_out <= rom_array(4229);
		when "1000010000110" => data_out <= rom_array(4230);
		when "1000010000111" => data_out <= rom_array(4231);
		when "1000010001000" => data_out <= rom_array(4232);
		when "1000010001001" => data_out <= rom_array(4233);
		when "1000010001010" => data_out <= rom_array(4234);
		when "1000010001011" => data_out <= rom_array(4235);
		when "1000010001100" => data_out <= rom_array(4236);
		when "1000010001101" => data_out <= rom_array(4237);
		when "1000010001110" => data_out <= rom_array(4238);
		when "1000010001111" => data_out <= rom_array(4239);
		when "1000010010000" => data_out <= rom_array(4240);
		when "1000010010001" => data_out <= rom_array(4241);
		when "1000010010010" => data_out <= rom_array(4242);
		when "1000010010011" => data_out <= rom_array(4243);
		when "1000010010100" => data_out <= rom_array(4244);
		when "1000010010101" => data_out <= rom_array(4245);
		when "1000010010110" => data_out <= rom_array(4246);
		when "1000010010111" => data_out <= rom_array(4247);
		when "1000010011000" => data_out <= rom_array(4248);
		when "1000010011001" => data_out <= rom_array(4249);
		when "1000010011010" => data_out <= rom_array(4250);
		when "1000010011011" => data_out <= rom_array(4251);
		when "1000010011100" => data_out <= rom_array(4252);
		when "1000010011101" => data_out <= rom_array(4253);
		when "1000010011110" => data_out <= rom_array(4254);
		when "1000010011111" => data_out <= rom_array(4255);
		when "1000010100000" => data_out <= rom_array(4256);
		when "1000010100001" => data_out <= rom_array(4257);
		when "1000010100010" => data_out <= rom_array(4258);
		when "1000010100011" => data_out <= rom_array(4259);
		when "1000010100100" => data_out <= rom_array(4260);
		when "1000010100101" => data_out <= rom_array(4261);
		when "1000010100110" => data_out <= rom_array(4262);
		when "1000010100111" => data_out <= rom_array(4263);
		when "1000010101000" => data_out <= rom_array(4264);
		when "1000010101001" => data_out <= rom_array(4265);
		when "1000010101010" => data_out <= rom_array(4266);
		when "1000010101011" => data_out <= rom_array(4267);
		when "1000010101100" => data_out <= rom_array(4268);
		when "1000010101101" => data_out <= rom_array(4269);
		when "1000010101110" => data_out <= rom_array(4270);
		when "1000010101111" => data_out <= rom_array(4271);
		when "1000010110000" => data_out <= rom_array(4272);
		when "1000010110001" => data_out <= rom_array(4273);
		when "1000010110010" => data_out <= rom_array(4274);
		when "1000010110011" => data_out <= rom_array(4275);
		when "1000010110100" => data_out <= rom_array(4276);
		when "1000010110101" => data_out <= rom_array(4277);
		when "1000010110110" => data_out <= rom_array(4278);
		when "1000010110111" => data_out <= rom_array(4279);
		when "1000010111000" => data_out <= rom_array(4280);
		when "1000010111001" => data_out <= rom_array(4281);
		when "1000010111010" => data_out <= rom_array(4282);
		when "1000010111011" => data_out <= rom_array(4283);
		when "1000010111100" => data_out <= rom_array(4284);
		when "1000010111101" => data_out <= rom_array(4285);
		when "1000010111110" => data_out <= rom_array(4286);
		when "1000010111111" => data_out <= rom_array(4287);
		when "1000011000000" => data_out <= rom_array(4288);
		when "1000011000001" => data_out <= rom_array(4289);
		when "1000011000010" => data_out <= rom_array(4290);
		when "1000011000011" => data_out <= rom_array(4291);
		when "1000011000100" => data_out <= rom_array(4292);
		when "1000011000101" => data_out <= rom_array(4293);
		when "1000011000110" => data_out <= rom_array(4294);
		when "1000011000111" => data_out <= rom_array(4295);
		when "1000011001000" => data_out <= rom_array(4296);
		when "1000011001001" => data_out <= rom_array(4297);
		when "1000011001010" => data_out <= rom_array(4298);
		when "1000011001011" => data_out <= rom_array(4299);
		when "1000011001100" => data_out <= rom_array(4300);
		when "1000011001101" => data_out <= rom_array(4301);
		when "1000011001110" => data_out <= rom_array(4302);
		when "1000011001111" => data_out <= rom_array(4303);
		when "1000011010000" => data_out <= rom_array(4304);
		when "1000011010001" => data_out <= rom_array(4305);
		when "1000011010010" => data_out <= rom_array(4306);
		when "1000011010011" => data_out <= rom_array(4307);
		when "1000011010100" => data_out <= rom_array(4308);
		when "1000011010101" => data_out <= rom_array(4309);
		when "1000011010110" => data_out <= rom_array(4310);
		when "1000011010111" => data_out <= rom_array(4311);
		when "1000011011000" => data_out <= rom_array(4312);
		when "1000011011001" => data_out <= rom_array(4313);
		when "1000011011010" => data_out <= rom_array(4314);
		when "1000011011011" => data_out <= rom_array(4315);
		when "1000011011100" => data_out <= rom_array(4316);
		when "1000011011101" => data_out <= rom_array(4317);
		when "1000011011110" => data_out <= rom_array(4318);
		when "1000011011111" => data_out <= rom_array(4319);
		when "1000011100000" => data_out <= rom_array(4320);
		when "1000011100001" => data_out <= rom_array(4321);
		when "1000011100010" => data_out <= rom_array(4322);
		when "1000011100011" => data_out <= rom_array(4323);
		when "1000011100100" => data_out <= rom_array(4324);
		when "1000011100101" => data_out <= rom_array(4325);
		when "1000011100110" => data_out <= rom_array(4326);
		when "1000011100111" => data_out <= rom_array(4327);
		when "1000011101000" => data_out <= rom_array(4328);
		when "1000011101001" => data_out <= rom_array(4329);
		when "1000011101010" => data_out <= rom_array(4330);
		when "1000011101011" => data_out <= rom_array(4331);
		when "1000011101100" => data_out <= rom_array(4332);
		when "1000011101101" => data_out <= rom_array(4333);
		when "1000011101110" => data_out <= rom_array(4334);
		when "1000011101111" => data_out <= rom_array(4335);
		when "1000011110000" => data_out <= rom_array(4336);
		when "1000011110001" => data_out <= rom_array(4337);
		when "1000011110010" => data_out <= rom_array(4338);
		when "1000011110011" => data_out <= rom_array(4339);
		when "1000011110100" => data_out <= rom_array(4340);
		when "1000011110101" => data_out <= rom_array(4341);
		when "1000011110110" => data_out <= rom_array(4342);
		when "1000011110111" => data_out <= rom_array(4343);
		when "1000011111000" => data_out <= rom_array(4344);
		when "1000011111001" => data_out <= rom_array(4345);
		when "1000011111010" => data_out <= rom_array(4346);
		when "1000011111011" => data_out <= rom_array(4347);
		when "1000011111100" => data_out <= rom_array(4348);
		when "1000011111101" => data_out <= rom_array(4349);
		when "1000011111110" => data_out <= rom_array(4350);
		when "1000011111111" => data_out <= rom_array(4351);
		when "1000100000000" => data_out <= rom_array(4352);
		when "1000100000001" => data_out <= rom_array(4353);
		when "1000100000010" => data_out <= rom_array(4354);
		when "1000100000011" => data_out <= rom_array(4355);
		when "1000100000100" => data_out <= rom_array(4356);
		when "1000100000101" => data_out <= rom_array(4357);
		when "1000100000110" => data_out <= rom_array(4358);
		when "1000100000111" => data_out <= rom_array(4359);
		when "1000100001000" => data_out <= rom_array(4360);
		when "1000100001001" => data_out <= rom_array(4361);
		when "1000100001010" => data_out <= rom_array(4362);
		when "1000100001011" => data_out <= rom_array(4363);
		when "1000100001100" => data_out <= rom_array(4364);
		when "1000100001101" => data_out <= rom_array(4365);
		when "1000100001110" => data_out <= rom_array(4366);
		when "1000100001111" => data_out <= rom_array(4367);
		when "1000100010000" => data_out <= rom_array(4368);
		when "1000100010001" => data_out <= rom_array(4369);
		when "1000100010010" => data_out <= rom_array(4370);
		when "1000100010011" => data_out <= rom_array(4371);
		when "1000100010100" => data_out <= rom_array(4372);
		when "1000100010101" => data_out <= rom_array(4373);
		when "1000100010110" => data_out <= rom_array(4374);
		when "1000100010111" => data_out <= rom_array(4375);
		when "1000100011000" => data_out <= rom_array(4376);
		when "1000100011001" => data_out <= rom_array(4377);
		when "1000100011010" => data_out <= rom_array(4378);
		when "1000100011011" => data_out <= rom_array(4379);
		when "1000100011100" => data_out <= rom_array(4380);
		when "1000100011101" => data_out <= rom_array(4381);
		when "1000100011110" => data_out <= rom_array(4382);
		when "1000100011111" => data_out <= rom_array(4383);
		when "1000100100000" => data_out <= rom_array(4384);
		when "1000100100001" => data_out <= rom_array(4385);
		when "1000100100010" => data_out <= rom_array(4386);
		when "1000100100011" => data_out <= rom_array(4387);
		when "1000100100100" => data_out <= rom_array(4388);
		when "1000100100101" => data_out <= rom_array(4389);
		when "1000100100110" => data_out <= rom_array(4390);
		when "1000100100111" => data_out <= rom_array(4391);
		when "1000100101000" => data_out <= rom_array(4392);
		when "1000100101001" => data_out <= rom_array(4393);
		when "1000100101010" => data_out <= rom_array(4394);
		when "1000100101011" => data_out <= rom_array(4395);
		when "1000100101100" => data_out <= rom_array(4396);
		when "1000100101101" => data_out <= rom_array(4397);
		when "1000100101110" => data_out <= rom_array(4398);
		when "1000100101111" => data_out <= rom_array(4399);
		when "1000100110000" => data_out <= rom_array(4400);
		when "1000100110001" => data_out <= rom_array(4401);
		when "1000100110010" => data_out <= rom_array(4402);
		when "1000100110011" => data_out <= rom_array(4403);
		when "1000100110100" => data_out <= rom_array(4404);
		when "1000100110101" => data_out <= rom_array(4405);
		when "1000100110110" => data_out <= rom_array(4406);
		when "1000100110111" => data_out <= rom_array(4407);
		when "1000100111000" => data_out <= rom_array(4408);
		when others => data_out <= (others => '0');
		end case;
	end process;
ClockProc: process (clk, rst) is
begin

if rising_edge(clk) then
	if rst = '1' then
		count <= (others => '0');
	
	elsif (ENABLE = '1') then
		if (unsigned(count) < rom_type'length) then
			count <= std_logic_vector(unsigned(count) + 1);
		else
			count <= (others => '0');
		end if;
	end if;
end if;

end process;
end Behavioral;
