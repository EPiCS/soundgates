../../../../../sndcomponents/nco/nco.vhd