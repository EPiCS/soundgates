../../../../../basic/amplifier/amplifier.vhd