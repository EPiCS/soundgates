--  ____                        _             _            
-- / ___|  ___  _   _ _ __   __| | __ _  __ _| |_ ___  ___ 
-- \___ \ / _ \| | | | '_ \ / _` |/ _` |/ _` | __/ _ \/ __|
--  ___) | (_) | |_| | | | | (_| | (_| | (_| | ||  __/\__ \
-- |____/ \___/ \__,_|_| |_|\__,_|\__, |\__,_|\__\___||___/
--                                |___/                    
-- ======================================================================
--
--   title:        VHDL module - hwt_fir
--
--   project:      PG-Soundgates
--   author:       Hendrik Hangmann, University of Paderborn
--
--   description:  Hardware thread for FIR Filter
-- ======================================================================

library ieee;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

--library proc_common_v3_00_a;
--use proc_common_v3_00_a.proc_common_pkg.all;

library reconos_v3_00_c;
use reconos_v3_00_c.reconos_pkg.all;

library soundgates_v1_00_a;
use soundgates_v1_00_a.soundgates_common_pkg.all;
use soundgates_v1_00_a.soundgates_reconos_pkg.all;

entity hwt_fir is
    generic(
    	SND_COMP_CLK_FREQ   : integer := 100_000_000;
		FIR_ORDER			  : integer := 7  -- 8 coefficients
	);
   port (
		-- OSIF FIFO ports
		OSIF_FIFO_Sw2Hw_Data    : in  std_logic_vector(31 downto 0);
		OSIF_FIFO_Sw2Hw_Fill    : in  std_logic_vector(15 downto 0);
		OSIF_FIFO_Sw2Hw_Empty   : in  std_logic;
		OSIF_FIFO_Sw2Hw_RE      : out std_logic;

		OSIF_FIFO_Hw2Sw_Data    : out std_logic_vector(31 downto 0);
		OSIF_FIFO_Hw2Sw_Rem     : in  std_logic_vector(15 downto 0);
		OSIF_FIFO_Hw2Sw_Full    : in  std_logic;
		OSIF_FIFO_Hw2Sw_WE      : out std_logic;

		-- MEMIF FIFO ports
		MEMIF_FIFO_Hwt2Mem_Data    : out std_logic_vector(31 downto 0);
		MEMIF_FIFO_Hwt2Mem_Rem     : in  std_logic_vector(15 downto 0);
		MEMIF_FIFO_Hwt2Mem_Full    : in  std_logic;
		MEMIF_FIFO_Hwt2Mem_WE      : out std_logic;

		MEMIF_FIFO_Mem2Hwt_Data    : in  std_logic_vector(31 downto 0);
		MEMIF_FIFO_Mem2Hwt_Fill    : in  std_logic_vector(15 downto 0);
		MEMIF_FIFO_Mem2Hwt_Empty   : in  std_logic;
		MEMIF_FIFO_Mem2Hwt_RE      : out std_logic;

		HWT_Clk   : in  std_logic;
		HWT_Rst   : in  std_logic
    );
end hwt_fir;

architecture Behavioral of hwt_fir is

    ----------------------------------------------------------------
    -- Subcomponent declarations
    ----------------------------------------------------------------

   -- ?? Was macht das hier?
   --  memif_read_word(i_memif, o_memif, rlse_amp_addr, rlse_amp, done);
   --                 if done then
   --                     refresh_state <= "0";
   --                     state <= STATE_PROCESS;
 
    signal clk   : std_logic;
	signal rst   : std_logic;

-- ReconOS Stuff
    signal i_osif   : i_osif_t;
    signal o_osif   : o_osif_t;
    signal i_memif  : i_memif_t;
    signal o_memif  : o_memif_t;
    
    signal i_ram    : i_ram_t;
    signal o_ram    : o_ram_t;
    
    constant MBOX_START   : std_logic_vector(31 downto 0) := x"00000000";
    constant MBOX_FINISH  : std_logic_vector(31 downto 0) := x"00000001";
-- /ReconOS Stuff

    type STATE_TYPE is (STATE_INIT, STATE_INIT_ADDRESSES, STATE_READ_COEFFICIENTS_ADRESSES, STATE_READ, STATE_WAITING, STATE_PROCESS, STATE_WRITE_MEM, STATE_NOTIFY, STATE_EXIT);
    signal state    : STATE_TYPE;
	 
	 
    
    ----------------------------------------------------------------
    -- Common sound component signals, constants and types
    ----------------------------------------------------------------
    
    constant C_MAX_SAMPLE_COUNT : integer := 64;
    
   	-- define size of local RAM here
	constant C_LOCAL_RAM_SIZE          : integer := C_MAX_SAMPLE_COUNT;
	constant C_LOCAL_RAM_ADDRESS_WIDTH : integer := 6;--clog2(C_LOCAL_RAM_SIZE);
	constant C_LOCAL_RAM_SIZE_IN_BYTES : integer := 4*C_LOCAL_RAM_SIZE;

    type LOCAL_MEMORY_T is array (0 to C_LOCAL_RAM_SIZE-1) of std_logic_vector(31 downto 0);
        
    signal o_RAMAddr_fir : std_logic_vector(0 to C_LOCAL_RAM_ADDRESS_WIDTH-1);
	signal o_RAMData_fir : std_logic_vector(0 to 31);   -- fir to local ram
	signal i_RAMData_fir : std_logic_vector(0 to 31);   -- local ram to fir
    signal o_RAMWE_fir   : std_logic;
	
  	signal o_RAMAddr_reconos   : std_logic_vector(0 to C_LOCAL_RAM_ADDRESS_WIDTH-1);
	signal o_RAMAddr_reconos_2 : std_logic_vector(0 to 31);
	signal o_RAMData_reconos   : std_logic_vector(0 to 31);
	signal o_RAMWE_reconos     : std_logic;
	signal i_RAMData_reconos   : std_logic_vector(0 to 31);
    
    signal osif_ctrl_signal : std_logic_vector(31 downto 0);
    signal ignore : std_logic_vector(31 downto 0);
    
    
    constant o_RAMAddr_max : std_logic_vector(0 to C_LOCAL_RAM_ADDRESS_WIDTH-1) := (others=>'1');

	shared variable local_ram : LOCAL_MEMORY_T;
    
    signal snd_comp_header : snd_comp_header_msg_t;  -- common sound component header
       
    signal sample_count            : unsigned(15 downto 0) := to_unsigned(C_MAX_SAMPLE_COUNT, 16);
    
    ----------------------------------------------------------------
    -- Component dependent signals
    ----------------------------------------------------------------
    signal fir_ce          : std_logic;           -- fir clock enable (like a start/stop signal)
    
    signal input_data       : signed(31 downto 0);
    signal fir_data         : signed(31 downto 0);

	 signal count 			    : signed (31 downto 0);
	 
	 signal process_state    : integer range 0 to 2;
	 
    type mem32 is array (natural range <>) of std_logic_vector(31 downto 0);
	 type smem32 is array (natural range <>) of signed(31 downto 0);
	 type mem64 is array (natural range <>) of signed(63 downto 0);
	 
    signal coeffs_mem32 : mem32(FIR_ORDER downto 0);
    signal coeff_index : signed(31 downto 0);

    signal inputs_mem32 : mem32(FIR_ORDER downto 0);

    signal mult_mem64 : mem64(FIR_ORDER downto 0);
	 
	 signal init_state : integer range 0 to 1;
	 
	 signal coefficients_addr : mem32(FIR_ORDER downto 0);
	 signal coefficients : mem32(FIR_ORDER downto 0);
	 
	 signal buffer_states_addr : mem32(FIR_ORDER downto 0);
	 signal buffer_states : mem32(FIR_ORDER downto 0);
	 
	 signal opt_arg : std_logic_vector(31 downto 0);
	 signal coefficient_count_addr : std_logic_vector(31 downto 0);
	 signal coefficient_count : std_logic_vector(31 downto 0);
	 
	 signal addr_counter : integer range 0 to FIR_ORDER + 1;
	 
	 signal input_mem32 : smem32(FIR_ORDER downto 0);
	 signal output_mem64 : mem64(FIR_ORDER downto 0);
	 
	 signal fir_data64 : signed(63 downto 0);
	     
    ----------------------------------------------------------------
    -- OS Communication
    ----------------------------------------------------------------
    
    constant fir_START : std_logic_vector(31 downto 0) := x"0000000F";
    constant fir_EXIT  : std_logic_vector(31 downto 0) := x"000000F0";
    
    constant C_START_BANG : std_logic_vector(31 downto 0) := x"00000001";
    constant C_STOP_BANG  : std_logic_vector(31 downto 0) := x"FFFFFFFF";

begin
    -----------------------------------
    -- Hard wirings
    -----------------------------------
    clk <= HWT_Clk;
	rst <= HWT_Rst;
--    o_RAMData_fir <= std_logic_vector(fir_data);
    
    
    
    o_RAMAddr_reconos(0 to C_LOCAL_RAM_ADDRESS_WIDTH-1) <= o_RAMAddr_reconos_2((32-C_LOCAL_RAM_ADDRESS_WIDTH) to 31);
    
        
    -- ReconOS Stuff
    osif_setup (
            i_osif,
            o_osif,
            OSIF_FIFO_Sw2Hw_Data,
            OSIF_FIFO_Sw2Hw_Fill,
            OSIF_FIFO_Sw2Hw_Empty,
            OSIF_FIFO_Hw2Sw_Rem,
            OSIF_FIFO_Hw2Sw_Full,
            OSIF_FIFO_Sw2Hw_RE,
            OSIF_FIFO_Hw2Sw_Data,
            OSIF_FIFO_Hw2Sw_WE
        );
                    
    memif_setup (
            i_memif,
            o_memif,
            MEMIF_FIFO_Mem2Hwt_Data,
            MEMIF_FIFO_Mem2Hwt_Fill,
            MEMIF_FIFO_Mem2Hwt_Empty,
            MEMIF_FIFO_Hwt2Mem_Rem,
            MEMIF_FIFO_Hwt2Mem_Full,
            MEMIF_FIFO_Mem2Hwt_RE,
            MEMIF_FIFO_Hwt2Mem_Data,
            MEMIF_FIFO_Hwt2Mem_WE
        );

    ram_setup (
		i_ram,
		o_ram,
		o_RAMAddr_reconos_2,
		o_RAMWE_reconos,
		o_RAMData_reconos,
		i_RAMData_reconos
	);
            
    -- /ReconOS Stuff
            
    local_ram_ctrl_1 : process (clk) is
	begin
		if (rising_edge(clk)) then
			if (o_RAMWE_reconos = '1') then
				local_ram(to_integer(unsigned(o_RAMAddr_reconos))) := o_RAMData_reconos;
			else
				i_RAMData_reconos <= local_ram(to_integer(unsigned(o_RAMAddr_reconos)));
			end if;
		end if;
	end process;
    
    local_ram_ctrl_2 : process (clk) is
	begin
		if (rising_edge(clk)) then		
			if (o_RAMWE_fir = '1') then
				local_ram(to_integer(unsigned(o_RAMAddr_fir))) := o_RAMData_fir;
         else      -- else needed, because fir is consuming samples
				i_RAMData_fir <= local_ram(to_integer(unsigned(o_RAMAddr_fir)));
			end if;
		end if;
	end process;
    
    
    fir_CTRL_FSM_PROC : process (clk, rst, o_osif, o_memif) is
        variable done : boolean;            
    begin
        if rst = '1' then
                    
            osif_reset(o_osif);
				memif_reset(o_memif);           
            ram_reset(o_ram);
            addr_counter <= 0;
            state           <= STATE_INIT;
            osif_ctrl_signal <= (others => '0');

            o_RAMWE_fir<= '0';

				count <= (others => '0');
            
            done := False;
				
				init_state <= 0;
              
            sample_count    <= to_unsigned(0, 16);
        elsif rising_edge(clk) then
            
            fir_ce      <= '0';
            o_RAMWE_fir <= '0';
            osif_ctrl_signal <= ( others => '0');
            
            case state is            
            -- INIT State gets the address of the header struct
            when STATE_INIT =>               
                snd_comp_get_header(i_osif, o_osif, i_memif, o_memif, snd_comp_header, done);         
                if done then
                    -- Initialize your signals
                        opt_arg  <= snd_comp_header.opt_arg_addr;
								coefficient_count_addr <= opt_arg; -- address to number of coefficients
								
                        state <= STATE_INIT_ADDRESSES;
                end if;    
					 
            when STATE_INIT_ADDRESSES =>
					case init_state is
					when 0 =>
						-- get number of coefficients
						memif_read_word(i_memif, o_memif, coefficient_count_addr, coefficient_count, done);
					  if done then
							init_state <= 1;
					  end if;
					  
					 when 1 =>					 
					 
					    coefficients_addr(addr_counter) <= std_logic_vector(unsigned(snd_comp_header.opt_arg_addr) + 4*(addr_counter+1));
						 addr_counter <= addr_counter + 1;
						 if addr_counter >= to_integer(signed(coefficient_count)) then
							init_state <= 0;
							state <= STATE_WAITING;
						 else
							init_state <= 1;
						 end if;
--						 for i in 0 to to_integer(signed(coefficient_count)) - 1 loop
--							  coefficients_addr(i) <= std_logic_vector(unsigned(snd_comp_header.opt_arg_addr) + 4*(i+1));
--							  --address to actual coefficients
--						 end loop;
--						 init_state <= 0;
--						 state <= STATE_WAITING;
					 
--					 when "2" =>
--					 
--						 buffer_state_count_addr <= std_logic_vector(unsigned(opt_arg + 4*(to_integer(signed(coefficient_count)) + 2)));
--						 -- address to number of buffer states
--						 
--						 for i in 0 to to_integer(signed(buffer_state_count_addr)) - 1 loop
--							  buffer_states_addr(i) <= std_logic_vector(unsigned(snd_comp_header.opt_arg_addr) + unsigned(4*(i+1)));
--							  --address to actual buffer states
--						 end loop;
						 
					end case;

            when STATE_WAITING =>
                -- Software process "Synthesizer" sends the start signal via mbox_start
                osif_mbox_get(i_osif, o_osif, MBOX_START, osif_ctrl_signal, done);
                if done then
                    if osif_ctrl_signal = fir_START then
                        state        <= STATE_READ_COEFFICIENTS_ADRESSES;

                    elsif osif_ctrl_signal = fir_EXIT then
                        
                        state   <= STATE_EXIT;

                    end if;    
                end if;
           					
			  
			  when STATE_READ_COEFFICIENTS_ADRESSES =>
			  -- read adresses to the fir coefficients values
                memif_read_word(i_memif, o_memif, coefficients_addr(to_integer(count)), coefficients(to_integer(count)), done);
					  if done then
						-- write values to FIR component
							count <= count + 1;
							
							if count > signed(coefficient_count) then
							  state <= STATE_READ;
							  count <= (others => '0');
							else
								state <= STATE_READ_COEFFICIENTS_ADRESSES;
							end if;
					  end if;
			  
--			 when STATE_READ_BUFFER_STATE_ADRESSES =>
--			 -- read adresses to the fir buffer state values
--                memif_read_word(i_memif, o_memif, buffer_states_addr(to_integer(count)), buffer_states(to_integer(count)), done);
--					  if done then
--							-- write values to the FIR component
--							count <= count + 1;
--							
--							config_buffer_state_valid <= '1';
--							config_buffer_state_index <= count;
--							config_buffer_state_data <= buffer_states(to_integer(count));
--							
--							if count > signed(buffer_states) then
--							  state <= STATE_READ;
--							  count <= (others => '0');
--							else
--								state <= STATE_READ_BUFFER_STATE_ADRESSES;
--							end if;
--					  end if;
			  
			  when STATE_READ => 
					-- store input samples in local ram
					memif_read(i_ram,o_ram,i_memif,o_memif,snd_comp_header.source_addr,X"00000000",std_logic_vector(to_unsigned(C_LOCAL_RAM_SIZE_IN_BYTES,24)),done);
					if done then
						state <= STATE_PROCESS;
					end if;
			 
            when STATE_PROCESS =>
                if sample_count < to_unsigned(C_MAX_SAMPLE_COUNT, 16) then
                    case process_state is

                    when 0 => 
								for i in 0 to FIR_ORDER - 1 loop
									input_mem32(i + 1) <= input_mem32(i);
								end loop;
								
								input_mem32(0) <= signed(i_RAMData_fir);
								
								for i in 0 to FIR_ORDER loop
									output_mem64(i) <= signed(coefficients(i)) * input_mem32(FIR_ORDER - i);
									fir_data64 <= fir_data64 + output_mem64(i);
								end loop;
								
								process_state  <= 1;

                    when 1 =>
								fir_data <= fir_data64(31 downto 0);
								o_RAMData_fir <= std_logic_vector(fir_data);
                        o_RAMWE_fir   <= '1';
								count <= count + 1;
                        process_state  <= 2;       

                    when 2 =>
                        o_RAMWE_fir   <= '0';
								fir_data64 <= (others => '0');
                        o_RAMAddr_fir <= std_logic_vector(unsigned(o_RAMAddr_fir) + 1);
                        sample_count  <= sample_count + 1;
								
                        process_state  <= 0;  
                    end case;

                else
                    -- Samples have been generated
                    o_RAMAddr_fir  <= (others => '0');
                    sample_count    <= to_unsigned(0, 16);
                    state <= STATE_WRITE_MEM;
                end if;


             when STATE_WRITE_MEM =>
        
                memif_write(i_ram, o_ram, i_memif, o_memif, X"00000000", snd_comp_header.dest_addr, std_logic_vector(to_unsigned(C_LOCAL_RAM_SIZE_IN_BYTES,24)), done);
                if done then
                    state <= STATE_NOTIFY;
					end if;
				
				when STATE_NOTIFY =>

                osif_mbox_put(i_osif, o_osif, MBOX_FINISH, snd_comp_header.dest_addr, ignore, done);
                if done then
                    state <= STATE_WAITING;
						end if;
                        
            when STATE_EXIT =>

                   osif_thread_exit(i_osif,o_osif);            
            end case;
        end if;
    end process;


end Behavioral;

-- ====================================
-- = RECONOS Function Library - Copy and Paste!
-- ====================================        
-- osif_mbox_put(i_osif, o_osif, MBOX_NAME, SOURCESIGNAL, ignore, done);
-- osif_mbox_get(i_osif, o_osif, MBOX_NAME, TARGETSIGNAL, done);

-- Read from shared memory:

-- Speicherzugriffe:
-- Wortzugriff:
-- memif_read_word(i_memif, o_memif, addr, TARGETSIGNAL, done);
-- memif_write_word(i_memif, o_memif, addr, SOURCESIGNAL, done);

-- Die Laenge ist bei Speicherzugriffen Byte adressiert!
-- memif_read(i_ram, o_ram, i_memif, o_memif, SRC_ADDR std_logic_vector(31 downto 0);
--            dst_addr std_logic_vector(31 downto 0);
--            BYTES std_logic_vector(23 downto 0);
--            done);
-- memif_write(i_ram, o_ram, i_memif, o_memif,
--             src_addr : in std_logic_vector(31 downto 0),
--             dst_addr : in std_logic_vector(31 downto 0);
--             len      : in std_logic_vector(23 downto 0);
--             done);

