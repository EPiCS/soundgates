../../../../basic/triangle/triangle.vhd