../../../../../basic/mul/mul.vhd