../../../../../basic/fir/fir_transposed.vhd