../../../../../basic/sawtooth/sawtooth.vhd