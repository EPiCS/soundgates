../../../../../basic/cordic/cordic.vhd